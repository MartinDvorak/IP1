
	library ieee;
use ieee.std_logic_1164.all;

architecture ./vtf_tests/backdoor-subset-4 of pattern_match is

--#################################################
-- start section fullgraph: 0

  -- state q345
  signal reg_q345        : std_logic;
  signal reg_q345_in     : std_logic;
  		

  -- state q2757
  signal reg_q2757        : std_logic;
  signal reg_q2757_in     : std_logic;
  		
  signal reg_fullgraph0       : std_logic_vector(1 downto 0);
  signal reg_fullgraph0_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph0_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph0_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph0
  --#################################################			
		
--#################################################
-- start section fullgraph: 1

  -- state q565
  signal reg_q565        : std_logic;
  signal reg_q565_in     : std_logic;
  		

  -- state q587
  signal reg_q587        : std_logic;
  signal reg_q587_in     : std_logic;
  		

  -- state q1323
  signal reg_q1323        : std_logic;
  signal reg_q1323_in     : std_logic;
  		

  -- state q494
  signal reg_q494        : std_logic;
  signal reg_q494_in     : std_logic;
  		

  -- state q2526
  signal reg_q2526        : std_logic;
  signal reg_q2526_in     : std_logic;
  		

  -- state q377
  signal reg_q377        : std_logic;
  signal reg_q377_in     : std_logic;
  		

  -- state q185
  signal reg_q185        : std_logic;
  signal reg_q185_in     : std_logic;
  		

  -- state q522
  signal reg_q522        : std_logic;
  signal reg_q522_in     : std_logic;
  		

  -- state q1719
  signal reg_q1719        : std_logic;
  signal reg_q1719_in     : std_logic;
  		

  -- state q2736
  signal reg_q2736        : std_logic;
  signal reg_q2736_in     : std_logic;
  		

  -- state q2738
  signal reg_q2738        : std_logic;
  signal reg_q2738_in     : std_logic;
  		

  -- state q876
  signal reg_q876        : std_logic;
  signal reg_q876_in     : std_logic;
  		

  -- state q942
  signal reg_q942        : std_logic;
  signal reg_q942_in     : std_logic;
  		

  -- state q2524
  signal reg_q2524        : std_logic;
  signal reg_q2524_in     : std_logic;
  		

  -- state q359
  signal reg_q359        : std_logic;
  signal reg_q359_in     : std_logic;
  		

  -- state q2034
  signal reg_q2034        : std_logic;
  signal reg_q2034_in     : std_logic;
  		

  -- state q2036
  signal reg_q2036        : std_logic;
  signal reg_q2036_in     : std_logic;
  		

  -- state q2623
  signal reg_q2623        : std_logic;
  signal reg_q2623_in     : std_logic;
  		

  -- state q675
  signal reg_q675        : std_logic;
  signal reg_q675_in     : std_logic;
  		

  -- state q149
  signal reg_q149        : std_logic;
  signal reg_q149_in     : std_logic;
  		

  -- state q151
  signal reg_q151        : std_logic;
  signal reg_q151_in     : std_logic;
  		

  -- state q480
  signal reg_q480        : std_logic;
  signal reg_q480_in     : std_logic;
  		

  -- state q40
  signal reg_q40        : std_logic;
  signal reg_q40_in     : std_logic;
  		

  -- state q732
  signal reg_q732        : std_logic;
  signal reg_q732_in     : std_logic;
  		

  -- state q1357
  signal reg_q1357        : std_logic;
  signal reg_q1357_in     : std_logic;
  		

  -- state q107
  signal reg_q107        : std_logic;
  signal reg_q107_in     : std_logic;
  		

  -- state q2290
  signal reg_q2290        : std_logic;
  signal reg_q2290_in     : std_logic;
  		

  -- state q2312
  signal reg_q2312        : std_logic;
  signal reg_q2312_in     : std_logic;
  		

  -- state q2314
  signal reg_q2314        : std_logic;
  signal reg_q2314_in     : std_logic;
  		

  -- state q2038
  signal reg_q2038        : std_logic;
  signal reg_q2038_in     : std_logic;
  		

  -- state q1502
  signal reg_q1502        : std_logic;
  signal reg_q1502_in     : std_logic;
  		

  -- state q1504
  signal reg_q1504        : std_logic;
  signal reg_q1504_in     : std_logic;
  		

  -- state q1996
  signal reg_q1996        : std_logic;
  signal reg_q1996_in     : std_logic;
  		

  -- state q1998
  signal reg_q1998        : std_logic;
  signal reg_q1998_in     : std_logic;
  		

  -- state q2006
  signal reg_q2006        : std_logic;
  signal reg_q2006_in     : std_logic;
  		

  -- state q2008
  signal reg_q2008        : std_logic;
  signal reg_q2008_in     : std_logic;
  		

  -- state q817
  signal reg_q817        : std_logic;
  signal reg_q817_in     : std_logic;
  		

  -- state q1128
  signal reg_q1128        : std_logic;
  signal reg_q1128_in     : std_logic;
  		

  -- state q1130
  signal reg_q1130        : std_logic;
  signal reg_q1130_in     : std_logic;
  		

  -- state q2050
  signal reg_q2050        : std_logic;
  signal reg_q2050_in     : std_logic;
  		

  -- state q2054
  signal reg_q2054        : std_logic;
  signal reg_q2054_in     : std_logic;
  		

  -- state q210
  signal reg_q210        : std_logic;
  signal reg_q210_in     : std_logic;
  		

  -- state q369
  signal reg_q369        : std_logic;
  signal reg_q369_in     : std_logic;
  		

  -- state q712
  signal reg_q712        : std_logic;
  signal reg_q712_in     : std_logic;
  		

  -- state q714
  signal reg_q714        : std_logic;
  signal reg_q714_in     : std_logic;
  		

  -- state q1924
  signal reg_q1924        : std_logic;
  signal reg_q1924_in     : std_logic;
  		

  -- state q1926
  signal reg_q1926        : std_logic;
  signal reg_q1926_in     : std_logic;
  		

  -- state q1709
  signal reg_q1709        : std_logic;
  signal reg_q1709_in     : std_logic;
  		

  -- state q1711
  signal reg_q1711        : std_logic;
  signal reg_q1711_in     : std_logic;
  		

  -- state q2280
  signal reg_q2280        : std_logic;
  signal reg_q2280_in     : std_logic;
  		

  -- state q2282
  signal reg_q2282        : std_logic;
  signal reg_q2282_in     : std_logic;
  		

  -- state q282
  signal reg_q282        : std_logic;
  signal reg_q282_in     : std_logic;
  		

  -- state q284
  signal reg_q284        : std_logic;
  signal reg_q284_in     : std_logic;
  		

  -- state q2387
  signal reg_q2387        : std_logic;
  signal reg_q2387_in     : std_logic;
  		

  -- state q2389
  signal reg_q2389        : std_logic;
  signal reg_q2389_in     : std_logic;
  		

  -- state q1500
  signal reg_q1500        : std_logic;
  signal reg_q1500_in     : std_logic;
  		

  -- state q2744
  signal reg_q2744        : std_logic;
  signal reg_q2744_in     : std_logic;
  		

  -- state q2746
  signal reg_q2746        : std_logic;
  signal reg_q2746_in     : std_logic;
  		

  -- state q1915
  signal reg_q1915        : std_logic;
  signal reg_q1915_in     : std_logic;
  		

  -- state q1498
  signal reg_q1498        : std_logic;
  signal reg_q1498_in     : std_logic;
  		

  -- state q218
  signal reg_q218        : std_logic;
  signal reg_q218_in     : std_logic;
  		

  -- state q220
  signal reg_q220        : std_logic;
  signal reg_q220_in     : std_logic;
  		

  -- state q1990
  signal reg_q1990        : std_logic;
  signal reg_q1990_in     : std_logic;
  		

  -- state q1992
  signal reg_q1992        : std_logic;
  signal reg_q1992_in     : std_logic;
  		

  -- state q2020
  signal reg_q2020        : std_logic;
  signal reg_q2020_in     : std_logic;
  		

  -- state q2022
  signal reg_q2022        : std_logic;
  signal reg_q2022_in     : std_logic;
  		

  -- state q214
  signal reg_q214        : std_logic;
  signal reg_q214_in     : std_logic;
  		

  -- state q2712
  signal reg_q2712        : std_logic;
  signal reg_q2712_in     : std_logic;
  		

  -- state q2714
  signal reg_q2714        : std_logic;
  signal reg_q2714_in     : std_logic;
  		

  -- state q2032
  signal reg_q2032        : std_logic;
  signal reg_q2032_in     : std_logic;
  		

  -- state q1945
  signal reg_q1945        : std_logic;
  signal reg_q1945_in     : std_logic;
  		

  -- state q1947
  signal reg_q1947        : std_logic;
  signal reg_q1947_in     : std_logic;
  		

  -- state q124
  signal reg_q124        : std_logic;
  signal reg_q124_in     : std_logic;
  		

  -- state q126
  signal reg_q126        : std_logic;
  signal reg_q126_in     : std_logic;
  		

  -- state q2272
  signal reg_q2272        : std_logic;
  signal reg_q2272_in     : std_logic;
  		

  -- state q2274
  signal reg_q2274        : std_logic;
  signal reg_q2274_in     : std_logic;
  		

  -- state q42
  signal reg_q42        : std_logic;
  signal reg_q42_in     : std_logic;
  		

  -- state q44
  signal reg_q44        : std_logic;
  signal reg_q44_in     : std_logic;
  		

  -- state q2028
  signal reg_q2028        : std_logic;
  signal reg_q2028_in     : std_logic;
  		

  -- state q2030
  signal reg_q2030        : std_logic;
  signal reg_q2030_in     : std_logic;
  		

  -- state q1315
  signal reg_q1315        : std_logic;
  signal reg_q1315_in     : std_logic;
  		

  -- state q2704
  signal reg_q2704        : std_logic;
  signal reg_q2704_in     : std_logic;
  		

  -- state q2706
  signal reg_q2706        : std_logic;
  signal reg_q2706_in     : std_logic;
  		

  -- state q1994
  signal reg_q1994        : std_logic;
  signal reg_q1994_in     : std_logic;
  		

  -- state q1804
  signal reg_q1804        : std_logic;
  signal reg_q1804_in     : std_logic;
  		

  -- state q1806
  signal reg_q1806        : std_logic;
  signal reg_q1806_in     : std_logic;
  		

  -- state q698
  signal reg_q698        : std_logic;
  signal reg_q698_in     : std_logic;
  		

  -- state q700
  signal reg_q700        : std_logic;
  signal reg_q700_in     : std_logic;
  		

  -- state q2617
  signal reg_q2617        : std_logic;
  signal reg_q2617_in     : std_logic;
  		

  -- state q768
  signal reg_q768        : std_logic;
  signal reg_q768_in     : std_logic;
  		

  -- state q2752
  signal reg_q2752        : std_logic;
  signal reg_q2752_in     : std_logic;
  		

  -- state q2754
  signal reg_q2754        : std_logic;
  signal reg_q2754_in     : std_logic;
  		

  -- state q1701
  signal reg_q1701        : std_logic;
  signal reg_q1701_in     : std_logic;
  		

  -- state q1703
  signal reg_q1703        : std_logic;
  signal reg_q1703_in     : std_logic;
  		

  -- state q120
  signal reg_q120        : std_logic;
  signal reg_q120_in     : std_logic;
  		

  -- state q122
  signal reg_q122        : std_logic;
  signal reg_q122_in     : std_logic;
  		

  -- state q2726
  signal reg_q2726        : std_logic;
  signal reg_q2726_in     : std_logic;
  		

  -- state q2728
  signal reg_q2728        : std_logic;
  signal reg_q2728_in     : std_logic;
  		

  -- state q2040
  signal reg_q2040        : std_logic;
  signal reg_q2040_in     : std_logic;
  		

  -- state q2042
  signal reg_q2042        : std_logic;
  signal reg_q2042_in     : std_logic;
  		

  -- state q208
  signal reg_q208        : std_logic;
  signal reg_q208_in     : std_logic;
  		

  -- state q1126
  signal reg_q1126        : std_logic;
  signal reg_q1126_in     : std_logic;
  		

  -- state q1212
  signal reg_q1212        : std_logic;
  signal reg_q1212_in     : std_logic;
  		

  -- state q1214
  signal reg_q1214        : std_logic;
  signal reg_q1214_in     : std_logic;
  		

  -- state q2316
  signal reg_q2316        : std_logic;
  signal reg_q2316_in     : std_logic;
  		

  -- state q2018
  signal reg_q2018        : std_logic;
  signal reg_q2018_in     : std_logic;
  		

  -- state q355
  signal reg_q355        : std_logic;
  signal reg_q355_in     : std_logic;
  		

  -- state q357
  signal reg_q357        : std_logic;
  signal reg_q357_in     : std_logic;
  		

  -- state q776
  signal reg_q776        : std_logic;
  signal reg_q776_in     : std_logic;
  		

  -- state q778
  signal reg_q778        : std_logic;
  signal reg_q778_in     : std_logic;
  		

  -- state q58
  signal reg_q58        : std_logic;
  signal reg_q58_in     : std_logic;
  		

  -- state q60
  signal reg_q60        : std_logic;
  signal reg_q60_in     : std_logic;
  		

  -- state q1183
  signal reg_q1183        : std_logic;
  signal reg_q1183_in     : std_logic;
  		

  -- state q718
  signal reg_q718        : std_logic;
  signal reg_q718_in     : std_logic;
  		

  -- state q972
  signal reg_q972        : std_logic;
  signal reg_q972_in     : std_logic;
  		

  -- state q974
  signal reg_q974        : std_logic;
  signal reg_q974_in     : std_logic;
  		

  -- state q2012
  signal reg_q2012        : std_logic;
  signal reg_q2012_in     : std_logic;
  		

  -- state q2014
  signal reg_q2014        : std_logic;
  signal reg_q2014_in     : std_logic;
  		

  -- state q2383
  signal reg_q2383        : std_logic;
  signal reg_q2383_in     : std_logic;
  		

  -- state q2385
  signal reg_q2385        : std_logic;
  signal reg_q2385_in     : std_logic;
  		

  -- state q782
  signal reg_q782        : std_logic;
  signal reg_q782_in     : std_logic;
  		

  -- state q784
  signal reg_q784        : std_logic;
  signal reg_q784_in     : std_logic;
  		

  -- state q501
  signal reg_q501        : std_logic;
  signal reg_q501_in     : std_logic;
  		

  -- state q1707
  signal reg_q1707        : std_logic;
  signal reg_q1707_in     : std_logic;
  		

  -- state q1949
  signal reg_q1949        : std_logic;
  signal reg_q1949_in     : std_logic;
  		

  -- state q52
  signal reg_q52        : std_logic;
  signal reg_q52_in     : std_logic;
  		

  -- state q54
  signal reg_q54        : std_logic;
  signal reg_q54_in     : std_logic;
  		

  -- state q2621
  signal reg_q2621        : std_logic;
  signal reg_q2621_in     : std_logic;
  		

  -- state q238
  signal reg_q238        : std_logic;
  signal reg_q238_in     : std_logic;
  		

  -- state q240
  signal reg_q240        : std_logic;
  signal reg_q240_in     : std_logic;
  		

  -- state q716
  signal reg_q716        : std_logic;
  signal reg_q716_in     : std_logic;
  		

  -- state q1187
  signal reg_q1187        : std_logic;
  signal reg_q1187_in     : std_logic;
  		

  -- state q1189
  signal reg_q1189        : std_logic;
  signal reg_q1189_in     : std_logic;
  		

  -- state q2597
  signal reg_q2597        : std_logic;
  signal reg_q2597_in     : std_logic;
  		

  -- state q2599
  signal reg_q2599        : std_logic;
  signal reg_q2599_in     : std_logic;
  		

  -- state q141
  signal reg_q141        : std_logic;
  signal reg_q141_in     : std_logic;
  		

  -- state q143
  signal reg_q143        : std_logic;
  signal reg_q143_in     : std_logic;
  		

  -- state q1768
  signal reg_q1768        : std_logic;
  signal reg_q1768_in     : std_logic;
  		

  -- state q1770
  signal reg_q1770        : std_logic;
  signal reg_q1770_in     : std_logic;
  		

  -- state q2288
  signal reg_q2288        : std_logic;
  signal reg_q2288_in     : std_logic;
  		

  -- state q2000
  signal reg_q2000        : std_logic;
  signal reg_q2000_in     : std_logic;
  		

  -- state q1717
  signal reg_q1717        : std_logic;
  signal reg_q1717_in     : std_logic;
  		

  -- state q2225
  signal reg_q2225        : std_logic;
  signal reg_q2225_in     : std_logic;
  		

  -- state q2227
  signal reg_q2227        : std_logic;
  signal reg_q2227_in     : std_logic;
  		

  -- state q50
  signal reg_q50        : std_logic;
  signal reg_q50_in     : std_logic;
  		

  -- state q557
  signal reg_q557        : std_logic;
  signal reg_q557_in     : std_logic;
  		

  -- state q559
  signal reg_q559        : std_logic;
  signal reg_q559_in     : std_logic;
  		

  -- state q478
  signal reg_q478        : std_logic;
  signal reg_q478_in     : std_logic;
  		

  -- state q2619
  signal reg_q2619        : std_logic;
  signal reg_q2619_in     : std_logic;
  		

  -- state q2004
  signal reg_q2004        : std_logic;
  signal reg_q2004_in     : std_logic;
  		

  -- state q212
  signal reg_q212        : std_logic;
  signal reg_q212_in     : std_logic;
  		

  -- state q2276
  signal reg_q2276        : std_logic;
  signal reg_q2276_in     : std_logic;
  		

  -- state q2278
  signal reg_q2278        : std_logic;
  signal reg_q2278_in     : std_logic;
  		

  -- state q1778
  signal reg_q1778        : std_logic;
  signal reg_q1778_in     : std_logic;
  		

  -- state q1780
  signal reg_q1780        : std_logic;
  signal reg_q1780_in     : std_logic;
  		

  -- state q2264
  signal reg_q2264        : std_logic;
  signal reg_q2264_in     : std_logic;
  		

  -- state q2266
  signal reg_q2266        : std_logic;
  signal reg_q2266_in     : std_logic;
  		

  -- state q1136
  signal reg_q1136        : std_logic;
  signal reg_q1136_in     : std_logic;
  		

  -- state q69
  signal reg_q69        : std_logic;
  signal reg_q69_in     : std_logic;
  		

  -- state q71
  signal reg_q71        : std_logic;
  signal reg_q71_in     : std_logic;
  		

  -- state q171
  signal reg_q171        : std_logic;
  signal reg_q171_in     : std_logic;
  		

  -- state q1721
  signal reg_q1721        : std_logic;
  signal reg_q1721_in     : std_logic;
  		

  -- state q2016
  signal reg_q2016        : std_logic;
  signal reg_q2016_in     : std_logic;
  		

  -- state q1100
  signal reg_q1100        : std_logic;
  signal reg_q1100_in     : std_logic;
  		

  -- state q1102
  signal reg_q1102        : std_logic;
  signal reg_q1102_in     : std_logic;
  		

  -- state q722
  signal reg_q722        : std_logic;
  signal reg_q722_in     : std_logic;
  		

  -- state q724
  signal reg_q724        : std_logic;
  signal reg_q724_in     : std_logic;
  		

  -- state q1073
  signal reg_q1073        : std_logic;
  signal reg_q1073_in     : std_logic;
  		

  -- state q1075
  signal reg_q1075        : std_logic;
  signal reg_q1075_in     : std_logic;
  		

  -- state q2044
  signal reg_q2044        : std_logic;
  signal reg_q2044_in     : std_logic;
  		

  -- state q2046
  signal reg_q2046        : std_logic;
  signal reg_q2046_in     : std_logic;
  		

  -- state q258
  signal reg_q258        : std_logic;
  signal reg_q258_in     : std_logic;
  		

  -- state q260
  signal reg_q260        : std_logic;
  signal reg_q260_in     : std_logic;
  		

  -- state q236
  signal reg_q236        : std_logic;
  signal reg_q236_in     : std_logic;
  		

  -- state q1800
  signal reg_q1800        : std_logic;
  signal reg_q1800_in     : std_logic;
  		

  -- state q1802
  signal reg_q1802        : std_logic;
  signal reg_q1802_in     : std_logic;
  		

  -- state q145
  signal reg_q145        : std_logic;
  signal reg_q145_in     : std_logic;
  		

  -- state q1723
  signal reg_q1723        : std_logic;
  signal reg_q1723_in     : std_logic;
  		

  -- state q511
  signal reg_q511        : std_logic;
  signal reg_q511_in     : std_logic;
  		

  -- state q1010
  signal reg_q1010        : std_logic;
  signal reg_q1010_in     : std_logic;
  		

  -- state q555
  signal reg_q555        : std_logic;
  signal reg_q555_in     : std_logic;
  		

  -- state q167
  signal reg_q167        : std_logic;
  signal reg_q167_in     : std_logic;
  		

  -- state q169
  signal reg_q169        : std_logic;
  signal reg_q169_in     : std_logic;
  		

  -- state q2304
  signal reg_q2304        : std_logic;
  signal reg_q2304_in     : std_logic;
  		

  -- state q2306
  signal reg_q2306        : std_logic;
  signal reg_q2306_in     : std_logic;
  		

  -- state q2223
  signal reg_q2223        : std_logic;
  signal reg_q2223_in     : std_logic;
  		

  -- state q1171
  signal reg_q1171        : std_logic;
  signal reg_q1171_in     : std_logic;
  		

  -- state q1173
  signal reg_q1173        : std_logic;
  signal reg_q1173_in     : std_logic;
  		

  -- state q1520
  signal reg_q1520        : std_logic;
  signal reg_q1520_in     : std_logic;
  		

  -- state q147
  signal reg_q147        : std_logic;
  signal reg_q147_in     : std_logic;
  		

  -- state q79
  signal reg_q79        : std_logic;
  signal reg_q79_in     : std_logic;
  		

  -- state q81
  signal reg_q81        : std_logic;
  signal reg_q81_in     : std_logic;
  		

  -- state q242
  signal reg_q242        : std_logic;
  signal reg_q242_in     : std_logic;
  		

  -- state q244
  signal reg_q244        : std_logic;
  signal reg_q244_in     : std_logic;
  		

  -- state q1911
  signal reg_q1911        : std_logic;
  signal reg_q1911_in     : std_logic;
  		

  -- state q1913
  signal reg_q1913        : std_logic;
  signal reg_q1913_in     : std_logic;
  		

  -- state q190
  signal reg_q190        : std_logic;
  signal reg_q190_in     : std_logic;
  		

  -- state q2024
  signal reg_q2024        : std_logic;
  signal reg_q2024_in     : std_logic;
  		

  -- state q2026
  signal reg_q2026        : std_logic;
  signal reg_q2026_in     : std_logic;
  		

  -- state q1159
  signal reg_q1159        : std_logic;
  signal reg_q1159_in     : std_logic;
  		

  -- state q1161
  signal reg_q1161        : std_logic;
  signal reg_q1161_in     : std_logic;
  		

  -- state q1918
  signal reg_q1918        : std_logic;
  signal reg_q1918_in     : std_logic;
  		

  -- state q1766
  signal reg_q1766        : std_logic;
  signal reg_q1766_in     : std_logic;
  		

  -- state q1715
  signal reg_q1715        : std_logic;
  signal reg_q1715_in     : std_logic;
  		

  -- state q530
  signal reg_q530        : std_logic;
  signal reg_q530_in     : std_logic;
  		

  -- state q32
  signal reg_q32        : std_logic;
  signal reg_q32_in     : std_logic;
  		

  -- state q34
  signal reg_q34        : std_logic;
  signal reg_q34_in     : std_logic;
  		

  -- state q990
  signal reg_q990        : std_logic;
  signal reg_q990_in     : std_logic;
  		

  -- state q992
  signal reg_q992        : std_logic;
  signal reg_q992_in     : std_logic;
  		

  -- state q18
  signal reg_q18        : std_logic;
  signal reg_q18_in     : std_logic;
  		

  -- state q20
  signal reg_q20        : std_logic;
  signal reg_q20_in     : std_logic;
  		

  -- state q9
  signal reg_q9        : std_logic;
  signal reg_q9_in     : std_logic;
  		

  -- state q11
  signal reg_q11        : std_logic;
  signal reg_q11_in     : std_logic;
  		

  -- state q1735
  signal reg_q1735        : std_logic;
  signal reg_q1735_in     : std_logic;
  		

  -- state q1737
  signal reg_q1737        : std_logic;
  signal reg_q1737_in     : std_logic;
  		

  -- state q1331
  signal reg_q1331        : std_logic;
  signal reg_q1331_in     : std_logic;
  		

  -- state q1333
  signal reg_q1333        : std_logic;
  signal reg_q1333_in     : std_logic;
  		

  -- state q1713
  signal reg_q1713        : std_logic;
  signal reg_q1713_in     : std_logic;
  		

  -- state q373
  signal reg_q373        : std_logic;
  signal reg_q373_in     : std_logic;
  		

  -- state q375
  signal reg_q375        : std_logic;
  signal reg_q375_in     : std_logic;
  		

  -- state q2395
  signal reg_q2395        : std_logic;
  signal reg_q2395_in     : std_logic;
  		

  -- state q2397
  signal reg_q2397        : std_logic;
  signal reg_q2397_in     : std_logic;
  		

  -- state q2601
  signal reg_q2601        : std_logic;
  signal reg_q2601_in     : std_logic;
  		

  -- state q77
  signal reg_q77        : std_logic;
  signal reg_q77_in     : std_logic;
  		

  -- state q2694
  signal reg_q2694        : std_logic;
  signal reg_q2694_in     : std_logic;
  		

  -- state q2696
  signal reg_q2696        : std_logic;
  signal reg_q2696_in     : std_logic;
  		

  -- state q2310
  signal reg_q2310        : std_logic;
  signal reg_q2310_in     : std_logic;
  		

  -- state q1012
  signal reg_q1012        : std_logic;
  signal reg_q1012_in     : std_logic;
  		

  -- state q1014
  signal reg_q1014        : std_logic;
  signal reg_q1014_in     : std_logic;
  		

  -- state q1193
  signal reg_q1193        : std_logic;
  signal reg_q1193_in     : std_logic;
  		

  -- state q1195
  signal reg_q1195        : std_logic;
  signal reg_q1195_in     : std_logic;
  		

  -- state q2407
  signal reg_q2407        : std_logic;
  signal reg_q2407_in     : std_logic;
  		

  -- state q2409
  signal reg_q2409        : std_logic;
  signal reg_q2409_in     : std_logic;
  		

  -- state q2718
  signal reg_q2718        : std_logic;
  signal reg_q2718_in     : std_logic;
  		

  -- state q2720
  signal reg_q2720        : std_logic;
  signal reg_q2720_in     : std_logic;
  		

  -- state q216
  signal reg_q216        : std_logic;
  signal reg_q216_in     : std_logic;
  		

  -- state q1327
  signal reg_q1327        : std_logic;
  signal reg_q1327_in     : std_logic;
  		

  -- state q551
  signal reg_q551        : std_logic;
  signal reg_q551_in     : std_logic;
  		

  -- state q2048
  signal reg_q2048        : std_logic;
  signal reg_q2048_in     : std_logic;
  		

  -- state q105
  signal reg_q105        : std_logic;
  signal reg_q105_in     : std_logic;
  		

  -- state q1484
  signal reg_q1484        : std_logic;
  signal reg_q1484_in     : std_logic;
  		

  -- state q250
  signal reg_q250        : std_logic;
  signal reg_q250_in     : std_logic;
  		

  -- state q252
  signal reg_q252        : std_logic;
  signal reg_q252_in     : std_logic;
  		

  -- state q2415
  signal reg_q2415        : std_logic;
  signal reg_q2415_in     : std_logic;
  		

  -- state q2010
  signal reg_q2010        : std_logic;
  signal reg_q2010_in     : std_logic;
  		

  -- state q2585
  signal reg_q2585        : std_logic;
  signal reg_q2585_in     : std_logic;
  		

  -- state q2682
  signal reg_q2682        : std_logic;
  signal reg_q2682_in     : std_logic;
  		

  -- state q996
  signal reg_q996        : std_logic;
  signal reg_q996_in     : std_logic;
  		

  -- state q998
  signal reg_q998        : std_logic;
  signal reg_q998_in     : std_logic;
  		

  -- state q1808
  signal reg_q1808        : std_logic;
  signal reg_q1808_in     : std_logic;
  		

  -- state q1810
  signal reg_q1810        : std_logic;
  signal reg_q1810_in     : std_logic;
  		

  -- state q1725
  signal reg_q1725        : std_logic;
  signal reg_q1725_in     : std_logic;
  		

  -- state q1727
  signal reg_q1727        : std_logic;
  signal reg_q1727_in     : std_logic;
  		

  -- state q1743
  signal reg_q1743        : std_logic;
  signal reg_q1743_in     : std_logic;
  		

  -- state q1745
  signal reg_q1745        : std_logic;
  signal reg_q1745_in     : std_logic;
  		

  -- state q204
  signal reg_q204        : std_logic;
  signal reg_q204_in     : std_logic;
  		

  -- state q206
  signal reg_q206        : std_logic;
  signal reg_q206_in     : std_logic;
  		

  -- state q2393
  signal reg_q2393        : std_logic;
  signal reg_q2393_in     : std_logic;
  		

  -- state q1762
  signal reg_q1762        : std_logic;
  signal reg_q1762_in     : std_logic;
  		

  -- state q1764
  signal reg_q1764        : std_logic;
  signal reg_q1764_in     : std_logic;
  		

  -- state q868
  signal reg_q868        : std_logic;
  signal reg_q868_in     : std_logic;
  		

  -- state q2684
  signal reg_q2684        : std_logic;
  signal reg_q2684_in     : std_logic;
  		

  -- state q2686
  signal reg_q2686        : std_logic;
  signal reg_q2686_in     : std_logic;
  		

  -- state q746
  signal reg_q746        : std_logic;
  signal reg_q746_in     : std_logic;
  		

  -- state q87
  signal reg_q87        : std_logic;
  signal reg_q87_in     : std_logic;
  		

  -- state q89
  signal reg_q89        : std_logic;
  signal reg_q89_in     : std_logic;
  		

  -- state q5
  signal reg_q5        : std_logic;
  signal reg_q5_in     : std_logic;
  		

  -- state q1165
  signal reg_q1165        : std_logic;
  signal reg_q1165_in     : std_logic;
  		

  -- state q1167
  signal reg_q1167        : std_logic;
  signal reg_q1167_in     : std_logic;
  		

  -- state q1208
  signal reg_q1208        : std_logic;
  signal reg_q1208_in     : std_logic;
  		

  -- state q1210
  signal reg_q1210        : std_logic;
  signal reg_q1210_in     : std_logic;
  		

  -- state q254
  signal reg_q254        : std_logic;
  signal reg_q254_in     : std_logic;
  		

  -- state q1313
  signal reg_q1313        : std_logic;
  signal reg_q1313_in     : std_logic;
  		

  -- state q1132
  signal reg_q1132        : std_logic;
  signal reg_q1132_in     : std_logic;
  		

  -- state q2308
  signal reg_q2308        : std_logic;
  signal reg_q2308_in     : std_logic;
  		

  -- state q702
  signal reg_q702        : std_logic;
  signal reg_q702_in     : std_logic;
  		

  -- state q1081
  signal reg_q1081        : std_logic;
  signal reg_q1081_in     : std_logic;
  		

  -- state q988
  signal reg_q988        : std_logic;
  signal reg_q988_in     : std_logic;
  		

  -- state q1689
  signal reg_q1689        : std_logic;
  signal reg_q1689_in     : std_logic;
  		

  -- state q1691
  signal reg_q1691        : std_logic;
  signal reg_q1691_in     : std_logic;
  		

  -- state q2615
  signal reg_q2615        : std_logic;
  signal reg_q2615_in     : std_logic;
  		

  -- state q1514
  signal reg_q1514        : std_logic;
  signal reg_q1514_in     : std_logic;
  		

  -- state q1516
  signal reg_q1516        : std_logic;
  signal reg_q1516_in     : std_logic;
  		

  -- state q740
  signal reg_q740        : std_logic;
  signal reg_q740_in     : std_logic;
  		

  -- state q563
  signal reg_q563        : std_logic;
  signal reg_q563_in     : std_logic;
  		

  -- state q994
  signal reg_q994        : std_logic;
  signal reg_q994_in     : std_logic;
  		

  -- state q2002
  signal reg_q2002        : std_logic;
  signal reg_q2002_in     : std_logic;
  		

  -- state q708
  signal reg_q708        : std_logic;
  signal reg_q708_in     : std_logic;
  		

  -- state q710
  signal reg_q710        : std_logic;
  signal reg_q710_in     : std_logic;
  		

  -- state q1185
  signal reg_q1185        : std_logic;
  signal reg_q1185_in     : std_logic;
  		

  -- state q2357
  signal reg_q2357        : std_logic;
  signal reg_q2357_in     : std_logic;
  		

  -- state q2359
  signal reg_q2359        : std_logic;
  signal reg_q2359_in     : std_logic;
  		

  -- state q226
  signal reg_q226        : std_logic;
  signal reg_q226_in     : std_logic;
  		

  -- state q228
  signal reg_q228        : std_logic;
  signal reg_q228_in     : std_logic;
  		

  -- state q1339
  signal reg_q1339        : std_logic;
  signal reg_q1339_in     : std_logic;
  		

  -- state q1341
  signal reg_q1341        : std_logic;
  signal reg_q1341_in     : std_logic;
  		

  -- state q1124
  signal reg_q1124        : std_logic;
  signal reg_q1124_in     : std_logic;
  		

  -- state q1317
  signal reg_q1317        : std_logic;
  signal reg_q1317_in     : std_logic;
  		

  -- state q38
  signal reg_q38        : std_logic;
  signal reg_q38_in     : std_logic;
  		

  -- state q673
  signal reg_q673        : std_logic;
  signal reg_q673_in     : std_logic;
  		

  -- state q1349
  signal reg_q1349        : std_logic;
  signal reg_q1349_in     : std_logic;
  		

  -- state q1351
  signal reg_q1351        : std_logic;
  signal reg_q1351_in     : std_logic;
  		

  -- state q1494
  signal reg_q1494        : std_logic;
  signal reg_q1494_in     : std_logic;
  		

  -- state q1496
  signal reg_q1496        : std_logic;
  signal reg_q1496_in     : std_logic;
  		

  -- state q532
  signal reg_q532        : std_logic;
  signal reg_q532_in     : std_logic;
  		

  -- state q534
  signal reg_q534        : std_logic;
  signal reg_q534_in     : std_logic;
  		

  -- state q967
  signal reg_q967        : std_logic;
  signal reg_q967_in     : std_logic;
  		

  -- state q955
  signal reg_q955        : std_logic;
  signal reg_q955_in     : std_logic;
  		

  -- state q270
  signal reg_q270        : std_logic;
  signal reg_q270_in     : std_logic;
  		

  -- state q272
  signal reg_q272        : std_logic;
  signal reg_q272_in     : std_logic;
  		

  -- state q734
  signal reg_q734        : std_logic;
  signal reg_q734_in     : std_logic;
  		

  -- state q736
  signal reg_q736        : std_logic;
  signal reg_q736_in     : std_logic;
  		

  -- state q1004
  signal reg_q1004        : std_logic;
  signal reg_q1004_in     : std_logic;
  		

  -- state q1006
  signal reg_q1006        : std_logic;
  signal reg_q1006_in     : std_logic;
  		

  -- state q1077
  signal reg_q1077        : std_logic;
  signal reg_q1077_in     : std_logic;
  		

  -- state q1079
  signal reg_q1079        : std_logic;
  signal reg_q1079_in     : std_logic;
  		

  -- state q2268
  signal reg_q2268        : std_logic;
  signal reg_q2268_in     : std_logic;
  		

  -- state q2270
  signal reg_q2270        : std_logic;
  signal reg_q2270_in     : std_logic;
  		

  -- state q2298
  signal reg_q2298        : std_logic;
  signal reg_q2298_in     : std_logic;
  		

  -- state q2300
  signal reg_q2300        : std_logic;
  signal reg_q2300_in     : std_logic;
  		

  -- state q1905
  signal reg_q1905        : std_logic;
  signal reg_q1905_in     : std_logic;
  		

  -- state q1163
  signal reg_q1163        : std_logic;
  signal reg_q1163_in     : std_logic;
  		

  -- state q1812
  signal reg_q1812        : std_logic;
  signal reg_q1812_in     : std_logic;
  		

  -- state q1814
  signal reg_q1814        : std_logic;
  signal reg_q1814_in     : std_logic;
  		

  -- state q1000
  signal reg_q1000        : std_logic;
  signal reg_q1000_in     : std_logic;
  		

  -- state q1069
  signal reg_q1069        : std_logic;
  signal reg_q1069_in     : std_logic;
  		

  -- state q274
  signal reg_q274        : std_logic;
  signal reg_q274_in     : std_logic;
  		

  -- state q1794
  signal reg_q1794        : std_logic;
  signal reg_q1794_in     : std_logic;
  		

  -- state q1796
  signal reg_q1796        : std_logic;
  signal reg_q1796_in     : std_logic;
  		

  -- state q280
  signal reg_q280        : std_logic;
  signal reg_q280_in     : std_logic;
  		

  -- state q2347
  signal reg_q2347        : std_logic;
  signal reg_q2347_in     : std_logic;
  		

  -- state q2349
  signal reg_q2349        : std_logic;
  signal reg_q2349_in     : std_logic;
  		

  -- state q387
  signal reg_q387        : std_logic;
  signal reg_q387_in     : std_logic;
  		

  -- state q389
  signal reg_q389        : std_logic;
  signal reg_q389_in     : std_logic;
  		

  -- state q1343
  signal reg_q1343        : std_logic;
  signal reg_q1343_in     : std_logic;
  		

  -- state q1729
  signal reg_q1729        : std_logic;
  signal reg_q1729_in     : std_logic;
  		

  -- state q2522
  signal reg_q2522        : std_logic;
  signal reg_q2522_in     : std_logic;
  		

  -- state q2722
  signal reg_q2722        : std_logic;
  signal reg_q2722_in     : std_logic;
  		

  -- state q2724
  signal reg_q2724        : std_logic;
  signal reg_q2724_in     : std_logic;
  		

  -- state q1776
  signal reg_q1776        : std_logic;
  signal reg_q1776_in     : std_logic;
  		

  -- state q2286
  signal reg_q2286        : std_logic;
  signal reg_q2286_in     : std_logic;
  		

  -- state q264
  signal reg_q264        : std_logic;
  signal reg_q264_in     : std_logic;
  		

  -- state q2373
  signal reg_q2373        : std_logic;
  signal reg_q2373_in     : std_logic;
  		

  -- state q2375
  signal reg_q2375        : std_logic;
  signal reg_q2375_in     : std_logic;
  		

  -- state q2702
  signal reg_q2702        : std_logic;
  signal reg_q2702_in     : std_logic;
  		

  -- state q276
  signal reg_q276        : std_logic;
  signal reg_q276_in     : std_logic;
  		

  -- state q278
  signal reg_q278        : std_logic;
  signal reg_q278_in     : std_logic;
  		

  -- state q383
  signal reg_q383        : std_logic;
  signal reg_q383_in     : std_logic;
  		

  -- state q385
  signal reg_q385        : std_logic;
  signal reg_q385_in     : std_logic;
  		

  -- state q679
  signal reg_q679        : std_logic;
  signal reg_q679_in     : std_logic;
  		

  -- state q2284
  signal reg_q2284        : std_logic;
  signal reg_q2284_in     : std_logic;
  		

  -- state q1008
  signal reg_q1008        : std_logic;
  signal reg_q1008_in     : std_logic;
  		

  -- state q83
  signal reg_q83        : std_logic;
  signal reg_q83_in     : std_logic;
  		

  -- state q85
  signal reg_q85        : std_logic;
  signal reg_q85_in     : std_logic;
  		

  -- state q1181
  signal reg_q1181        : std_logic;
  signal reg_q1181_in     : std_logic;
  		

  -- state q1345
  signal reg_q1345        : std_logic;
  signal reg_q1345_in     : std_logic;
  		

  -- state q730
  signal reg_q730        : std_logic;
  signal reg_q730_in     : std_logic;
  		

  -- state q2341
  signal reg_q2341        : std_logic;
  signal reg_q2341_in     : std_logic;
  		

  -- state q2343
  signal reg_q2343        : std_logic;
  signal reg_q2343_in     : std_logic;
  		

  -- state q669
  signal reg_q669        : std_logic;
  signal reg_q669_in     : std_logic;
  		

  -- state q1518
  signal reg_q1518        : std_logic;
  signal reg_q1518_in     : std_logic;
  		

  -- state q1112
  signal reg_q1112        : std_logic;
  signal reg_q1112_in     : std_logic;
  		

  -- state q1114
  signal reg_q1114        : std_logic;
  signal reg_q1114_in     : std_logic;
  		

  -- state q230
  signal reg_q230        : std_logic;
  signal reg_q230_in     : std_logic;
  		

  -- state q1118
  signal reg_q1118        : std_logic;
  signal reg_q1118_in     : std_logic;
  		

  -- state q1120
  signal reg_q1120        : std_logic;
  signal reg_q1120_in     : std_logic;
  		

  -- state q14
  signal reg_q14        : std_logic;
  signal reg_q14_in     : std_logic;
  		

  -- state q16
  signal reg_q16        : std_logic;
  signal reg_q16_in     : std_logic;
  		

  -- state q1071
  signal reg_q1071        : std_logic;
  signal reg_q1071_in     : std_logic;
  		

  -- state q2256
  signal reg_q2256        : std_logic;
  signal reg_q2256_in     : std_logic;
  		

  -- state q2258
  signal reg_q2258        : std_logic;
  signal reg_q2258_in     : std_logic;
  		

  -- state q1335
  signal reg_q1335        : std_logic;
  signal reg_q1335_in     : std_logic;
  		

  -- state q681
  signal reg_q681        : std_logic;
  signal reg_q681_in     : std_logic;
  		

  -- state q683
  signal reg_q683        : std_logic;
  signal reg_q683_in     : std_logic;
  		

  -- state q1984
  signal reg_q1984        : std_logic;
  signal reg_q1984_in     : std_logic;
  		

  -- state q1986
  signal reg_q1986        : std_logic;
  signal reg_q1986_in     : std_logic;
  		

  -- state q26
  signal reg_q26        : std_logic;
  signal reg_q26_in     : std_logic;
  		

  -- state q28
  signal reg_q28        : std_logic;
  signal reg_q28_in     : std_logic;
  		

  -- state q22
  signal reg_q22        : std_logic;
  signal reg_q22_in     : std_logic;
  		

  -- state q1699
  signal reg_q1699        : std_logic;
  signal reg_q1699_in     : std_logic;
  		

  -- state q1175
  signal reg_q1175        : std_logic;
  signal reg_q1175_in     : std_logic;
  		

  -- state q1177
  signal reg_q1177        : std_logic;
  signal reg_q1177_in     : std_logic;
  		

  -- state q381
  signal reg_q381        : std_logic;
  signal reg_q381_in     : std_logic;
  		

  -- state q2365
  signal reg_q2365        : std_logic;
  signal reg_q2365_in     : std_logic;
  		

  -- state q2367
  signal reg_q2367        : std_logic;
  signal reg_q2367_in     : std_logic;
  		

  -- state q192
  signal reg_q192        : std_logic;
  signal reg_q192_in     : std_logic;
  		

  -- state q194
  signal reg_q194        : std_logic;
  signal reg_q194_in     : std_logic;
  		

  -- state q1488
  signal reg_q1488        : std_logic;
  signal reg_q1488_in     : std_logic;
  		

  -- state q1490
  signal reg_q1490        : std_logic;
  signal reg_q1490_in     : std_logic;
  		

  -- state q1758
  signal reg_q1758        : std_logic;
  signal reg_q1758_in     : std_logic;
  		

  -- state q1760
  signal reg_q1760        : std_logic;
  signal reg_q1760_in     : std_logic;
  		

  -- state q2331
  signal reg_q2331        : std_logic;
  signal reg_q2331_in     : std_logic;
  		

  -- state q2333
  signal reg_q2333        : std_logic;
  signal reg_q2333_in     : std_logic;
  		

  -- state q163
  signal reg_q163        : std_logic;
  signal reg_q163_in     : std_logic;
  		

  -- state q165
  signal reg_q165        : std_logic;
  signal reg_q165_in     : std_logic;
  		

  -- state q2252
  signal reg_q2252        : std_logic;
  signal reg_q2252_in     : std_logic;
  		

  -- state q2254
  signal reg_q2254        : std_logic;
  signal reg_q2254_in     : std_logic;
  		

  -- state q1988
  signal reg_q1988        : std_logic;
  signal reg_q1988_in     : std_logic;
  		

  -- state q553
  signal reg_q553        : std_logic;
  signal reg_q553_in     : std_logic;
  		

  -- state q671
  signal reg_q671        : std_logic;
  signal reg_q671_in     : std_logic;
  		

  -- state q2716
  signal reg_q2716        : std_logic;
  signal reg_q2716_in     : std_logic;
  		

  -- state q2690
  signal reg_q2690        : std_logic;
  signal reg_q2690_in     : std_logic;
  		

  -- state q2692
  signal reg_q2692        : std_logic;
  signal reg_q2692_in     : std_logic;
  		

  -- state q1741
  signal reg_q1741        : std_logic;
  signal reg_q1741_in     : std_logic;
  		

  -- state q1337
  signal reg_q1337        : std_logic;
  signal reg_q1337_in     : std_logic;
  		

  -- state q75
  signal reg_q75        : std_logic;
  signal reg_q75_in     : std_logic;
  		

  -- state q24
  signal reg_q24        : std_logic;
  signal reg_q24_in     : std_logic;
  		

  -- state q1191
  signal reg_q1191        : std_logic;
  signal reg_q1191_in     : std_logic;
  		

  -- state q2603
  signal reg_q2603        : std_logic;
  signal reg_q2603_in     : std_logic;
  		

  -- state q2605
  signal reg_q2605        : std_logic;
  signal reg_q2605_in     : std_logic;
  		

  -- state q1932
  signal reg_q1932        : std_logic;
  signal reg_q1932_in     : std_logic;
  		

  -- state q950
  signal reg_q950        : std_logic;
  signal reg_q950_in     : std_logic;
  		

  -- state q2710
  signal reg_q2710        : std_logic;
  signal reg_q2710_in     : std_logic;
  		

  -- state q36
  signal reg_q36        : std_logic;
  signal reg_q36_in     : std_logic;
  		

  -- state q1155
  signal reg_q1155        : std_logic;
  signal reg_q1155_in     : std_logic;
  		

  -- state q1157
  signal reg_q1157        : std_logic;
  signal reg_q1157_in     : std_logic;
  		

  -- state q153
  signal reg_q153        : std_logic;
  signal reg_q153_in     : std_logic;
  		

  -- state q1169
  signal reg_q1169        : std_logic;
  signal reg_q1169_in     : std_logic;
  		

  -- state q266
  signal reg_q266        : std_logic;
  signal reg_q266_in     : std_logic;
  		

  -- state q507
  signal reg_q507        : std_logic;
  signal reg_q507_in     : std_logic;
  		

  -- state q509
  signal reg_q509        : std_logic;
  signal reg_q509_in     : std_logic;
  		

  -- state q2611
  signal reg_q2611        : std_logic;
  signal reg_q2611_in     : std_logic;
  		

  -- state q2613
  signal reg_q2613        : std_logic;
  signal reg_q2613_in     : std_logic;
  		

  -- state q2700
  signal reg_q2700        : std_logic;
  signal reg_q2700_in     : std_logic;
  		

  -- state q196
  signal reg_q196        : std_logic;
  signal reg_q196_in     : std_logic;
  		

  -- state q2708
  signal reg_q2708        : std_logic;
  signal reg_q2708_in     : std_logic;
  		

  -- state q561
  signal reg_q561        : std_logic;
  signal reg_q561_in     : std_logic;
  		

  -- state q161
  signal reg_q161        : std_logic;
  signal reg_q161_in     : std_logic;
  		

  -- state q224
  signal reg_q224        : std_logic;
  signal reg_q224_in     : std_logic;
  		

  -- state q232
  signal reg_q232        : std_logic;
  signal reg_q232_in     : std_logic;
  		

  -- state q234
  signal reg_q234        : std_logic;
  signal reg_q234_in     : std_logic;
  		

  -- state q2593
  signal reg_q2593        : std_logic;
  signal reg_q2593_in     : std_logic;
  		

  -- state q2595
  signal reg_q2595        : std_logic;
  signal reg_q2595_in     : std_logic;
  		

  -- state q594
  signal reg_q594        : std_logic;
  signal reg_q594_in     : std_logic;
  		

  -- state q2698
  signal reg_q2698        : std_logic;
  signal reg_q2698_in     : std_logic;
  		

  -- state q67
  signal reg_q67        : std_logic;
  signal reg_q67_in     : std_logic;
  		

  -- state q2302
  signal reg_q2302        : std_logic;
  signal reg_q2302_in     : std_logic;
  		

  -- state q2351
  signal reg_q2351        : std_logic;
  signal reg_q2351_in     : std_logic;
  		

  -- state q2353
  signal reg_q2353        : std_logic;
  signal reg_q2353_in     : std_logic;
  		

  -- state q1930
  signal reg_q1930        : std_logic;
  signal reg_q1930_in     : std_logic;
  		

  -- state q1695
  signal reg_q1695        : std_logic;
  signal reg_q1695_in     : std_logic;
  		

  -- state q1697
  signal reg_q1697        : std_logic;
  signal reg_q1697_in     : std_logic;
  		

  -- state q268
  signal reg_q268        : std_logic;
  signal reg_q268_in     : std_logic;
  		

  -- state q1085
  signal reg_q1085        : std_logic;
  signal reg_q1085_in     : std_logic;
  		

  -- state q685
  signal reg_q685        : std_logic;
  signal reg_q685_in     : std_logic;
  		

  -- state q1739
  signal reg_q1739        : std_logic;
  signal reg_q1739_in     : std_logic;
  		

  -- state q2361
  signal reg_q2361        : std_logic;
  signal reg_q2361_in     : std_logic;
  		

  -- state q262
  signal reg_q262        : std_logic;
  signal reg_q262_in     : std_logic;
  		

  -- state q46
  signal reg_q46        : std_logic;
  signal reg_q46_in     : std_logic;
  		

  -- state q1747
  signal reg_q1747        : std_logic;
  signal reg_q1747_in     : std_logic;
  		

  -- state q2371
  signal reg_q2371        : std_logic;
  signal reg_q2371_in     : std_logic;
  		

  -- state q2324
  signal reg_q2324        : std_logic;
  signal reg_q2324_in     : std_logic;
  		

  -- state q1980
  signal reg_q1980        : std_logic;
  signal reg_q1980_in     : std_logic;
  		

  -- state q2379
  signal reg_q2379        : std_logic;
  signal reg_q2379_in     : std_logic;
  		

  -- state q139
  signal reg_q139        : std_logic;
  signal reg_q139_in     : std_logic;
  		

  -- state q2377
  signal reg_q2377        : std_logic;
  signal reg_q2377_in     : std_logic;
  		

  -- state q93
  signal reg_q93        : std_logic;
  signal reg_q93_in     : std_logic;
  		

  -- state q95
  signal reg_q95        : std_logic;
  signal reg_q95_in     : std_logic;
  		

  -- state q1798
  signal reg_q1798        : std_logic;
  signal reg_q1798_in     : std_logic;
  		

  -- state q2730
  signal reg_q2730        : std_logic;
  signal reg_q2730_in     : std_logic;
  		

  -- state q2732
  signal reg_q2732        : std_logic;
  signal reg_q2732_in     : std_logic;
  		

  -- state q1329
  signal reg_q1329        : std_logic;
  signal reg_q1329_in     : std_logic;
  		

  -- state q155
  signal reg_q155        : std_logic;
  signal reg_q155_in     : std_logic;
  		

  -- state q157
  signal reg_q157        : std_logic;
  signal reg_q157_in     : std_logic;
  		

  -- state q1784
  signal reg_q1784        : std_logic;
  signal reg_q1784_in     : std_logic;
  		

  -- state q202
  signal reg_q202        : std_logic;
  signal reg_q202_in     : std_logic;
  		

  -- state q1002
  signal reg_q1002        : std_logic;
  signal reg_q1002_in     : std_logic;
  		

  -- state q2335
  signal reg_q2335        : std_logic;
  signal reg_q2335_in     : std_logic;
  		

  -- state q1792
  signal reg_q1792        : std_logic;
  signal reg_q1792_in     : std_logic;
  		

  -- state q1134
  signal reg_q1134        : std_logic;
  signal reg_q1134_in     : std_logic;
  		

  -- state q677
  signal reg_q677        : std_logic;
  signal reg_q677_in     : std_logic;
  		

  -- state q2734
  signal reg_q2734        : std_logic;
  signal reg_q2734_in     : std_logic;
  		

  -- state q2322
  signal reg_q2322        : std_logic;
  signal reg_q2322_in     : std_logic;
  		

  -- state q1140
  signal reg_q1140        : std_logic;
  signal reg_q1140_in     : std_logic;
  		

  -- state q2403
  signal reg_q2403        : std_logic;
  signal reg_q2403_in     : std_logic;
  		

  -- state q2405
  signal reg_q2405        : std_logic;
  signal reg_q2405_in     : std_logic;
  		

  -- state q2320
  signal reg_q2320        : std_logic;
  signal reg_q2320_in     : std_logic;
  		

  -- state q1153
  signal reg_q1153        : std_logic;
  signal reg_q1153_in     : std_logic;
  		

  -- state q505
  signal reg_q505        : std_logic;
  signal reg_q505_in     : std_logic;
  		

  -- state q1687
  signal reg_q1687        : std_logic;
  signal reg_q1687_in     : std_logic;
  		

  -- state q65
  signal reg_q65        : std_logic;
  signal reg_q65_in     : std_logic;
  		

  -- state q56
  signal reg_q56        : std_logic;
  signal reg_q56_in     : std_logic;
  		

  -- state q687
  signal reg_q687        : std_logic;
  signal reg_q687_in     : std_logic;
  		

  -- state q365
  signal reg_q365        : std_logic;
  signal reg_q365_in     : std_logic;
  		

  -- state q367
  signal reg_q367        : std_logic;
  signal reg_q367_in     : std_logic;
  		

  -- state q2260
  signal reg_q2260        : std_logic;
  signal reg_q2260_in     : std_logic;
  		

  -- state q2262
  signal reg_q2262        : std_logic;
  signal reg_q2262_in     : std_logic;
  		

  -- state q363
  signal reg_q363        : std_logic;
  signal reg_q363_in     : std_logic;
  		

  -- state q1104
  signal reg_q1104        : std_logic;
  signal reg_q1104_in     : std_logic;
  		

  -- state q1106
  signal reg_q1106        : std_logic;
  signal reg_q1106_in     : std_logic;
  		

  -- state q728
  signal reg_q728        : std_logic;
  signal reg_q728_in     : std_logic;
  		

  -- state q957
  signal reg_q957        : std_logic;
  signal reg_q957_in     : std_logic;
  		

  -- state q1506
  signal reg_q1506        : std_logic;
  signal reg_q1506_in     : std_logic;
  		

  -- state q137
  signal reg_q137        : std_logic;
  signal reg_q137_in     : std_logic;
  		

  -- state q2337
  signal reg_q2337        : std_logic;
  signal reg_q2337_in     : std_logic;
  		

  -- state q2339
  signal reg_q2339        : std_logic;
  signal reg_q2339_in     : std_logic;
  		

  -- state q986
  signal reg_q986        : std_logic;
  signal reg_q986_in     : std_logic;
  		

  -- state q738
  signal reg_q738        : std_logic;
  signal reg_q738_in     : std_logic;
  		

  -- state q1116
  signal reg_q1116        : std_logic;
  signal reg_q1116_in     : std_logic;
  		

  -- state q91
  signal reg_q91        : std_logic;
  signal reg_q91_in     : std_logic;
  		

  -- state q1179
  signal reg_q1179        : std_logic;
  signal reg_q1179_in     : std_logic;
  		

  -- state q1693
  signal reg_q1693        : std_logic;
  signal reg_q1693_in     : std_logic;
  		

  -- state q2391
  signal reg_q2391        : std_logic;
  signal reg_q2391_in     : std_logic;
  		

  -- state q2607
  signal reg_q2607        : std_logic;
  signal reg_q2607_in     : std_logic;
  		

  -- state q2609
  signal reg_q2609        : std_logic;
  signal reg_q2609_in     : std_logic;
  		

  -- state q1087
  signal reg_q1087        : std_logic;
  signal reg_q1087_in     : std_logic;
  		

  -- state q1786
  signal reg_q1786        : std_logic;
  signal reg_q1786_in     : std_logic;
  		

  -- state q1788
  signal reg_q1788        : std_logic;
  signal reg_q1788_in     : std_logic;
  		

  -- state q1016
  signal reg_q1016        : std_logic;
  signal reg_q1016_in     : std_logic;
  		

  -- state q706
  signal reg_q706        : std_logic;
  signal reg_q706_in     : std_logic;
  		

  -- state q2355
  signal reg_q2355        : std_logic;
  signal reg_q2355_in     : std_logic;
  		

  -- state q2688
  signal reg_q2688        : std_logic;
  signal reg_q2688_in     : std_logic;
  		

  -- state q222
  signal reg_q222        : std_logic;
  signal reg_q222_in     : std_logic;
  		

  -- state q248
  signal reg_q248        : std_logic;
  signal reg_q248_in     : std_logic;
  		

  -- state q1353
  signal reg_q1353        : std_logic;
  signal reg_q1353_in     : std_logic;
  		

  -- state q63
  signal reg_q63        : std_logic;
  signal reg_q63_in     : std_logic;
  		

  -- state q984
  signal reg_q984        : std_logic;
  signal reg_q984_in     : std_logic;
  		

  -- state q2748
  signal reg_q2748        : std_logic;
  signal reg_q2748_in     : std_logic;
  		

  -- state q1018
  signal reg_q1018        : std_logic;
  signal reg_q1018_in     : std_logic;
  		

  -- state q2411
  signal reg_q2411        : std_logic;
  signal reg_q2411_in     : std_logic;
  		

  -- state q2589
  signal reg_q2589        : std_logic;
  signal reg_q2589_in     : std_logic;
  		

  -- state q2591
  signal reg_q2591        : std_logic;
  signal reg_q2591_in     : std_logic;
  		

  -- state q1982
  signal reg_q1982        : std_logic;
  signal reg_q1982_in     : std_logic;
  		

  -- state q2401
  signal reg_q2401        : std_logic;
  signal reg_q2401_in     : std_logic;
  		

  -- state q1319
  signal reg_q1319        : std_logic;
  signal reg_q1319_in     : std_logic;
  		

  -- state q726
  signal reg_q726        : std_logic;
  signal reg_q726_in     : std_logic;
  		

  -- state q1108
  signal reg_q1108        : std_logic;
  signal reg_q1108_in     : std_logic;
  		

  -- state q1110
  signal reg_q1110        : std_logic;
  signal reg_q1110_in     : std_logic;
  		

  -- state q1355
  signal reg_q1355        : std_logic;
  signal reg_q1355_in     : std_logic;
  		

  -- state q704
  signal reg_q704        : std_logic;
  signal reg_q704_in     : std_logic;
  		

  -- state q1122
  signal reg_q1122        : std_logic;
  signal reg_q1122_in     : std_logic;
  		

  -- state q1749
  signal reg_q1749        : std_logic;
  signal reg_q1749_in     : std_logic;
  		

  -- state q159
  signal reg_q159        : std_logic;
  signal reg_q159_in     : std_logic;
  		

  -- state q2587
  signal reg_q2587        : std_logic;
  signal reg_q2587_in     : std_logic;
  		

  -- state q2345
  signal reg_q2345        : std_logic;
  signal reg_q2345_in     : std_logic;
  		

  -- state q2750
  signal reg_q2750        : std_logic;
  signal reg_q2750_in     : std_logic;
  		

  -- state q1937
  signal reg_q1937        : std_logic;
  signal reg_q1937_in     : std_logic;
  		

  -- state q1705
  signal reg_q1705        : std_logic;
  signal reg_q1705_in     : std_logic;
  		

  -- state q748
  signal reg_q748        : std_logic;
  signal reg_q748_in     : std_logic;
  		

  -- state q2369
  signal reg_q2369        : std_logic;
  signal reg_q2369_in     : std_logic;
  		

  -- state q596
  signal reg_q596        : std_logic;
  signal reg_q596_in     : std_logic;
  		

  -- state q598
  signal reg_q598        : std_logic;
  signal reg_q598_in     : std_logic;
  		

  -- state q1321
  signal reg_q1321        : std_logic;
  signal reg_q1321_in     : std_logic;
  		

  -- state q2318
  signal reg_q2318        : std_logic;
  signal reg_q2318_in     : std_logic;
  		

  -- state q976
  signal reg_q976        : std_logic;
  signal reg_q976_in     : std_logic;
  		

  -- state q1782
  signal reg_q1782        : std_logic;
  signal reg_q1782_in     : std_logic;
  		

  -- state q7
  signal reg_q7        : std_logic;
  signal reg_q7_in     : std_logic;
  		

  -- state q2248
  signal reg_q2248        : std_logic;
  signal reg_q2248_in     : std_logic;
  		

  -- state q103
  signal reg_q103        : std_logic;
  signal reg_q103_in     : std_logic;
  		

  -- state q513
  signal reg_q513        : std_logic;
  signal reg_q513_in     : std_logic;
  		

  -- state q980
  signal reg_q980        : std_logic;
  signal reg_q980_in     : std_logic;
  		

  -- state q982
  signal reg_q982        : std_logic;
  signal reg_q982_in     : std_logic;
  		

  -- state q246
  signal reg_q246        : std_logic;
  signal reg_q246_in     : std_logic;
  		

  -- state q965
  signal reg_q965        : std_logic;
  signal reg_q965_in     : std_logic;
  		

  -- state q1508
  signal reg_q1508        : std_logic;
  signal reg_q1508_in     : std_logic;
  		

  -- state q1067
  signal reg_q1067        : std_logic;
  signal reg_q1067_in     : std_logic;
  		

  -- state q48
  signal reg_q48        : std_logic;
  signal reg_q48_in     : std_logic;
  		

  -- state q1347
  signal reg_q1347        : std_logic;
  signal reg_q1347_in     : std_logic;
  		

  -- state q1091
  signal reg_q1091        : std_logic;
  signal reg_q1091_in     : std_logic;
  		

  -- state q1093
  signal reg_q1093        : std_logic;
  signal reg_q1093_in     : std_logic;
  		

  -- state q1751
  signal reg_q1751        : std_logic;
  signal reg_q1751_in     : std_logic;
  		

  -- state q1790
  signal reg_q1790        : std_logic;
  signal reg_q1790_in     : std_logic;
  		

  -- state q750
  signal reg_q750        : std_logic;
  signal reg_q750_in     : std_logic;
  		

  -- state q1492
  signal reg_q1492        : std_logic;
  signal reg_q1492_in     : std_logic;
  		

  -- state q1928
  signal reg_q1928        : std_logic;
  signal reg_q1928_in     : std_logic;
  		

  -- state q1089
  signal reg_q1089        : std_logic;
  signal reg_q1089_in     : std_logic;
  		

  -- state q1197
  signal reg_q1197        : std_logic;
  signal reg_q1197_in     : std_logic;
  		

  -- state q600
  signal reg_q600        : std_logic;
  signal reg_q600_in     : std_logic;
  		

  -- state q602
  signal reg_q602        : std_logic;
  signal reg_q602_in     : std_logic;
  		

  -- state q536
  signal reg_q536        : std_logic;
  signal reg_q536_in     : std_logic;
  		

  -- state q538
  signal reg_q538        : std_logic;
  signal reg_q538_in     : std_logic;
  		

  -- state q2250
  signal reg_q2250        : std_logic;
  signal reg_q2250_in     : std_logic;
  		

  -- state q73
  signal reg_q73        : std_logic;
  signal reg_q73_in     : std_logic;
  		

  -- state q978
  signal reg_q978        : std_logic;
  signal reg_q978_in     : std_logic;
  		

  -- state q256
  signal reg_q256        : std_logic;
  signal reg_q256_in     : std_logic;
  		

  -- state q128
  signal reg_q128        : std_logic;
  signal reg_q128_in     : std_logic;
  		

  -- state q130
  signal reg_q130        : std_logic;
  signal reg_q130_in     : std_logic;
  		

  -- state q959
  signal reg_q959        : std_logic;
  signal reg_q959_in     : std_logic;
  		

  -- state q960
  signal reg_q960        : std_logic;
  signal reg_q960_in     : std_logic;
  		

  -- state q2413
  signal reg_q2413        : std_logic;
  signal reg_q2413_in     : std_logic;
  		

  -- state q752
  signal reg_q752        : std_logic;
  signal reg_q752_in     : std_logic;
  		

  -- state q1216
  signal reg_q1216        : std_logic;
  signal reg_q1216_in     : std_logic;
  		

  -- state q198
  signal reg_q198        : std_logic;
  signal reg_q198_in     : std_logic;
  		

  -- state q1142
  signal reg_q1142        : std_logic;
  signal reg_q1142_in     : std_logic;
  		

  -- state q2755
  signal reg_q2755        : std_logic;
  signal reg_q2755_in     : std_logic;
  		

  -- state q689
  signal reg_q689        : std_logic;
  signal reg_q689_in     : std_logic;
  		

  -- state q97
  signal reg_q97        : std_logic;
  signal reg_q97_in     : std_logic;
  		

  -- state q754
  signal reg_q754        : std_logic;
  signal reg_q754_in     : std_logic;
  		

  -- state q1753
  signal reg_q1753        : std_logic;
  signal reg_q1753_in     : std_logic;
  		

  -- state q691
  signal reg_q691        : std_logic;
  signal reg_q691_in     : std_logic;
  		

  -- state q200
  signal reg_q200        : std_logic;
  signal reg_q200_in     : std_logic;
  		

  -- state q1020
  signal reg_q1020        : std_logic;
  signal reg_q1020_in     : std_logic;
  		
  signal reg_fullgraph1       : std_logic_vector(9 downto 0);
  signal reg_fullgraph1_in    : std_logic_vector(9 downto 0);
  signal reg_fullgraph1_init  : std_logic_vector(9 downto 0);
  signal reg_fullgraph1_sel   : std_logic_vector(1023 downto 0); 	
  -- end section fullgraph1
  --#################################################			
		

  -- state q772
  signal reg_q772        : std_logic;
  signal reg_q772_in     : std_logic;
  signal reg_q772_init   : std_logic;
		

  -- state q590
  signal reg_q590        : std_logic;
  signal reg_q590_in     : std_logic;
  signal reg_q590_init   : std_logic;
		

  -- state q545
  signal reg_q545        : std_logic;
  signal reg_q545_in     : std_logic;
  signal reg_q545_init   : std_logic;
		
--#################################################
-- start section fullgraph: 5

  -- state q2231
  signal reg_q2231        : std_logic;
  signal reg_q2231_in     : std_logic;
  		

  -- state q2233
  signal reg_q2233        : std_logic;
  signal reg_q2233_in     : std_logic;
  		

  -- state q1961
  signal reg_q1961        : std_logic;
  signal reg_q1961_in     : std_logic;
  		

  -- state q1672
  signal reg_q1672        : std_logic;
  signal reg_q1672_in     : std_logic;
  		

  -- state q2429
  signal reg_q2429        : std_logic;
  signal reg_q2429_in     : std_logic;
  		

  -- state q1602
  signal reg_q1602        : std_logic;
  signal reg_q1602_in     : std_logic;
  		

  -- state q1604
  signal reg_q1604        : std_logic;
  signal reg_q1604_in     : std_logic;
  		

  -- state q308
  signal reg_q308        : std_logic;
  signal reg_q308_in     : std_logic;
  		

  -- state q2651
  signal reg_q2651        : std_logic;
  signal reg_q2651_in     : std_logic;
  		

  -- state q1443
  signal reg_q1443        : std_logic;
  signal reg_q1443_in     : std_logic;
  		

  -- state q644
  signal reg_q644        : std_logic;
  signal reg_q644_in     : std_logic;
  		

  -- state q646
  signal reg_q646        : std_logic;
  signal reg_q646_in     : std_logic;
  		

  -- state q179
  signal reg_q179        : std_logic;
  signal reg_q179_in     : std_logic;
  		

  -- state q634
  signal reg_q634        : std_logic;
  signal reg_q634_in     : std_logic;
  		

  -- state q636
  signal reg_q636        : std_logic;
  signal reg_q636_in     : std_logic;
  		

  -- state q2570
  signal reg_q2570        : std_logic;
  signal reg_q2570_in     : std_logic;
  		

  -- state q2572
  signal reg_q2572        : std_logic;
  signal reg_q2572_in     : std_logic;
  		

  -- state q2451
  signal reg_q2451        : std_logic;
  signal reg_q2451_in     : std_logic;
  		

  -- state q2453
  signal reg_q2453        : std_logic;
  signal reg_q2453_in     : std_logic;
  		

  -- state q819
  signal reg_q819        : std_logic;
  signal reg_q819_in     : std_logic;
  		

  -- state q1377
  signal reg_q1377        : std_logic;
  signal reg_q1377_in     : std_logic;
  		

  -- state q1379
  signal reg_q1379        : std_logic;
  signal reg_q1379_in     : std_logic;
  		

  -- state q2534
  signal reg_q2534        : std_logic;
  signal reg_q2534_in     : std_logic;
  		

  -- state q1890
  signal reg_q1890        : std_logic;
  signal reg_q1890_in     : std_logic;
  		

  -- state q1892
  signal reg_q1892        : std_logic;
  signal reg_q1892_in     : std_logic;
  		

  -- state q2082
  signal reg_q2082        : std_logic;
  signal reg_q2082_in     : std_logic;
  		

  -- state q2627
  signal reg_q2627        : std_logic;
  signal reg_q2627_in     : std_logic;
  		

  -- state q2150
  signal reg_q2150        : std_logic;
  signal reg_q2150_in     : std_logic;
  		

  -- state q316
  signal reg_q316        : std_logic;
  signal reg_q316_in     : std_logic;
  		

  -- state q318
  signal reg_q318        : std_logic;
  signal reg_q318_in     : std_logic;
  		

  -- state q620
  signal reg_q620        : std_logic;
  signal reg_q620_in     : std_logic;
  		

  -- state q622
  signal reg_q622        : std_logic;
  signal reg_q622_in     : std_logic;
  		

  -- state q1616
  signal reg_q1616        : std_logic;
  signal reg_q1616_in     : std_logic;
  		

  -- state q2112
  signal reg_q2112        : std_logic;
  signal reg_q2112_in     : std_logic;
  		

  -- state q2439
  signal reg_q2439        : std_logic;
  signal reg_q2439_in     : std_logic;
  		

  -- state q2441
  signal reg_q2441        : std_logic;
  signal reg_q2441_in     : std_logic;
  		

  -- state q2192
  signal reg_q2192        : std_logic;
  signal reg_q2192_in     : std_logic;
  		

  -- state q2194
  signal reg_q2194        : std_logic;
  signal reg_q2194_in     : std_logic;
  		

  -- state q1524
  signal reg_q1524        : std_logic;
  signal reg_q1524_in     : std_logic;
  		

  -- state q2092
  signal reg_q2092        : std_logic;
  signal reg_q2092_in     : std_logic;
  		

  -- state q2094
  signal reg_q2094        : std_logic;
  signal reg_q2094_in     : std_logic;
  		

  -- state q439
  signal reg_q439        : std_logic;
  signal reg_q439_in     : std_logic;
  		

  -- state q441
  signal reg_q441        : std_logic;
  signal reg_q441_in     : std_logic;
  		

  -- state q488
  signal reg_q488        : std_logic;
  signal reg_q488_in     : std_logic;
  		

  -- state q490
  signal reg_q490        : std_logic;
  signal reg_q490_in     : std_logic;
  		

  -- state q173
  signal reg_q173        : std_logic;
  signal reg_q173_in     : std_logic;
  		

  -- state q2576
  signal reg_q2576        : std_logic;
  signal reg_q2576_in     : std_logic;
  		

  -- state q2578
  signal reg_q2578        : std_logic;
  signal reg_q2578_in     : std_logic;
  		

  -- state q1042
  signal reg_q1042        : std_logic;
  signal reg_q1042_in     : std_logic;
  		

  -- state q1044
  signal reg_q1044        : std_logic;
  signal reg_q1044_in     : std_logic;
  		

  -- state q2235
  signal reg_q2235        : std_logic;
  signal reg_q2235_in     : std_logic;
  		

  -- state q608
  signal reg_q608        : std_logic;
  signal reg_q608_in     : std_logic;
  		

  -- state q1658
  signal reg_q1658        : std_logic;
  signal reg_q1658_in     : std_logic;
  		

  -- state q1660
  signal reg_q1660        : std_logic;
  signal reg_q1660_in     : std_logic;
  		

  -- state q792
  signal reg_q792        : std_logic;
  signal reg_q792_in     : std_logic;
  		

  -- state q794
  signal reg_q794        : std_logic;
  signal reg_q794_in     : std_logic;
  		

  -- state q1606
  signal reg_q1606        : std_logic;
  signal reg_q1606_in     : std_logic;
  		

  -- state q312
  signal reg_q312        : std_logic;
  signal reg_q312_in     : std_logic;
  		

  -- state q314
  signal reg_q314        : std_logic;
  signal reg_q314_in     : std_logic;
  		

  -- state q2479
  signal reg_q2479        : std_logic;
  signal reg_q2479_in     : std_logic;
  		

  -- state q1526
  signal reg_q1526        : std_logic;
  signal reg_q1526_in     : std_logic;
  		

  -- state q1528
  signal reg_q1528        : std_logic;
  signal reg_q1528_in     : std_logic;
  		

  -- state q1844
  signal reg_q1844        : std_logic;
  signal reg_q1844_in     : std_logic;
  		

  -- state q890
  signal reg_q890        : std_logic;
  signal reg_q890_in     : std_logic;
  		

  -- state q892
  signal reg_q892        : std_logic;
  signal reg_q892_in     : std_logic;
  		

  -- state q183
  signal reg_q183        : std_logic;
  signal reg_q183_in     : std_logic;
  		

  -- state q2509
  signal reg_q2509        : std_logic;
  signal reg_q2509_in     : std_logic;
  		

  -- state q2511
  signal reg_q2511        : std_logic;
  signal reg_q2511_in     : std_logic;
  		

  -- state q1858
  signal reg_q1858        : std_logic;
  signal reg_q1858_in     : std_logic;
  		

  -- state q1860
  signal reg_q1860        : std_logic;
  signal reg_q1860_in     : std_logic;
  		

  -- state q290
  signal reg_q290        : std_logic;
  signal reg_q290_in     : std_logic;
  		

  -- state q292
  signal reg_q292        : std_logic;
  signal reg_q292_in     : std_logic;
  		

  -- state q2437
  signal reg_q2437        : std_logic;
  signal reg_q2437_in     : std_logic;
  		

  -- state q1473
  signal reg_q1473        : std_logic;
  signal reg_q1473_in     : std_logic;
  		

  -- state q1475
  signal reg_q1475        : std_logic;
  signal reg_q1475_in     : std_logic;
  		

  -- state q1260
  signal reg_q1260        : std_logic;
  signal reg_q1260_in     : std_logic;
  		

  -- state q1262
  signal reg_q1262        : std_logic;
  signal reg_q1262_in     : std_logic;
  		

  -- state q575
  signal reg_q575        : std_logic;
  signal reg_q575_in     : std_logic;
  		

  -- state q1427
  signal reg_q1427        : std_logic;
  signal reg_q1427_in     : std_logic;
  		

  -- state q1429
  signal reg_q1429        : std_logic;
  signal reg_q1429_in     : std_logic;
  		

  -- state q904
  signal reg_q904        : std_logic;
  signal reg_q904_in     : std_logic;
  		

  -- state q906
  signal reg_q906        : std_logic;
  signal reg_q906_in     : std_logic;
  		

  -- state q862
  signal reg_q862        : std_logic;
  signal reg_q862_in     : std_logic;
  		

  -- state q1832
  signal reg_q1832        : std_logic;
  signal reg_q1832_in     : std_logic;
  		

  -- state q1834
  signal reg_q1834        : std_logic;
  signal reg_q1834_in     : std_logic;
  		

  -- state q1610
  signal reg_q1610        : std_logic;
  signal reg_q1610_in     : std_logic;
  		

  -- state q1612
  signal reg_q1612        : std_logic;
  signal reg_q1612_in     : std_logic;
  		

  -- state q767
  signal reg_q767        : std_logic;
  signal reg_q767_in     : std_logic;
  		

  -- state q1546
  signal reg_q1546        : std_logic;
  signal reg_q1546_in     : std_logic;
  		

  -- state q1548
  signal reg_q1548        : std_logic;
  signal reg_q1548_in     : std_logic;
  		

  -- state q1854
  signal reg_q1854        : std_logic;
  signal reg_q1854_in     : std_logic;
  		

  -- state q1856
  signal reg_q1856        : std_logic;
  signal reg_q1856_in     : std_logic;
  		

  -- state q437
  signal reg_q437        : std_logic;
  signal reg_q437_in     : std_logic;
  		

  -- state q328
  signal reg_q328        : std_logic;
  signal reg_q328_in     : std_logic;
  		

  -- state q330
  signal reg_q330        : std_logic;
  signal reg_q330_in     : std_logic;
  		

  -- state q2190
  signal reg_q2190        : std_logic;
  signal reg_q2190_in     : std_logic;
  		

  -- state q1600
  signal reg_q1600        : std_logic;
  signal reg_q1600_in     : std_logic;
  		

  -- state q2560
  signal reg_q2560        : std_logic;
  signal reg_q2560_in     : std_logic;
  		

  -- state q2562
  signal reg_q2562        : std_logic;
  signal reg_q2562_in     : std_logic;
  		

  -- state q2168
  signal reg_q2168        : std_logic;
  signal reg_q2168_in     : std_logic;
  		

  -- state q2170
  signal reg_q2170        : std_logic;
  signal reg_q2170_in     : std_logic;
  		

  -- state q583
  signal reg_q583        : std_logic;
  signal reg_q583_in     : std_logic;
  		

  -- state q2568
  signal reg_q2568        : std_logic;
  signal reg_q2568_in     : std_logic;
  		

  -- state q1431
  signal reg_q1431        : std_logic;
  signal reg_q1431_in     : std_logic;
  		

  -- state q419
  signal reg_q419        : std_logic;
  signal reg_q419_in     : std_logic;
  		

  -- state q415
  signal reg_q415        : std_logic;
  signal reg_q415_in     : std_logic;
  		

  -- state q417
  signal reg_q417        : std_logic;
  signal reg_q417_in     : std_logic;
  		

  -- state q1266
  signal reg_q1266        : std_logic;
  signal reg_q1266_in     : std_logic;
  		

  -- state q2108
  signal reg_q2108        : std_logic;
  signal reg_q2108_in     : std_logic;
  		

  -- state q2110
  signal reg_q2110        : std_logic;
  signal reg_q2110_in     : std_logic;
  		

  -- state q1371
  signal reg_q1371        : std_logic;
  signal reg_q1371_in     : std_logic;
  		

  -- state q1373
  signal reg_q1373        : std_logic;
  signal reg_q1373_in     : std_logic;
  		

  -- state q786
  signal reg_q786        : std_logic;
  signal reg_q786_in     : std_logic;
  		

  -- state q2659
  signal reg_q2659        : std_logic;
  signal reg_q2659_in     : std_logic;
  		

  -- state q2661
  signal reg_q2661        : std_logic;
  signal reg_q2661_in     : std_logic;
  		

  -- state q1274
  signal reg_q1274        : std_logic;
  signal reg_q1274_in     : std_logic;
  		

  -- state q1276
  signal reg_q1276        : std_logic;
  signal reg_q1276_in     : std_logic;
  		

  -- state q2493
  signal reg_q2493        : std_logic;
  signal reg_q2493_in     : std_logic;
  		

  -- state q1375
  signal reg_q1375        : std_logic;
  signal reg_q1375_in     : std_logic;
  		

  -- state q1405
  signal reg_q1405        : std_logic;
  signal reg_q1405_in     : std_logic;
  		

  -- state q1407
  signal reg_q1407        : std_logic;
  signal reg_q1407_in     : std_logic;
  		

  -- state q916
  signal reg_q916        : std_logic;
  signal reg_q916_in     : std_logic;
  		

  -- state q918
  signal reg_q918        : std_logic;
  signal reg_q918_in     : std_logic;
  		

  -- state q2467
  signal reg_q2467        : std_logic;
  signal reg_q2467_in     : std_logic;
  		

  -- state q2469
  signal reg_q2469        : std_logic;
  signal reg_q2469_in     : std_logic;
  		

  -- state q1943
  signal reg_q1943        : std_logic;
  signal reg_q1943_in     : std_logic;
  		

  -- state q1232
  signal reg_q1232        : std_logic;
  signal reg_q1232_in     : std_logic;
  		

  -- state q1234
  signal reg_q1234        : std_logic;
  signal reg_q1234_in     : std_logic;
  		

  -- state q1477
  signal reg_q1477        : std_logic;
  signal reg_q1477_in     : std_logic;
  		

  -- state q1230
  signal reg_q1230        : std_logic;
  signal reg_q1230_in     : std_logic;
  		

  -- state q1250
  signal reg_q1250        : std_logic;
  signal reg_q1250_in     : std_logic;
  		

  -- state q1252
  signal reg_q1252        : std_logic;
  signal reg_q1252_in     : std_logic;
  		

  -- state q1423
  signal reg_q1423        : std_logic;
  signal reg_q1423_in     : std_logic;
  		

  -- state q1425
  signal reg_q1425        : std_logic;
  signal reg_q1425_in     : std_logic;
  		

  -- state q2212
  signal reg_q2212        : std_logic;
  signal reg_q2212_in     : std_logic;
  		

  -- state q2214
  signal reg_q2214        : std_logic;
  signal reg_q2214_in     : std_logic;
  		

  -- state q1288
  signal reg_q1288        : std_logic;
  signal reg_q1288_in     : std_logic;
  		

  -- state q1290
  signal reg_q1290        : std_logic;
  signal reg_q1290_in     : std_logic;
  		

  -- state q340
  signal reg_q340        : std_logic;
  signal reg_q340_in     : std_logic;
  		

  -- state q1622
  signal reg_q1622        : std_logic;
  signal reg_q1622_in     : std_logic;
  		

  -- state q624
  signal reg_q624        : std_logic;
  signal reg_q624_in     : std_logic;
  		

  -- state q423
  signal reg_q423        : std_logic;
  signal reg_q423_in     : std_logic;
  		

  -- state q425
  signal reg_q425        : std_logic;
  signal reg_q425_in     : std_logic;
  		

  -- state q1588
  signal reg_q1588        : std_logic;
  signal reg_q1588_in     : std_logic;
  		

  -- state q1590
  signal reg_q1590        : std_logic;
  signal reg_q1590_in     : std_logic;
  		

  -- state q332
  signal reg_q332        : std_logic;
  signal reg_q332_in     : std_logic;
  		

  -- state q2076
  signal reg_q2076        : std_logic;
  signal reg_q2076_in     : std_logic;
  		

  -- state q2078
  signal reg_q2078        : std_logic;
  signal reg_q2078_in     : std_logic;
  		

  -- state q1248
  signal reg_q1248        : std_logic;
  signal reg_q1248_in     : std_logic;
  		

  -- state q181
  signal reg_q181        : std_logic;
  signal reg_q181_in     : std_logic;
  		

  -- state q585
  signal reg_q585        : std_logic;
  signal reg_q585_in     : std_logic;
  		

  -- state q334
  signal reg_q334        : std_logic;
  signal reg_q334_in     : std_logic;
  		

  -- state q2124
  signal reg_q2124        : std_logic;
  signal reg_q2124_in     : std_logic;
  		

  -- state q2126
  signal reg_q2126        : std_logic;
  signal reg_q2126_in     : std_logic;
  		

  -- state q2558
  signal reg_q2558        : std_logic;
  signal reg_q2558_in     : std_logic;
  		

  -- state q1449
  signal reg_q1449        : std_logic;
  signal reg_q1449_in     : std_logic;
  		

  -- state q1451
  signal reg_q1451        : std_logic;
  signal reg_q1451_in     : std_logic;
  		

  -- state q835
  signal reg_q835        : std_logic;
  signal reg_q835_in     : std_logic;
  		

  -- state q837
  signal reg_q837        : std_logic;
  signal reg_q837_in     : std_logic;
  		

  -- state q626
  signal reg_q626        : std_logic;
  signal reg_q626_in     : std_logic;
  		

  -- state q628
  signal reg_q628        : std_logic;
  signal reg_q628_in     : std_logic;
  		

  -- state q1258
  signal reg_q1258        : std_logic;
  signal reg_q1258_in     : std_logic;
  		

  -- state q1558
  signal reg_q1558        : std_logic;
  signal reg_q1558_in     : std_logic;
  		

  -- state q1668
  signal reg_q1668        : std_logic;
  signal reg_q1668_in     : std_logic;
  		

  -- state q1670
  signal reg_q1670        : std_logic;
  signal reg_q1670_in     : std_logic;
  		

  -- state q1570
  signal reg_q1570        : std_logic;
  signal reg_q1570_in     : std_logic;
  		

  -- state q1572
  signal reg_q1572        : std_logic;
  signal reg_q1572_in     : std_logic;
  		

  -- state q1580
  signal reg_q1580        : std_logic;
  signal reg_q1580_in     : std_logic;
  		

  -- state q1582
  signal reg_q1582        : std_logic;
  signal reg_q1582_in     : std_logic;
  		

  -- state q841
  signal reg_q841        : std_logic;
  signal reg_q841_in     : std_logic;
  		

  -- state q652
  signal reg_q652        : std_logic;
  signal reg_q652_in     : std_logic;
  		

  -- state q654
  signal reg_q654        : std_logic;
  signal reg_q654_in     : std_logic;
  		

  -- state q1409
  signal reg_q1409        : std_logic;
  signal reg_q1409_in     : std_logic;
  		

  -- state q839
  signal reg_q839        : std_logic;
  signal reg_q839_in     : std_logic;
  		

  -- state q1421
  signal reg_q1421        : std_logic;
  signal reg_q1421_in     : std_logic;
  		

  -- state q912
  signal reg_q912        : std_logic;
  signal reg_q912_in     : std_logic;
  		

  -- state q1272
  signal reg_q1272        : std_logic;
  signal reg_q1272_in     : std_logic;
  		

  -- state q1614
  signal reg_q1614        : std_logic;
  signal reg_q1614_in     : std_logic;
  		

  -- state q2530
  signal reg_q2530        : std_logic;
  signal reg_q2530_in     : std_logic;
  		

  -- state q2532
  signal reg_q2532        : std_logic;
  signal reg_q2532_in     : std_logic;
  		

  -- state q928
  signal reg_q928        : std_logic;
  signal reg_q928_in     : std_logic;
  		

  -- state q930
  signal reg_q930        : std_logic;
  signal reg_q930_in     : std_logic;
  		

  -- state q2198
  signal reg_q2198        : std_logic;
  signal reg_q2198_in     : std_logic;
  		

  -- state q2200
  signal reg_q2200        : std_logic;
  signal reg_q2200_in     : std_logic;
  		

  -- state q503
  signal reg_q503        : std_logic;
  signal reg_q503_in     : std_logic;
  		

  -- state q2146
  signal reg_q2146        : std_logic;
  signal reg_q2146_in     : std_logic;
  		

  -- state q2148
  signal reg_q2148        : std_logic;
  signal reg_q2148_in     : std_logic;
  		

  -- state q926
  signal reg_q926        : std_logic;
  signal reg_q926_in     : std_logic;
  		

  -- state q1325
  signal reg_q1325        : std_logic;
  signal reg_q1325_in     : std_logic;
  		

  -- state q549
  signal reg_q549        : std_logic;
  signal reg_q549_in     : std_logic;
  		

  -- state q403
  signal reg_q403        : std_logic;
  signal reg_q403_in     : std_logic;
  		

  -- state q2188
  signal reg_q2188        : std_logic;
  signal reg_q2188_in     : std_logic;
  		

  -- state q898
  signal reg_q898        : std_logic;
  signal reg_q898_in     : std_logic;
  		

  -- state q900
  signal reg_q900        : std_logic;
  signal reg_q900_in     : std_logic;
  		

  -- state q630
  signal reg_q630        : std_logic;
  signal reg_q630_in     : std_logic;
  		

  -- state q632
  signal reg_q632        : std_logic;
  signal reg_q632_in     : std_logic;
  		

  -- state q1455
  signal reg_q1455        : std_logic;
  signal reg_q1455_in     : std_logic;
  		

  -- state q1254
  signal reg_q1254        : std_logic;
  signal reg_q1254_in     : std_logic;
  		

  -- state q1256
  signal reg_q1256        : std_logic;
  signal reg_q1256_in     : std_logic;
  		

  -- state q1138
  signal reg_q1138        : std_logic;
  signal reg_q1138_in     : std_logic;
  		

  -- state q1278
  signal reg_q1278        : std_logic;
  signal reg_q1278_in     : std_logic;
  		

  -- state q1280
  signal reg_q1280        : std_logic;
  signal reg_q1280_in     : std_logic;
  		

  -- state q656
  signal reg_q656        : std_logic;
  signal reg_q656_in     : std_logic;
  		

  -- state q2540
  signal reg_q2540        : std_logic;
  signal reg_q2540_in     : std_logic;
  		

  -- state q2542
  signal reg_q2542        : std_logic;
  signal reg_q2542_in     : std_logic;
  		

  -- state q910
  signal reg_q910        : std_logic;
  signal reg_q910_in     : std_logic;
  		

  -- state q2176
  signal reg_q2176        : std_logic;
  signal reg_q2176_in     : std_logic;
  		

  -- state q2178
  signal reg_q2178        : std_logic;
  signal reg_q2178_in     : std_logic;
  		

  -- state q2070
  signal reg_q2070        : std_logic;
  signal reg_q2070_in     : std_logic;
  		

  -- state q2072
  signal reg_q2072        : std_logic;
  signal reg_q2072_in     : std_logic;
  		

  -- state q1242
  signal reg_q1242        : std_logic;
  signal reg_q1242_in     : std_logic;
  		

  -- state q1244
  signal reg_q1244        : std_logic;
  signal reg_q1244_in     : std_logic;
  		

  -- state q2156
  signal reg_q2156        : std_logic;
  signal reg_q2156_in     : std_logic;
  		

  -- state q2158
  signal reg_q2158        : std_logic;
  signal reg_q2158_in     : std_logic;
  		

  -- state q2465
  signal reg_q2465        : std_logic;
  signal reg_q2465_in     : std_logic;
  		

  -- state q924
  signal reg_q924        : std_logic;
  signal reg_q924_in     : std_logic;
  		

  -- state q2088
  signal reg_q2088        : std_logic;
  signal reg_q2088_in     : std_logic;
  		

  -- state q2090
  signal reg_q2090        : std_logic;
  signal reg_q2090_in     : std_logic;
  		

  -- state q2066
  signal reg_q2066        : std_logic;
  signal reg_q2066_in     : std_logic;
  		

  -- state q870
  signal reg_q870        : std_logic;
  signal reg_q870_in     : std_logic;
  		

  -- state q2184
  signal reg_q2184        : std_logic;
  signal reg_q2184_in     : std_logic;
  		

  -- state q2186
  signal reg_q2186        : std_logic;
  signal reg_q2186_in     : std_logic;
  		

  -- state q864
  signal reg_q864        : std_logic;
  signal reg_q864_in     : std_logic;
  		

  -- state q866
  signal reg_q866        : std_logic;
  signal reg_q866_in     : std_logic;
  		

  -- state q2497
  signal reg_q2497        : std_logic;
  signal reg_q2497_in     : std_logic;
  		

  -- state q433
  signal reg_q433        : std_logic;
  signal reg_q433_in     : std_logic;
  		

  -- state q1822
  signal reg_q1822        : std_logic;
  signal reg_q1822_in     : std_logic;
  		

  -- state q1662
  signal reg_q1662        : std_logic;
  signal reg_q1662_in     : std_logic;
  		

  -- state q2120
  signal reg_q2120        : std_logic;
  signal reg_q2120_in     : std_logic;
  		

  -- state q1236
  signal reg_q1236        : std_logic;
  signal reg_q1236_in     : std_logic;
  		

  -- state q1036
  signal reg_q1036        : std_logic;
  signal reg_q1036_in     : std_logic;
  		

  -- state q1538
  signal reg_q1538        : std_logic;
  signal reg_q1538_in     : std_logic;
  		

  -- state q1540
  signal reg_q1540        : std_logic;
  signal reg_q1540_in     : std_logic;
  		

  -- state q1550
  signal reg_q1550        : std_logic;
  signal reg_q1550_in     : std_logic;
  		

  -- state q1552
  signal reg_q1552        : std_logic;
  signal reg_q1552_in     : std_logic;
  		

  -- state q742
  signal reg_q742        : std_logic;
  signal reg_q742_in     : std_logic;
  		

  -- state q2671
  signal reg_q2671        : std_logic;
  signal reg_q2671_in     : std_logic;
  		

  -- state q1284
  signal reg_q1284        : std_logic;
  signal reg_q1284_in     : std_logic;
  		

  -- state q1286
  signal reg_q1286        : std_logic;
  signal reg_q1286_in     : std_logic;
  		

  -- state q1850
  signal reg_q1850        : std_logic;
  signal reg_q1850_in     : std_logic;
  		

  -- state q1852
  signal reg_q1852        : std_logic;
  signal reg_q1852_in     : std_logic;
  		

  -- state q1731
  signal reg_q1731        : std_logic;
  signal reg_q1731_in     : std_logic;
  		

  -- state q1733
  signal reg_q1733        : std_logic;
  signal reg_q1733_in     : std_logic;
  		

  -- state q612
  signal reg_q612        : std_logic;
  signal reg_q612_in     : std_logic;
  		

  -- state q614
  signal reg_q614        : std_logic;
  signal reg_q614_in     : std_logic;
  		

  -- state q825
  signal reg_q825        : std_logic;
  signal reg_q825_in     : std_logic;
  		

  -- state q2206
  signal reg_q2206        : std_logic;
  signal reg_q2206_in     : std_logic;
  		

  -- state q2208
  signal reg_q2208        : std_logic;
  signal reg_q2208_in     : std_logic;
  		

  -- state q1648
  signal reg_q1648        : std_logic;
  signal reg_q1648_in     : std_logic;
  		

  -- state q1650
  signal reg_q1650        : std_logic;
  signal reg_q1650_in     : std_logic;
  		

  -- state q1401
  signal reg_q1401        : std_logic;
  signal reg_q1401_in     : std_logic;
  		

  -- state q1888
  signal reg_q1888        : std_logic;
  signal reg_q1888_in     : std_logic;
  		

  -- state q2471
  signal reg_q2471        : std_logic;
  signal reg_q2471_in     : std_logic;
  		

  -- state q2473
  signal reg_q2473        : std_logic;
  signal reg_q2473_in     : std_logic;
  		

  -- state q326
  signal reg_q326        : std_logic;
  signal reg_q326_in     : std_logic;
  		

  -- state q1471
  signal reg_q1471        : std_logic;
  signal reg_q1471_in     : std_logic;
  		

  -- state q1246
  signal reg_q1246        : std_logic;
  signal reg_q1246_in     : std_logic;
  		

  -- state q2742
  signal reg_q2742        : std_logic;
  signal reg_q2742_in     : std_logic;
  		

  -- state q2421
  signal reg_q2421        : std_logic;
  signal reg_q2421_in     : std_logic;
  		

  -- state q2423
  signal reg_q2423        : std_logic;
  signal reg_q2423_in     : std_logic;
  		

  -- state q579
  signal reg_q579        : std_logic;
  signal reg_q579_in     : std_logic;
  		

  -- state q932
  signal reg_q932        : std_logic;
  signal reg_q932_in     : std_logic;
  		

  -- state q934
  signal reg_q934        : std_logic;
  signal reg_q934_in     : std_logic;
  		

  -- state q1907
  signal reg_q1907        : std_logic;
  signal reg_q1907_in     : std_logic;
  		

  -- state q1367
  signal reg_q1367        : std_logic;
  signal reg_q1367_in     : std_logic;
  		

  -- state q2665
  signal reg_q2665        : std_logic;
  signal reg_q2665_in     : std_logic;
  		

  -- state q2667
  signal reg_q2667        : std_logic;
  signal reg_q2667_in     : std_logic;
  		

  -- state q1638
  signal reg_q1638        : std_logic;
  signal reg_q1638_in     : std_logic;
  		

  -- state q1967
  signal reg_q1967        : std_logic;
  signal reg_q1967_in     : std_logic;
  		

  -- state q1866
  signal reg_q1866        : std_logic;
  signal reg_q1866_in     : std_logic;
  		

  -- state q1868
  signal reg_q1868        : std_logic;
  signal reg_q1868_in     : std_logic;
  		

  -- state q1304
  signal reg_q1304        : std_logic;
  signal reg_q1304_in     : std_logic;
  		

  -- state q1306
  signal reg_q1306        : std_logic;
  signal reg_q1306_in     : std_logic;
  		

  -- state q2513
  signal reg_q2513        : std_logic;
  signal reg_q2513_in     : std_logic;
  		

  -- state q1870
  signal reg_q1870        : std_logic;
  signal reg_q1870_in     : std_logic;
  		

  -- state q1872
  signal reg_q1872        : std_logic;
  signal reg_q1872_in     : std_logic;
  		

  -- state q1969
  signal reg_q1969        : std_logic;
  signal reg_q1969_in     : std_logic;
  		

  -- state q1971
  signal reg_q1971        : std_logic;
  signal reg_q1971_in     : std_logic;
  		

  -- state q577
  signal reg_q577        : std_logic;
  signal reg_q577_in     : std_logic;
  		

  -- state q413
  signal reg_q413        : std_logic;
  signal reg_q413_in     : std_logic;
  		

  -- state q405
  signal reg_q405        : std_logic;
  signal reg_q405_in     : std_logic;
  		

  -- state q407
  signal reg_q407        : std_logic;
  signal reg_q407_in     : std_logic;
  		

  -- state q2564
  signal reg_q2564        : std_logic;
  signal reg_q2564_in     : std_logic;
  		

  -- state q2740
  signal reg_q2740        : std_logic;
  signal reg_q2740_in     : std_logic;
  		

  -- state q2477
  signal reg_q2477        : std_logic;
  signal reg_q2477_in     : std_logic;
  		

  -- state q1632
  signal reg_q1632        : std_logic;
  signal reg_q1632_in     : std_logic;
  		

  -- state q306
  signal reg_q306        : std_logic;
  signal reg_q306_in     : std_logic;
  		

  -- state q2174
  signal reg_q2174        : std_logic;
  signal reg_q2174_in     : std_logic;
  		

  -- state q1282
  signal reg_q1282        : std_logic;
  signal reg_q1282_in     : std_logic;
  		

  -- state q2084
  signal reg_q2084        : std_logic;
  signal reg_q2084_in     : std_logic;
  		

  -- state q1955
  signal reg_q1955        : std_logic;
  signal reg_q1955_in     : std_logic;
  		

  -- state q1957
  signal reg_q1957        : std_logic;
  signal reg_q1957_in     : std_logic;
  		

  -- state q1238
  signal reg_q1238        : std_logic;
  signal reg_q1238_in     : std_logic;
  		

  -- state q922
  signal reg_q922        : std_logic;
  signal reg_q922_in     : std_logic;
  		

  -- state q2457
  signal reg_q2457        : std_logic;
  signal reg_q2457_in     : std_logic;
  		

  -- state q2459
  signal reg_q2459        : std_logic;
  signal reg_q2459_in     : std_logic;
  		

  -- state q463
  signal reg_q463        : std_logic;
  signal reg_q463_in     : std_logic;
  		

  -- state q465
  signal reg_q465        : std_logic;
  signal reg_q465_in     : std_logic;
  		

  -- state q320
  signal reg_q320        : std_logic;
  signal reg_q320_in     : std_logic;
  		

  -- state q322
  signal reg_q322        : std_logic;
  signal reg_q322_in     : std_logic;
  		

  -- state q2475
  signal reg_q2475        : std_logic;
  signal reg_q2475_in     : std_logic;
  		

  -- state q1901
  signal reg_q1901        : std_logic;
  signal reg_q1901_in     : std_logic;
  		

  -- state q457
  signal reg_q457        : std_logic;
  signal reg_q457_in     : std_logic;
  		

  -- state q459
  signal reg_q459        : std_logic;
  signal reg_q459_in     : std_logic;
  		

  -- state q1560
  signal reg_q1560        : std_logic;
  signal reg_q1560_in     : std_logic;
  		

  -- state q1562
  signal reg_q1562        : std_logic;
  signal reg_q1562_in     : std_logic;
  		

  -- state q336
  signal reg_q336        : std_logic;
  signal reg_q336_in     : std_logic;
  		

  -- state q338
  signal reg_q338        : std_logic;
  signal reg_q338_in     : std_logic;
  		

  -- state q300
  signal reg_q300        : std_logic;
  signal reg_q300_in     : std_logic;
  		

  -- state q573
  signal reg_q573        : std_logic;
  signal reg_q573_in     : std_logic;
  		

  -- state q765
  signal reg_q765        : std_logic;
  signal reg_q765_in     : std_logic;
  		

  -- state q1264
  signal reg_q1264        : std_logic;
  signal reg_q1264_in     : std_logic;
  		

  -- state q610
  signal reg_q610        : std_logic;
  signal reg_q610_in     : std_logic;
  		

  -- state q1512
  signal reg_q1512        : std_logic;
  signal reg_q1512_in     : std_logic;
  		

  -- state q453
  signal reg_q453        : std_logic;
  signal reg_q453_in     : std_logic;
  		

  -- state q2491
  signal reg_q2491        : std_logic;
  signal reg_q2491_in     : std_logic;
  		

  -- state q1536
  signal reg_q1536        : std_logic;
  signal reg_q1536_in     : std_logic;
  		

  -- state q2202
  signal reg_q2202        : std_logic;
  signal reg_q2202_in     : std_logic;
  		

  -- state q2204
  signal reg_q2204        : std_logic;
  signal reg_q2204_in     : std_logic;
  		

  -- state q2663
  signal reg_q2663        : std_logic;
  signal reg_q2663_in     : std_logic;
  		

  -- state q2566
  signal reg_q2566        : std_logic;
  signal reg_q2566_in     : std_logic;
  		

  -- state q2580
  signal reg_q2580        : std_logic;
  signal reg_q2580_in     : std_logic;
  		

  -- state q1959
  signal reg_q1959        : std_logic;
  signal reg_q1959_in     : std_logic;
  		

  -- state q920
  signal reg_q920        : std_logic;
  signal reg_q920_in     : std_logic;
  		

  -- state q1654
  signal reg_q1654        : std_logic;
  signal reg_q1654_in     : std_logic;
  		

  -- state q1656
  signal reg_q1656        : std_logic;
  signal reg_q1656_in     : std_logic;
  		

  -- state q1224
  signal reg_q1224        : std_logic;
  signal reg_q1224_in     : std_logic;
  		

  -- state q2106
  signal reg_q2106        : std_logic;
  signal reg_q2106_in     : std_logic;
  		

  -- state q2182
  signal reg_q2182        : std_logic;
  signal reg_q2182_in     : std_logic;
  		

  -- state q1864
  signal reg_q1864        : std_logic;
  signal reg_q1864_in     : std_logic;
  		

  -- state q1586
  signal reg_q1586        : std_logic;
  signal reg_q1586_in     : std_logic;
  		

  -- state q2455
  signal reg_q2455        : std_logic;
  signal reg_q2455_in     : std_logic;
  		

  -- state q914
  signal reg_q914        : std_logic;
  signal reg_q914_in     : std_logic;
  		

  -- state q451
  signal reg_q451        : std_logic;
  signal reg_q451_in     : std_logic;
  		

  -- state q1556
  signal reg_q1556        : std_logic;
  signal reg_q1556_in     : std_logic;
  		

  -- state q2132
  signal reg_q2132        : std_logic;
  signal reg_q2132_in     : std_logic;
  		

  -- state q2134
  signal reg_q2134        : std_logic;
  signal reg_q2134_in     : std_logic;
  		

  -- state q1417
  signal reg_q1417        : std_logic;
  signal reg_q1417_in     : std_logic;
  		

  -- state q1419
  signal reg_q1419        : std_logic;
  signal reg_q1419_in     : std_logic;
  		

  -- state q872
  signal reg_q872        : std_logic;
  signal reg_q872_in     : std_logic;
  		

  -- state q638
  signal reg_q638        : std_logic;
  signal reg_q638_in     : std_logic;
  		

  -- state q640
  signal reg_q640        : std_logic;
  signal reg_q640_in     : std_logic;
  		

  -- state q431
  signal reg_q431        : std_logic;
  signal reg_q431_in     : std_logic;
  		

  -- state q1646
  signal reg_q1646        : std_logic;
  signal reg_q1646_in     : std_logic;
  		

  -- state q1532
  signal reg_q1532        : std_logic;
  signal reg_q1532_in     : std_logic;
  		

  -- state q1624
  signal reg_q1624        : std_logic;
  signal reg_q1624_in     : std_logic;
  		

  -- state q1292
  signal reg_q1292        : std_logic;
  signal reg_q1292_in     : std_logic;
  		

  -- state q1298
  signal reg_q1298        : std_logic;
  signal reg_q1298_in     : std_logic;
  		

  -- state q2196
  signal reg_q2196        : std_logic;
  signal reg_q2196_in     : std_logic;
  		

  -- state q936
  signal reg_q936        : std_logic;
  signal reg_q936_in     : std_logic;
  		

  -- state q938
  signal reg_q938        : std_logic;
  signal reg_q938_in     : std_logic;
  		

  -- state q1083
  signal reg_q1083        : std_logic;
  signal reg_q1083_in     : std_logic;
  		

  -- state q1403
  signal reg_q1403        : std_logic;
  signal reg_q1403_in     : std_logic;
  		

  -- state q2140
  signal reg_q2140        : std_logic;
  signal reg_q2140_in     : std_logic;
  		

  -- state q2142
  signal reg_q2142        : std_logic;
  signal reg_q2142_in     : std_logic;
  		

  -- state q1886
  signal reg_q1886        : std_logic;
  signal reg_q1886_in     : std_logic;
  		

  -- state q1828
  signal reg_q1828        : std_logic;
  signal reg_q1828_in     : std_logic;
  		

  -- state q1830
  signal reg_q1830        : std_logic;
  signal reg_q1830_in     : std_logic;
  		

  -- state q2515
  signal reg_q2515        : std_logic;
  signal reg_q2515_in     : std_logic;
  		

  -- state q1381
  signal reg_q1381        : std_logic;
  signal reg_q1381_in     : std_logic;
  		

  -- state q1383
  signal reg_q1383        : std_logic;
  signal reg_q1383_in     : std_logic;
  		

  -- state q2489
  signal reg_q2489        : std_logic;
  signal reg_q2489_in     : std_logic;
  		

  -- state q650
  signal reg_q650        : std_logic;
  signal reg_q650_in     : std_logic;
  		

  -- state q744
  signal reg_q744        : std_logic;
  signal reg_q744_in     : std_logic;
  		

  -- state q1953
  signal reg_q1953        : std_logic;
  signal reg_q1953_in     : std_logic;
  		

  -- state q581
  signal reg_q581        : std_logic;
  signal reg_q581_in     : std_logic;
  		

  -- state q1542
  signal reg_q1542        : std_logic;
  signal reg_q1542_in     : std_logic;
  		

  -- state q1544
  signal reg_q1544        : std_logic;
  signal reg_q1544_in     : std_logic;
  		

  -- state q1842
  signal reg_q1842        : std_logic;
  signal reg_q1842_in     : std_logic;
  		

  -- state q2443
  signal reg_q2443        : std_logic;
  signal reg_q2443_in     : std_logic;
  		

  -- state q618
  signal reg_q618        : std_logic;
  signal reg_q618_in     : std_logic;
  		

  -- state q1413
  signal reg_q1413        : std_logic;
  signal reg_q1413_in     : std_logic;
  		

  -- state q1415
  signal reg_q1415        : std_logic;
  signal reg_q1415_in     : std_logic;
  		

  -- state q2548
  signal reg_q2548        : std_logic;
  signal reg_q2548_in     : std_logic;
  		

  -- state q1040
  signal reg_q1040        : std_logic;
  signal reg_q1040_in     : std_logic;
  		

  -- state q2096
  signal reg_q2096        : std_logic;
  signal reg_q2096_in     : std_logic;
  		

  -- state q2098
  signal reg_q2098        : std_logic;
  signal reg_q2098_in     : std_logic;
  		

  -- state q827
  signal reg_q827        : std_logic;
  signal reg_q827_in     : std_logic;
  		

  -- state q1151
  signal reg_q1151        : std_logic;
  signal reg_q1151_in     : std_logic;
  		

  -- state q2144
  signal reg_q2144        : std_logic;
  signal reg_q2144_in     : std_logic;
  		

  -- state q888
  signal reg_q888        : std_logic;
  signal reg_q888_in     : std_logic;
  		

  -- state q616
  signal reg_q616        : std_logic;
  signal reg_q616_in     : std_logic;
  		

  -- state q1608
  signal reg_q1608        : std_logic;
  signal reg_q1608_in     : std_logic;
  		

  -- state q1294
  signal reg_q1294        : std_logic;
  signal reg_q1294_in     : std_logic;
  		

  -- state q1240
  signal reg_q1240        : std_logic;
  signal reg_q1240_in     : std_logic;
  		

  -- state q658
  signal reg_q658        : std_logic;
  signal reg_q658_in     : std_logic;
  		

  -- state q886
  signal reg_q886        : std_logic;
  signal reg_q886_in     : std_logic;
  		

  -- state q1894
  signal reg_q1894        : std_logic;
  signal reg_q1894_in     : std_logic;
  		

  -- state q2445
  signal reg_q2445        : std_logic;
  signal reg_q2445_in     : std_logic;
  		

  -- state q2138
  signal reg_q2138        : std_logic;
  signal reg_q2138_in     : std_logic;
  		

  -- state q2485
  signal reg_q2485        : std_logic;
  signal reg_q2485_in     : std_logic;
  		

  -- state q1564
  signal reg_q1564        : std_logic;
  signal reg_q1564_in     : std_logic;
  		

  -- state q1566
  signal reg_q1566        : std_logic;
  signal reg_q1566_in     : std_logic;
  		

  -- state q1862
  signal reg_q1862        : std_logic;
  signal reg_q1862_in     : std_logic;
  		

  -- state q443
  signal reg_q443        : std_logic;
  signal reg_q443_in     : std_logic;
  		

  -- state q2210
  signal reg_q2210        : std_logic;
  signal reg_q2210_in     : std_logic;
  		

  -- state q447
  signal reg_q447        : std_logic;
  signal reg_q447_in     : std_logic;
  		

  -- state q449
  signal reg_q449        : std_logic;
  signal reg_q449_in     : std_logic;
  		

  -- state q1840
  signal reg_q1840        : std_logic;
  signal reg_q1840_in     : std_logic;
  		

  -- state q1824
  signal reg_q1824        : std_logic;
  signal reg_q1824_in     : std_logic;
  		

  -- state q1774
  signal reg_q1774        : std_logic;
  signal reg_q1774_in     : std_logic;
  		

  -- state q720
  signal reg_q720        : std_logic;
  signal reg_q720_in     : std_logic;
  		

  -- state q2483
  signal reg_q2483        : std_logic;
  signal reg_q2483_in     : std_logic;
  		

  -- state q2481
  signal reg_q2481        : std_logic;
  signal reg_q2481_in     : std_logic;
  		

  -- state q1568
  signal reg_q1568        : std_logic;
  signal reg_q1568_in     : std_logic;
  		

  -- state q2128
  signal reg_q2128        : std_logic;
  signal reg_q2128_in     : std_logic;
  		

  -- state q1666
  signal reg_q1666        : std_logic;
  signal reg_q1666_in     : std_logic;
  		

  -- state q2517
  signal reg_q2517        : std_logic;
  signal reg_q2517_in     : std_logic;
  		

  -- state q391
  signal reg_q391        : std_logic;
  signal reg_q391_in     : std_logic;
  		

  -- state q796
  signal reg_q796        : std_logic;
  signal reg_q796_in     : std_logic;
  		

  -- state q798
  signal reg_q798        : std_logic;
  signal reg_q798_in     : std_logic;
  		

  -- state q1878
  signal reg_q1878        : std_logic;
  signal reg_q1878_in     : std_logic;
  		

  -- state q1880
  signal reg_q1880        : std_logic;
  signal reg_q1880_in     : std_logic;
  		

  -- state q2499
  signal reg_q2499        : std_logic;
  signal reg_q2499_in     : std_logic;
  		

  -- state q2086
  signal reg_q2086        : std_logic;
  signal reg_q2086_in     : std_logic;
  		

  -- state q2180
  signal reg_q2180        : std_logic;
  signal reg_q2180_in     : std_logic;
  		

  -- state q421
  signal reg_q421        : std_logic;
  signal reg_q421_in     : std_logic;
  		

  -- state q2136
  signal reg_q2136        : std_logic;
  signal reg_q2136_in     : std_logic;
  		

  -- state q2507
  signal reg_q2507        : std_logic;
  signal reg_q2507_in     : std_logic;
  		

  -- state q2399
  signal reg_q2399        : std_logic;
  signal reg_q2399_in     : std_logic;
  		

  -- state q2501
  signal reg_q2501        : std_logic;
  signal reg_q2501_in     : std_logic;
  		

  -- state q304
  signal reg_q304        : std_logic;
  signal reg_q304_in     : std_logic;
  		

  -- state q2100
  signal reg_q2100        : std_logic;
  signal reg_q2100_in     : std_logic;
  		

  -- state q1664
  signal reg_q1664        : std_logic;
  signal reg_q1664_in     : std_logic;
  		

  -- state q896
  signal reg_q896        : std_logic;
  signal reg_q896_in     : std_logic;
  		

  -- state q2675
  signal reg_q2675        : std_logic;
  signal reg_q2675_in     : std_logic;
  		

  -- state q429
  signal reg_q429        : std_logic;
  signal reg_q429_in     : std_logic;
  		

  -- state q2657
  signal reg_q2657        : std_logic;
  signal reg_q2657_in     : std_logic;
  		

  -- state q2461
  signal reg_q2461        : std_logic;
  signal reg_q2461_in     : std_logic;
  		

  -- state q1226
  signal reg_q1226        : std_logic;
  signal reg_q1226_in     : std_logic;
  		

  -- state q1228
  signal reg_q1228        : std_logic;
  signal reg_q1228_in     : std_logic;
  		

  -- state q642
  signal reg_q642        : std_logic;
  signal reg_q642_in     : std_logic;
  		

  -- state q302
  signal reg_q302        : std_logic;
  signal reg_q302_in     : std_logic;
  		

  -- state q1939
  signal reg_q1939        : std_logic;
  signal reg_q1939_in     : std_logic;
  		

  -- state q2425
  signal reg_q2425        : std_logic;
  signal reg_q2425_in     : std_logic;
  		

  -- state q2427
  signal reg_q2427        : std_logic;
  signal reg_q2427_in     : std_logic;
  		

  -- state q1054
  signal reg_q1054        : std_logic;
  signal reg_q1054_in     : std_logic;
  		

  -- state q1056
  signal reg_q1056        : std_logic;
  signal reg_q1056_in     : std_logic;
  		

  -- state q1826
  signal reg_q1826        : std_logic;
  signal reg_q1826_in     : std_logic;
  		

  -- state q1302
  signal reg_q1302        : std_logic;
  signal reg_q1302_in     : std_logic;
  		

  -- state q1268
  signal reg_q1268        : std_logic;
  signal reg_q1268_in     : std_logic;
  		

  -- state q1874
  signal reg_q1874        : std_logic;
  signal reg_q1874_in     : std_logic;
  		

  -- state q2574
  signal reg_q2574        : std_logic;
  signal reg_q2574_in     : std_logic;
  		

  -- state q467
  signal reg_q467        : std_logic;
  signal reg_q467_in     : std_logic;
  		

  -- state q1510
  signal reg_q1510        : std_logic;
  signal reg_q1510_in     : std_logic;
  		

  -- state q1199
  signal reg_q1199        : std_logic;
  signal reg_q1199_in     : std_logic;
  		

  -- state q1201
  signal reg_q1201        : std_logic;
  signal reg_q1201_in     : std_logic;
  		

  -- state q1876
  signal reg_q1876        : std_logic;
  signal reg_q1876_in     : std_logic;
  		

  -- state q1435
  signal reg_q1435        : std_logic;
  signal reg_q1435_in     : std_logic;
  		

  -- state q1437
  signal reg_q1437        : std_logic;
  signal reg_q1437_in     : std_logic;
  		

  -- state q833
  signal reg_q833        : std_logic;
  signal reg_q833_in     : std_logic;
  		

  -- state q445
  signal reg_q445        : std_logic;
  signal reg_q445_in     : std_logic;
  		

  -- state q780
  signal reg_q780        : std_logic;
  signal reg_q780_in     : std_logic;
  		

  -- state q2463
  signal reg_q2463        : std_logic;
  signal reg_q2463_in     : std_logic;
  		

  -- state q409
  signal reg_q409        : std_logic;
  signal reg_q409_in     : std_logic;
  		

  -- state q1920
  signal reg_q1920        : std_logic;
  signal reg_q1920_in     : std_logic;
  		

  -- state q829
  signal reg_q829        : std_logic;
  signal reg_q829_in     : std_logic;
  		

  -- state q831
  signal reg_q831        : std_logic;
  signal reg_q831_in     : std_logic;
  		

  -- state q1439
  signal reg_q1439        : std_logic;
  signal reg_q1439_in     : std_logic;
  		

  -- state q1441
  signal reg_q1441        : std_logic;
  signal reg_q1441_in     : std_logic;
  		

  -- state q1678
  signal reg_q1678        : std_logic;
  signal reg_q1678_in     : std_logic;
  		

  -- state q1038
  signal reg_q1038        : std_logic;
  signal reg_q1038_in     : std_logic;
  		

  -- state q2068
  signal reg_q2068        : std_logic;
  signal reg_q2068_in     : std_logic;
  		

  -- state q1048
  signal reg_q1048        : std_logic;
  signal reg_q1048_in     : std_logic;
  		

  -- state q1050
  signal reg_q1050        : std_logic;
  signal reg_q1050_in     : std_logic;
  		

  -- state q2130
  signal reg_q2130        : std_logic;
  signal reg_q2130_in     : std_logic;
  		

  -- state q2166
  signal reg_q2166        : std_logic;
  signal reg_q2166_in     : std_logic;
  		

  -- state q324
  signal reg_q324        : std_logic;
  signal reg_q324_in     : std_logic;
  		

  -- state q1882
  signal reg_q1882        : std_logic;
  signal reg_q1882_in     : std_logic;
  		

  -- state q2669
  signal reg_q2669        : std_logic;
  signal reg_q2669_in     : std_logic;
  		

  -- state q2102
  signal reg_q2102        : std_logic;
  signal reg_q2102_in     : std_logic;
  		

  -- state q908
  signal reg_q908        : std_logic;
  signal reg_q908_in     : std_logic;
  		

  -- state q1149
  signal reg_q1149        : std_logic;
  signal reg_q1149_in     : std_logic;
  		

  -- state q2104
  signal reg_q2104        : std_logic;
  signal reg_q2104_in     : std_logic;
  		

  -- state q1838
  signal reg_q1838        : std_logic;
  signal reg_q1838_in     : std_logic;
  		

  -- state q1896
  signal reg_q1896        : std_logic;
  signal reg_q1896_in     : std_logic;
  		

  -- state q1772
  signal reg_q1772        : std_logic;
  signal reg_q1772_in     : std_logic;
  		

  -- state q1433
  signal reg_q1433        : std_logic;
  signal reg_q1433_in     : std_logic;
  		

  -- state q1554
  signal reg_q1554        : std_logic;
  signal reg_q1554_in     : std_logic;
  		

  -- state q940
  signal reg_q940        : std_logic;
  signal reg_q940_in     : std_logic;
  		

  -- state q1300
  signal reg_q1300        : std_logic;
  signal reg_q1300_in     : std_logic;
  		

  -- state q1836
  signal reg_q1836        : std_logic;
  signal reg_q1836_in     : std_logic;
  		

  -- state q2546
  signal reg_q2546        : std_logic;
  signal reg_q2546_in     : std_logic;
  		

  -- state q902
  signal reg_q902        : std_logic;
  signal reg_q902_in     : std_logic;
  		

  -- state q1680
  signal reg_q1680        : std_logic;
  signal reg_q1680_in     : std_logic;
  		

  -- state q1030
  signal reg_q1030        : std_logic;
  signal reg_q1030_in     : std_logic;
  		

  -- state q1032
  signal reg_q1032        : std_logic;
  signal reg_q1032_in     : std_logic;
  		

  -- state q1052
  signal reg_q1052        : std_logic;
  signal reg_q1052_in     : std_logic;
  		

  -- state q1898
  signal reg_q1898        : std_logic;
  signal reg_q1898_in     : std_logic;
  		

  -- state q1058
  signal reg_q1058        : std_logic;
  signal reg_q1058_in     : std_logic;
  		

  -- state q427
  signal reg_q427        : std_logic;
  signal reg_q427_in     : std_logic;
  		

  -- state q2544
  signal reg_q2544        : std_logic;
  signal reg_q2544_in     : std_logic;
  		
  signal reg_fullgraph5       : std_logic_vector(8 downto 0);
  signal reg_fullgraph5_in    : std_logic_vector(8 downto 0);
  signal reg_fullgraph5_init  : std_logic_vector(8 downto 0);
  signal reg_fullgraph5_sel   : std_logic_vector(511 downto 0); 	
  -- end section fullgraph5
  --#################################################			
		

  -- state q470
  signal reg_q470        : std_logic;
  signal reg_q470_in     : std_logic;
  signal reg_q470_init   : std_logic;
		

  -- state q694
  signal reg_q694        : std_logic;
  signal reg_q694_in     : std_logic;
  signal reg_q694_init   : std_logic;
		

  -- state q2229
  signal reg_q2229        : std_logic;
  signal reg_q2229_in     : std_logic;
  signal reg_q2229_init   : std_logic;
		

  -- state q1756
  signal reg_q1756        : std_logic;
  signal reg_q1756_in     : std_logic;
  signal reg_q1756_init   : std_logic;
		

  -- state q860
  signal reg_q860        : std_logic;
  signal reg_q860_in     : std_logic;
  signal reg_q860_init   : std_logic;
		
--#################################################
-- start section fullgraph: 11

  -- state q1975
  signal reg_q1975        : std_logic;
  signal reg_q1975_in     : std_logic;
  		

  -- state q1686
  signal reg_q1686        : std_logic;
  signal reg_q1686_in     : std_logic;
  		

  -- state q788
  signal reg_q788        : std_logic;
  signal reg_q788_in     : std_logic;
  		

  -- state q2631
  signal reg_q2631        : std_logic;
  signal reg_q2631_in     : std_logic;
  		

  -- state q518
  signal reg_q518        : std_logic;
  signal reg_q518_in     : std_logic;
  		

  -- state q474
  signal reg_q474        : std_logic;
  signal reg_q474_in     : std_logic;
  		

  -- state q1311
  signal reg_q1311        : std_logic;
  signal reg_q1311_in     : std_logic;
  		

  -- state q3
  signal reg_q3        : std_logic;
  signal reg_q3_in     : std_logic;
  		

  -- state q118
  signal reg_q118        : std_logic;
  signal reg_q118_in     : std_logic;
  		

  -- state q2246
  signal reg_q2246        : std_logic;
  signal reg_q2246_in     : std_logic;
  		

  -- state q476
  signal reg_q476        : std_logic;
  signal reg_q476_in     : std_logic;
  		

  -- state q763
  signal reg_q763        : std_logic;
  signal reg_q763_in     : std_logic;
  		

  -- state q761
  signal reg_q761        : std_logic;
  signal reg_q761_in     : std_logic;
  		

  -- state q952
  signal reg_q952        : std_logic;
  signal reg_q952_in     : std_logic;
  		

  -- state q1098
  signal reg_q1098        : std_logic;
  signal reg_q1098_in     : std_logic;
  		

  -- state q349
  signal reg_q349        : std_logic;
  signal reg_q349_in     : std_logic;
  		

  -- state q1909
  signal reg_q1909        : std_logic;
  signal reg_q1909_in     : std_logic;
  		

  -- state q1147
  signal reg_q1147        : std_logic;
  signal reg_q1147_in     : std_logic;
  		

  -- state q874
  signal reg_q874        : std_logic;
  signal reg_q874_in     : std_logic;
  		

  -- state q1486
  signal reg_q1486        : std_logic;
  signal reg_q1486_in     : std_logic;
  		

  -- state q1935
  signal reg_q1935        : std_logic;
  signal reg_q1935_in     : std_logic;
  		

  -- state q813
  signal reg_q813        : std_logic;
  signal reg_q813_in     : std_logic;
  		

  -- state q815
  signal reg_q815        : std_logic;
  signal reg_q815_in     : std_logic;
  		

  -- state q1941
  signal reg_q1941        : std_logic;
  signal reg_q1941_in     : std_logic;
  		

  -- state q353
  signal reg_q353        : std_logic;
  signal reg_q353_in     : std_logic;
  		

  -- state q351
  signal reg_q351        : std_logic;
  signal reg_q351_in     : std_logic;
  		

  -- state q1065
  signal reg_q1065        : std_logic;
  signal reg_q1065_in     : std_logic;
  		

  -- state q811
  signal reg_q811        : std_logic;
  signal reg_q811_in     : std_logic;
  		

  -- state q1903
  signal reg_q1903        : std_logic;
  signal reg_q1903_in     : std_logic;
  		

  -- state q807
  signal reg_q807        : std_logic;
  signal reg_q807_in     : std_logic;
  		

  -- state q809
  signal reg_q809        : std_logic;
  signal reg_q809_in     : std_logic;
  		

  -- state q1922
  signal reg_q1922        : std_logic;
  signal reg_q1922_in     : std_logic;
  		
  signal reg_fullgraph11       : std_logic_vector(5 downto 0);
  signal reg_fullgraph11_in    : std_logic_vector(5 downto 0);
  signal reg_fullgraph11_init  : std_logic_vector(5 downto 0);
  signal reg_fullgraph11_sel   : std_logic_vector(63 downto 0); 	
  -- end section fullgraph11
  --#################################################			
		

  -- state q286
  signal reg_q286        : std_logic;
  signal reg_q286_in     : std_logic;
  signal reg_q286_init   : std_logic;
		

  -- state q1309
  signal reg_q1309        : std_logic;
  signal reg_q1309_in     : std_logic;
  signal reg_q1309_init   : std_logic;
		

  -- state q2244
  signal reg_q2244        : std_logic;
  signal reg_q2244_in     : std_logic;
  signal reg_q2244_init   : std_logic;
		
--#################################################
-- start section fullgraph: 15

  -- state q1682
  signal reg_q1682        : std_logic;
  signal reg_q1682_in     : std_logic;
  		

  -- state q2625
  signal reg_q2625        : std_logic;
  signal reg_q2625_in     : std_logic;
  		

  -- state q499
  signal reg_q499        : std_logic;
  signal reg_q499_in     : std_logic;
  		

  -- state q663
  signal reg_q663        : std_logic;
  signal reg_q663_in     : std_logic;
  		

  -- state q520
  signal reg_q520        : std_logic;
  signal reg_q520_in     : std_logic;
  		

  -- state q667
  signal reg_q667        : std_logic;
  signal reg_q667_in     : std_logic;
  		

  -- state q101
  signal reg_q101        : std_logic;
  signal reg_q101_in     : std_logic;
  		

  -- state q1206
  signal reg_q1206        : std_logic;
  signal reg_q1206_in     : std_logic;
  		

  -- state q1978
  signal reg_q1978        : std_logic;
  signal reg_q1978_in     : std_logic;
  		

  -- state q30
  signal reg_q30        : std_logic;
  signal reg_q30_in     : std_logic;
  		

  -- state q1063
  signal reg_q1063        : std_logic;
  signal reg_q1063_in     : std_logic;
  		
  signal reg_fullgraph15       : std_logic_vector(3 downto 0);
  signal reg_fullgraph15_in    : std_logic_vector(3 downto 0);
  signal reg_fullgraph15_init  : std_logic_vector(3 downto 0);
  signal reg_fullgraph15_sel   : std_logic_vector(15 downto 0); 	
  -- end section fullgraph15
  --#################################################			
		

  -- state q945
  signal reg_q945        : std_logic;
  signal reg_q945_in     : std_logic;
  signal reg_q945_init   : std_logic;
		

  -- state q2554
  signal reg_q2554        : std_logic;
  signal reg_q2554_in     : std_logic;
  signal reg_q2554_init   : std_logic;
		

  -- state q1479
  signal reg_q1479        : std_logic;
  signal reg_q1479_in     : std_logic;
  signal reg_q1479_init   : std_logic;
		

  -- state q2583
  signal reg_q2583        : std_logic;
  signal reg_q2583_in     : std_logic;
  signal reg_q2583_init   : std_logic;
		
--#################################################
-- start section fullgraph: 20

  -- state q393
  signal reg_q393        : std_logic;
  signal reg_q393_in     : std_logic;
  		

  -- state q542
  signal reg_q542        : std_logic;
  signal reg_q542_in     : std_logic;
  		

  -- state q857
  signal reg_q857        : std_logic;
  signal reg_q857_in     : std_logic;
  		

  -- state q2629
  signal reg_q2629        : std_logic;
  signal reg_q2629_in     : std_logic;
  		

  -- state q569
  signal reg_q569        : std_logic;
  signal reg_q569_in     : std_logic;
  		

  -- state q571
  signal reg_q571        : std_logic;
  signal reg_q571_in     : std_logic;
  		

  -- state q696
  signal reg_q696        : std_logic;
  signal reg_q696_in     : std_logic;
  		

  -- state q177
  signal reg_q177        : std_logic;
  signal reg_q177_in     : std_logic;
  		

  -- state q665
  signal reg_q665        : std_logic;
  signal reg_q665_in     : std_logic;
  		

  -- state q948
  signal reg_q948        : std_logic;
  signal reg_q948_in     : std_logic;
  		

  -- state q135
  signal reg_q135        : std_logic;
  signal reg_q135_in     : std_logic;
  		
  signal reg_fullgraph20       : std_logic_vector(3 downto 0);
  signal reg_fullgraph20_in    : std_logic_vector(3 downto 0);
  signal reg_fullgraph20_init  : std_logic_vector(3 downto 0);
  signal reg_fullgraph20_sel   : std_logic_vector(15 downto 0); 	
  -- end section fullgraph20
  --#################################################			
		

  -- state q2520
  signal reg_q2520        : std_logic;
  signal reg_q2520_in     : std_logic;
  signal reg_q2520_init   : std_logic;
		
--#################################################
-- start section fullgraph: 22

  -- state q2447
  signal reg_q2447        : std_logic;
  signal reg_q2447_in     : std_logic;
  		

  -- state q773
  signal reg_q773        : std_logic;
  signal reg_q773_in     : std_logic;
  		

  -- state q472
  signal reg_q472        : std_logic;
  signal reg_q472_in     : std_logic;
  		
  signal reg_fullgraph22       : std_logic_vector(1 downto 0);
  signal reg_fullgraph22_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph22_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph22_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph22
  --#################################################			
		

  -- state q1218
  signal reg_q1218        : std_logic;
  signal reg_q1218_in     : std_logic;
  signal reg_q1218_init   : std_logic;
		

  -- state q1061
  signal reg_q1061        : std_logic;
  signal reg_q1061_in     : std_logic;
  signal reg_q1061_init   : std_logic;
		

  -- state q2449
  signal reg_q2449        : std_logic;
  signal reg_q2449_in     : std_logic;
  signal reg_q2449_init   : std_logic;
		

  -- state q497
  signal reg_q497        : std_logic;
  signal reg_q497_in     : std_logic;
  signal reg_q497_init   : std_logic;
		

  -- state q757
  signal reg_q757        : std_logic;
  signal reg_q757_in     : std_logic;
  signal reg_q757_init   : std_logic;
		
--#################################################
-- start section fullgraph: 28

  -- state q1626
  signal reg_q1626        : std_logic;
  signal reg_q1626_in     : std_logic;
  		

  -- state q471
  signal reg_q471        : std_logic;
  signal reg_q471_in     : std_logic;
  		

  -- state q759
  signal reg_q759        : std_logic;
  signal reg_q759_in     : std_logic;
  		
  signal reg_fullgraph28       : std_logic_vector(1 downto 0);
  signal reg_fullgraph28_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph28_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph28_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph28
  --#################################################			
		

  -- state q1951
  signal reg_q1951        : std_logic;
  signal reg_q1951_in     : std_logic;
  signal reg_q1951_init   : std_logic;
		

  -- state q2680
  signal reg_q2680        : std_logic;
  signal reg_q2680_in     : std_logic;
  signal reg_q2680_init   : std_logic;
		

  -- state q2417
  signal reg_q2417        : std_logic;
  signal reg_q2417_in     : std_logic;
  signal reg_q2417_init   : std_logic;
		

  -- state q99
  signal reg_q99        : std_logic;
  signal reg_q99_in     : std_logic;
  signal reg_q99_init   : std_logic;
		
--#################################################
-- start section fullgraph: 33

  -- state q395
  signal reg_q395        : std_logic;
  signal reg_q395_in     : std_logic;
  		

  -- state q526
  signal reg_q526        : std_logic;
  signal reg_q526_in     : std_logic;
  		

  -- state q800
  signal reg_q800        : std_logic;
  signal reg_q800_in     : std_logic;
  		

  -- state q486
  signal reg_q486        : std_logic;
  signal reg_q486_in     : std_logic;
  		

  -- state q1757
  signal reg_q1757        : std_logic;
  signal reg_q1757_in     : std_logic;
  		

  -- state q484
  signal reg_q484        : std_logic;
  signal reg_q484_in     : std_logic;
  		

  -- state q774
  signal reg_q774        : std_logic;
  signal reg_q774_in     : std_logic;
  		
  signal reg_fullgraph33       : std_logic_vector(2 downto 0);
  signal reg_fullgraph33_in    : std_logic_vector(2 downto 0);
  signal reg_fullgraph33_init  : std_logic_vector(2 downto 0);
  signal reg_fullgraph33_sel   : std_logic_vector(7 downto 0); 	
  -- end section fullgraph33
  --#################################################			
		

  -- state q2677
  signal reg_q2677        : std_logic;
  signal reg_q2677_in     : std_logic;
  signal reg_q2677_init   : std_logic;
		

  -- state q1145
  signal reg_q1145        : std_logic;
  signal reg_q1145_in     : std_logic;
  signal reg_q1145_init   : std_logic;
		

  -- state q133
  signal reg_q133        : std_logic;
  signal reg_q133_in     : std_logic;
  signal reg_q133_init   : std_logic;
		

  -- state q1204
  signal reg_q1204        : std_logic;
  signal reg_q1204_in     : std_logic;
  signal reg_q1204_init   : std_logic;
		
--#################################################
-- start section fullgraph: 38

  -- state q2216
  signal reg_q2216        : std_logic;
  signal reg_q2216_in     : std_logic;
  		

  -- state q117
  signal reg_q117        : std_logic;
  signal reg_q117_in     : std_logic;
  		

  -- state q805
  signal reg_q805        : std_logic;
  signal reg_q805_in     : std_logic;
  		
  signal reg_fullgraph38       : std_logic_vector(1 downto 0);
  signal reg_fullgraph38_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph38_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph38_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph38
  --#################################################			
		
--#################################################
-- start section fullgraph: 39

  -- state q397
  signal reg_q397        : std_logic;
  signal reg_q397_in     : std_logic;
  		

  -- state q540
  signal reg_q540        : std_logic;
  signal reg_q540_in     : std_logic;
  		

  -- state q847
  signal reg_q847        : std_logic;
  signal reg_q847_in     : std_logic;
  		

  -- state q855
  signal reg_q855        : std_logic;
  signal reg_q855_in     : std_logic;
  		

  -- state q823
  signal reg_q823        : std_logic;
  signal reg_q823_in     : std_logic;
  		

  -- state q853
  signal reg_q853        : std_logic;
  signal reg_q853_in     : std_logic;
  		

  -- state q845
  signal reg_q845        : std_logic;
  signal reg_q845_in     : std_logic;
  		

  -- state q843
  signal reg_q843        : std_logic;
  signal reg_q843_in     : std_logic;
  		

  -- state q1146
  signal reg_q1146        : std_logic;
  signal reg_q1146_in     : std_logic;
  		

  -- state q849
  signal reg_q849        : std_logic;
  signal reg_q849_in     : std_logic;
  		

  -- state q851
  signal reg_q851        : std_logic;
  signal reg_q851_in     : std_logic;
  		

  -- state q347
  signal reg_q347        : std_logic;
  signal reg_q347_in     : std_logic;
  		

  -- state q880
  signal reg_q880        : std_logic;
  signal reg_q880_in     : std_logic;
  		

  -- state q884
  signal reg_q884        : std_logic;
  signal reg_q884_in     : std_logic;
  		

  -- state q882
  signal reg_q882        : std_logic;
  signal reg_q882_in     : std_logic;
  		
  signal reg_fullgraph39       : std_logic_vector(3 downto 0);
  signal reg_fullgraph39_in    : std_logic_vector(3 downto 0);
  signal reg_fullgraph39_init  : std_logic_vector(3 downto 0);
  signal reg_fullgraph39_sel   : std_logic_vector(15 downto 0); 	
  -- end section fullgraph39
  --#################################################			
		

  -- state q970
  signal reg_q970        : std_logic;
  signal reg_q970_in     : std_logic;
  signal reg_q970_init   : std_logic;
		

  -- state q1096
  signal reg_q1096        : std_logic;
  signal reg_q1096_in     : std_logic;
  signal reg_q1096_init   : std_logic;
		
--#################################################
-- start section fullgraph: 42

  -- state q2218
  signal reg_q2218        : std_logic;
  signal reg_q2218_in     : std_logic;
  		

  -- state q546
  signal reg_q546        : std_logic;
  signal reg_q546_in     : std_logic;
  		

  -- state q592
  signal reg_q592        : std_logic;
  signal reg_q592_in     : std_logic;
  		
  signal reg_fullgraph42       : std_logic_vector(1 downto 0);
  signal reg_fullgraph42_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph42_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph42_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph42
  --#################################################			
		

  -- state q2056
  signal reg_q2056        : std_logic;
  signal reg_q2056_in     : std_logic;
  signal reg_q2056_init   : std_logic;
		

  -- state q1393
  signal reg_q1393        : std_logic;
  signal reg_q1393_in     : std_logic;
  signal reg_q1393_init   : std_logic;
		

  -- state q1685
  signal reg_q1685        : std_logic;
  signal reg_q1685_in     : std_logic;
  signal reg_q1685_init   : std_logic;
		

  -- state q2633
  signal reg_q2633        : std_logic;
  signal reg_q2633_in     : std_logic;
  signal reg_q2633_init   : std_logic;
		

  -- state q1395
  signal reg_q1395        : std_logic;
  signal reg_q1395_in     : std_logic;
  signal reg_q1395_init   : std_logic;
		

  -- state q516
  signal reg_q516        : std_logic;
  signal reg_q516_in     : std_logic;
  signal reg_q516_init   : std_logic;
		

  -- state q1
  signal reg_q1        : std_logic;
  signal reg_q1_in     : std_logic;
  signal reg_q1_init   : std_logic;
		

  -- state q2556
  signal reg_q2556        : std_logic;
  signal reg_q2556_in     : std_logic;
  signal reg_q2556_init   : std_logic;
		

  -- state q399
  signal reg_q399        : std_logic;
  signal reg_q399_in     : std_logic;
  signal reg_q399_init   : std_logic;
		

  -- state q1628
  signal reg_q1628        : std_logic;
  signal reg_q1628_in     : std_logic;
  signal reg_q1628_init   : std_logic;
		

  -- state q2552
  signal reg_q2552        : std_logic;
  signal reg_q2552_in     : std_logic;
  signal reg_q2552_init   : std_logic;
		

  -- state q1482
  signal reg_q1482        : std_logic;
  signal reg_q1482_in     : std_logic;
  signal reg_q1482_init   : std_logic;
		
--#################################################
-- start section fullgraph: 55

  -- state q2080
  signal reg_q2080        : std_logic;
  signal reg_q2080_in     : std_logic;
  		

  -- state q606
  signal reg_q606        : std_logic;
  signal reg_q606_in     : std_logic;
  		

  -- state q342
  signal reg_q342        : std_logic;
  signal reg_q342_in     : std_logic;
  		

  -- state q2435
  signal reg_q2435        : std_logic;
  signal reg_q2435_in     : std_logic;
  		

  -- state q2641
  signal reg_q2641        : std_logic;
  signal reg_q2641_in     : std_logic;
  		

  -- state q435
  signal reg_q435        : std_logic;
  signal reg_q435_in     : std_logic;
  		

  -- state q2116
  signal reg_q2116        : std_logic;
  signal reg_q2116_in     : std_logic;
  		

  -- state q1465
  signal reg_q1465        : std_logic;
  signal reg_q1465_in     : std_logic;
  		

  -- state q2643
  signal reg_q2643        : std_logic;
  signal reg_q2643_in     : std_logic;
  		

  -- state q296
  signal reg_q296        : std_logic;
  signal reg_q296_in     : std_logic;
  		

  -- state q2241
  signal reg_q2241        : std_logic;
  signal reg_q2241_in     : std_logic;
  		

  -- state q2237
  signal reg_q2237        : std_logic;
  signal reg_q2237_in     : std_logic;
  		

  -- state q2647
  signal reg_q2647        : std_logic;
  signal reg_q2647_in     : std_logic;
  		

  -- state q2649
  signal reg_q2649        : std_logic;
  signal reg_q2649_in     : std_logic;
  		

  -- state q1457
  signal reg_q1457        : std_logic;
  signal reg_q1457_in     : std_logic;
  		

  -- state q1411
  signal reg_q1411        : std_logic;
  signal reg_q1411_in     : std_logic;
  		

  -- state q2064
  signal reg_q2064        : std_logic;
  signal reg_q2064_in     : std_logic;
  		

  -- state q1820
  signal reg_q1820        : std_logic;
  signal reg_q1820_in     : std_logic;
  		

  -- state q1463
  signal reg_q1463        : std_logic;
  signal reg_q1463_in     : std_logic;
  		

  -- state q2118
  signal reg_q2118        : std_logic;
  signal reg_q2118_in     : std_logic;
  		

  -- state q294
  signal reg_q294        : std_logic;
  signal reg_q294_in     : std_logic;
  		

  -- state q1034
  signal reg_q1034        : std_logic;
  signal reg_q1034_in     : std_logic;
  		

  -- state q2673
  signal reg_q2673        : std_logic;
  signal reg_q2673_in     : std_logic;
  		

  -- state q2635
  signal reg_q2635        : std_logic;
  signal reg_q2635_in     : std_logic;
  		

  -- state q2637
  signal reg_q2637        : std_logic;
  signal reg_q2637_in     : std_logic;
  		

  -- state q2060
  signal reg_q2060        : std_logic;
  signal reg_q2060_in     : std_logic;
  		

  -- state q2062
  signal reg_q2062        : std_logic;
  signal reg_q2062_in     : std_logic;
  		

  -- state q1369
  signal reg_q1369        : std_logic;
  signal reg_q1369_in     : std_logic;
  		

  -- state q1636
  signal reg_q1636        : std_logic;
  signal reg_q1636_in     : std_logic;
  		

  -- state q2645
  signal reg_q2645        : std_logic;
  signal reg_q2645_in     : std_logic;
  		

  -- state q2433
  signal reg_q2433        : std_logic;
  signal reg_q2433_in     : std_logic;
  		

  -- state q1399
  signal reg_q1399        : std_logic;
  signal reg_q1399_in     : std_logic;
  		

  -- state q2239
  signal reg_q2239        : std_logic;
  signal reg_q2239_in     : std_logic;
  		

  -- state q2122
  signal reg_q2122        : std_logic;
  signal reg_q2122_in     : std_logic;
  		

  -- state q1578
  signal reg_q1578        : std_logic;
  signal reg_q1578_in     : std_logic;
  		

  -- state q1848
  signal reg_q1848        : std_logic;
  signal reg_q1848_in     : std_logic;
  		

  -- state q1389
  signal reg_q1389        : std_logic;
  signal reg_q1389_in     : std_logic;
  		

  -- state q1385
  signal reg_q1385        : std_logic;
  signal reg_q1385_in     : std_logic;
  		

  -- state q1387
  signal reg_q1387        : std_logic;
  signal reg_q1387_in     : std_logic;
  		

  -- state q1644
  signal reg_q1644        : std_logic;
  signal reg_q1644_in     : std_logic;
  		

  -- state q1530
  signal reg_q1530        : std_logic;
  signal reg_q1530_in     : std_logic;
  		

  -- state q1592
  signal reg_q1592        : std_logic;
  signal reg_q1592_in     : std_logic;
  		

  -- state q1884
  signal reg_q1884        : std_logic;
  signal reg_q1884_in     : std_logic;
  		

  -- state q1026
  signal reg_q1026        : std_logic;
  signal reg_q1026_in     : std_logic;
  		

  -- state q2639
  signal reg_q2639        : std_logic;
  signal reg_q2639_in     : std_logic;
  		

  -- state q2074
  signal reg_q2074        : std_logic;
  signal reg_q2074_in     : std_logic;
  		

  -- state q1818
  signal reg_q1818        : std_logic;
  signal reg_q1818_in     : std_logic;
  		

  -- state q1461
  signal reg_q1461        : std_logic;
  signal reg_q1461_in     : std_logic;
  		

  -- state q1634
  signal reg_q1634        : std_logic;
  signal reg_q1634_in     : std_logic;
  		

  -- state q1467
  signal reg_q1467        : std_logic;
  signal reg_q1467_in     : std_logic;
  		

  -- state q2172
  signal reg_q2172        : std_logic;
  signal reg_q2172_in     : std_logic;
  		

  -- state q1640
  signal reg_q1640        : std_logic;
  signal reg_q1640_in     : std_logic;
  		

  -- state q1642
  signal reg_q1642        : std_logic;
  signal reg_q1642_in     : std_logic;
  		

  -- state q1594
  signal reg_q1594        : std_logic;
  signal reg_q1594_in     : std_logic;
  		

  -- state q1365
  signal reg_q1365        : std_logic;
  signal reg_q1365_in     : std_logic;
  		

  -- state q2538
  signal reg_q2538        : std_logic;
  signal reg_q2538_in     : std_logic;
  		

  -- state q1598
  signal reg_q1598        : std_logic;
  signal reg_q1598_in     : std_logic;
  		

  -- state q1270
  signal reg_q1270        : std_logic;
  signal reg_q1270_in     : std_logic;
  		

  -- state q411
  signal reg_q411        : std_logic;
  signal reg_q411_in     : std_logic;
  		

  -- state q1453
  signal reg_q1453        : std_logic;
  signal reg_q1453_in     : std_logic;
  		

  -- state q1469
  signal reg_q1469        : std_logic;
  signal reg_q1469_in     : std_logic;
  		

  -- state q1534
  signal reg_q1534        : std_logic;
  signal reg_q1534_in     : std_logic;
  		

  -- state q461
  signal reg_q461        : std_logic;
  signal reg_q461_in     : std_logic;
  		

  -- state q492
  signal reg_q492        : std_logic;
  signal reg_q492_in     : std_logic;
  		

  -- state q1973
  signal reg_q1973        : std_logic;
  signal reg_q1973_in     : std_logic;
  		

  -- state q2160
  signal reg_q2160        : std_logic;
  signal reg_q2160_in     : std_logic;
  		

  -- state q1028
  signal reg_q1028        : std_logic;
  signal reg_q1028_in     : std_logic;
  		

  -- state q2164
  signal reg_q2164        : std_logic;
  signal reg_q2164_in     : std_logic;
  		
  signal reg_fullgraph55       : std_logic_vector(6 downto 0);
  signal reg_fullgraph55_in    : std_logic_vector(6 downto 0);
  signal reg_fullgraph55_init  : std_logic_vector(6 downto 0);
  signal reg_fullgraph55_sel   : std_logic_vector(127 downto 0); 	
  -- end section fullgraph55
  --#################################################			
		

  -- state q1522
  signal reg_q1522        : std_logic;
  signal reg_q1522_in     : std_logic;
  signal reg_q1522_init   : std_logic;
		

  -- state q661
  signal reg_q661        : std_logic;
  signal reg_q661_in     : std_logic;
  signal reg_q661_init   : std_logic;
		

  -- state q2329
  signal reg_q2329        : std_logic;
  signal reg_q2329_in     : std_logic;
  signal reg_q2329_init   : std_logic;
		

  -- state q803
  signal reg_q803        : std_logic;
  signal reg_q803_in     : std_logic;
  signal reg_q803_init   : std_logic;
		

  -- state q604
  signal reg_q604        : std_logic;
  signal reg_q604_in     : std_logic;
  signal reg_q604_init   : std_logic;
		

  -- state q1574
  signal reg_q1574        : std_logic;
  signal reg_q1574_in     : std_logic;
  signal reg_q1574_init   : std_logic;
		
--#################################################
-- start section fullgraph: 62

  -- state q113
  signal reg_q113        : std_logic;
  signal reg_q113_in     : std_logic;
  		

  -- state q498
  signal reg_q498        : std_logic;
  signal reg_q498_in     : std_logic;
  		
  signal reg_fullgraph62       : std_logic_vector(1 downto 0);
  signal reg_fullgraph62_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph62_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph62_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph62
  --#################################################			
		

  -- state q116
  signal reg_q116        : std_logic;
  signal reg_q116_in     : std_logic;
  signal reg_q116_init   : std_logic;
		
--#################################################
-- start section fullgraph: 64

  -- state q2326
  signal reg_q2326        : std_logic;
  signal reg_q2326_in     : std_logic;
  		

  -- state q2584
  signal reg_q2584        : std_logic;
  signal reg_q2584_in     : std_logic;
  		
  signal reg_fullgraph64       : std_logic_vector(1 downto 0);
  signal reg_fullgraph64_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph64_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph64_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph64
  --#################################################			
		

  -- state q1022
  signal reg_q1022        : std_logic;
  signal reg_q1022_in     : std_logic;
  signal reg_q1022_init   : std_logic;
		

  -- state q2221
  signal reg_q2221        : std_logic;
  signal reg_q2221_in     : std_logic;
  signal reg_q2221_init   : std_logic;
		

  -- state q188
  signal reg_q188        : std_logic;
  signal reg_q188_in     : std_logic;
  signal reg_q188_init   : std_logic;
		

  -- state q1816
  signal reg_q1816        : std_logic;
  signal reg_q1816_in     : std_logic;
  signal reg_q1816_init   : std_logic;
		
--#################################################
-- start section fullgraph: 69

  -- state q298
  signal reg_q298        : std_logic;
  signal reg_q298_in     : std_logic;
  		

  -- state q1620
  signal reg_q1620        : std_logic;
  signal reg_q1620_in     : std_logic;
  		

  -- state q288
  signal reg_q288        : std_logic;
  signal reg_q288_in     : std_logic;
  		

  -- state q2681
  signal reg_q2681        : std_logic;
  signal reg_q2681_in     : std_logic;
  		

  -- state q1965
  signal reg_q1965        : std_logic;
  signal reg_q1965_in     : std_logic;
  		

  -- state q1630
  signal reg_q1630        : std_logic;
  signal reg_q1630_in     : std_logic;
  		

  -- state q1361
  signal reg_q1361        : std_logic;
  signal reg_q1361_in     : std_logic;
  		

  -- state q1391
  signal reg_q1391        : std_logic;
  signal reg_q1391_in     : std_logic;
  		

  -- state q2058
  signal reg_q2058        : std_logic;
  signal reg_q2058_in     : std_logic;
  		

  -- state q2419
  signal reg_q2419        : std_logic;
  signal reg_q2419_in     : std_logic;
  		

  -- state q1584
  signal reg_q1584        : std_logic;
  signal reg_q1584_in     : std_logic;
  		

  -- state q1222
  signal reg_q1222        : std_logic;
  signal reg_q1222_in     : std_logic;
  		

  -- state q1024
  signal reg_q1024        : std_logic;
  signal reg_q1024_in     : std_logic;
  		

  -- state q1459
  signal reg_q1459        : std_logic;
  signal reg_q1459_in     : std_logic;
  		

  -- state q2162
  signal reg_q2162        : std_logic;
  signal reg_q2162_in     : std_logic;
  		
  signal reg_fullgraph69       : std_logic_vector(3 downto 0);
  signal reg_fullgraph69_in    : std_logic_vector(3 downto 0);
  signal reg_fullgraph69_init  : std_logic_vector(3 downto 0);
  signal reg_fullgraph69_sel   : std_logic_vector(15 downto 0); 	
  -- end section fullgraph69
  --#################################################			
		
--#################################################
-- start section fullgraph: 70

  -- state q401
  signal reg_q401        : std_logic;
  signal reg_q401_in     : std_logic;
  		

  -- state q695
  signal reg_q695        : std_logic;
  signal reg_q695_in     : std_logic;
  		

  -- state q1397
  signal reg_q1397        : std_logic;
  signal reg_q1397_in     : std_logic;
  		

  -- state q1676
  signal reg_q1676        : std_logic;
  signal reg_q1676_in     : std_logic;
  		

  -- state q2154
  signal reg_q2154        : std_logic;
  signal reg_q2154_in     : std_logic;
  		

  -- state q2550
  signal reg_q2550        : std_logic;
  signal reg_q2550_in     : std_logic;
  		

  -- state q2505
  signal reg_q2505        : std_logic;
  signal reg_q2505_in     : std_logic;
  		

  -- state q2655
  signal reg_q2655        : std_logic;
  signal reg_q2655_in     : std_logic;
  		

  -- state q2503
  signal reg_q2503        : std_logic;
  signal reg_q2503_in     : std_logic;
  		

  -- state q1652
  signal reg_q1652        : std_logic;
  signal reg_q1652_in     : std_logic;
  		
  signal reg_fullgraph70       : std_logic_vector(3 downto 0);
  signal reg_fullgraph70_in    : std_logic_vector(3 downto 0);
  signal reg_fullgraph70_init  : std_logic_vector(3 downto 0);
  signal reg_fullgraph70_sel   : std_logic_vector(15 downto 0); 	
  -- end section fullgraph70
  --#################################################			
		
--#################################################
-- start section fullgraph: 71

  -- state q2495
  signal reg_q2495        : std_logic;
  signal reg_q2495_in     : std_logic;
  		

  -- state q946
  signal reg_q946        : std_logic;
  signal reg_q946_in     : std_logic;
  		

  -- state q648
  signal reg_q648        : std_logic;
  signal reg_q648_in     : std_logic;
  		

  -- state q310
  signal reg_q310        : std_logic;
  signal reg_q310_in     : std_logic;
  		

  -- state q1576
  signal reg_q1576        : std_logic;
  signal reg_q1576_in     : std_logic;
  		

  -- state q1846
  signal reg_q1846        : std_logic;
  signal reg_q1846_in     : std_logic;
  		

  -- state q455
  signal reg_q455        : std_logic;
  signal reg_q455_in     : std_logic;
  		

  -- state q1447
  signal reg_q1447        : std_logic;
  signal reg_q1447_in     : std_logic;
  		

  -- state q1296
  signal reg_q1296        : std_logic;
  signal reg_q1296_in     : std_logic;
  		

  -- state q894
  signal reg_q894        : std_logic;
  signal reg_q894_in     : std_logic;
  		

  -- state q2487
  signal reg_q2487        : std_logic;
  signal reg_q2487_in     : std_logic;
  		

  -- state q1046
  signal reg_q1046        : std_logic;
  signal reg_q1046_in     : std_logic;
  		

  -- state q1596
  signal reg_q1596        : std_logic;
  signal reg_q1596_in     : std_logic;
  		

  -- state q1363
  signal reg_q1363        : std_logic;
  signal reg_q1363_in     : std_logic;
  		
  signal reg_fullgraph71       : std_logic_vector(3 downto 0);
  signal reg_fullgraph71_in    : std_logic_vector(3 downto 0);
  signal reg_fullgraph71_init  : std_logic_vector(3 downto 0);
  signal reg_fullgraph71_sel   : std_logic_vector(15 downto 0); 	
  -- end section fullgraph71
  --#################################################			
		
--#################################################
-- start section fullgraph: 72

  -- state q1483
  signal reg_q1483        : std_logic;
  signal reg_q1483_in     : std_logic;
  		

  -- state q963
  signal reg_q963        : std_logic;
  signal reg_q963_in     : std_logic;
  		

  -- state q1220
  signal reg_q1220        : std_logic;
  signal reg_q1220_in     : std_logic;
  		
  signal reg_fullgraph72       : std_logic_vector(1 downto 0);
  signal reg_fullgraph72_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph72_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph72_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph72
  --#################################################			
		
--#################################################
-- start section fullgraph: 73

  -- state q861
  signal reg_q861        : std_logic;
  signal reg_q861_in     : std_logic;
  		

  -- state q547
  signal reg_q547        : std_logic;
  signal reg_q547_in     : std_logic;
  		
  signal reg_fullgraph73       : std_logic_vector(1 downto 0);
  signal reg_fullgraph73_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph73_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph73_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph73
  --#################################################			
		

  -- state q134
  signal reg_q134        : std_logic;
  signal reg_q134_in     : std_logic;
  signal reg_q134_init   : std_logic;
		

  -- state q2330
  signal reg_q2330        : std_logic;
  signal reg_q2330_in     : std_logic;
  signal reg_q2330_init   : std_logic;
		

  -- state q346
  signal reg_q346        : std_logic;
  signal reg_q346_in     : std_logic;
  signal reg_q346_init   : std_logic;
		
--#################################################
-- start section fullgraph: 77

  -- state q2294
  signal reg_q2294        : std_logic;
  signal reg_q2294_in     : std_logic;
  		

  -- state q2296
  signal reg_q2296        : std_logic;
  signal reg_q2296_in     : std_logic;
  		
  signal reg_fullgraph77       : std_logic_vector(1 downto 0);
  signal reg_fullgraph77_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph77_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph77_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph77
  --#################################################			
		

  -- state q2521
  signal reg_q2521        : std_logic;
  signal reg_q2521_in     : std_logic;
  signal reg_q2521_init   : std_logic;
		

  -- state q662
  signal reg_q662        : std_logic;
  signal reg_q662_in     : std_logic;
  signal reg_q662_init   : std_logic;
		

  -- state q758
  signal reg_q758        : std_logic;
  signal reg_q758_in     : std_logic;
  signal reg_q758_init   : std_logic;
		

  -- state q189
  signal reg_q189        : std_logic;
  signal reg_q189_in     : std_logic;
  signal reg_q189_init   : std_logic;
		

  -- state q2245
  signal reg_q2245        : std_logic;
  signal reg_q2245_in     : std_logic;
  signal reg_q2245_init   : std_logic;
		

  -- state q1097
  signal reg_q1097        : std_logic;
  signal reg_q1097_in     : std_logic;
  signal reg_q1097_init   : std_logic;
		

  -- state q100
  signal reg_q100        : std_logic;
  signal reg_q100_in     : std_logic;
  signal reg_q100_init   : std_logic;
		

  -- state q804
  signal reg_q804        : std_logic;
  signal reg_q804_in     : std_logic;
  signal reg_q804_init   : std_logic;
		

  -- state q591
  signal reg_q591        : std_logic;
  signal reg_q591_in     : std_logic;
  signal reg_q591_init   : std_logic;
		

  -- state q1310
  signal reg_q1310        : std_logic;
  signal reg_q1310_in     : std_logic;
  signal reg_q1310_init   : std_logic;
		

  -- state q1205
  signal reg_q1205        : std_logic;
  signal reg_q1205_in     : std_logic;
  signal reg_q1205_init   : std_logic;
		

  -- state q517
  signal reg_q517        : std_logic;
  signal reg_q517_in     : std_logic;
  signal reg_q517_init   : std_logic;
		

  -- state q2
  signal reg_q2        : std_logic;
  signal reg_q2_in     : std_logic;
  signal reg_q2_init   : std_logic;
		

  -- state q2222
  signal reg_q2222        : std_logic;
  signal reg_q2222_in     : std_logic;
  signal reg_q2222_init   : std_logic;
		

  -- state q1062
  signal reg_q1062        : std_logic;
  signal reg_q1062_in     : std_logic;
  signal reg_q1062_init   : std_logic;
		

  -- state q971
  signal reg_q971        : std_logic;
  signal reg_q971_in     : std_logic;
  signal reg_q971_init   : std_logic;
		

  -- state q111
  signal reg_q111        : std_logic;
  signal reg_q111_in     : std_logic;
  signal reg_q111_init   : std_logic;
		

  -- symbol decoder
  signal symb_decoder : std_logic_vector(2**DATA_WIDTH - 1 downto 0);

  -- intialization signal
  signal initialize   : std_logic;

	begin
	-- initialization
  	initialize <= INIT OR INPUT_EOF; 
	 
		symb_decoder(16#ca#) <= '1' when (INPUT = X"ca") else
                          '0';
		symb_decoder(16#f4#) <= '1' when (INPUT = X"f4") else
                          '0';
		symb_decoder(16#fa#) <= '1' when (INPUT = X"fa") else
                          '0';
		symb_decoder(16#a0#) <= '1' when (INPUT = X"a0") else
                          '0';
		symb_decoder(16#60#) <= '1' when (INPUT = X"60") else
                          '0';
		symb_decoder(16#f5#) <= '1' when (INPUT = X"f5") else
                          '0';
		symb_decoder(16#cd#) <= '1' when (INPUT = X"cd") else
                          '0';
		symb_decoder(16#98#) <= '1' when (INPUT = X"98") else
                          '0';
		symb_decoder(16#27#) <= '1' when (INPUT = X"27") else
                          '0';
		symb_decoder(16#48#) <= '1' when (INPUT = X"48") else
                          '0';
		symb_decoder(16#7e#) <= '1' when (INPUT = X"7e") else
                          '0';
		symb_decoder(16#20#) <= '1' when (INPUT = X"20") else
                          '0';
		symb_decoder(16#fd#) <= '1' when (INPUT = X"fd") else
                          '0';
		symb_decoder(16#0d#) <= '1' when (INPUT = X"0d") else
                          '0';
		symb_decoder(16#9a#) <= '1' when (INPUT = X"9a") else
                          '0';
		symb_decoder(16#08#) <= '1' when (INPUT = X"08") else
                          '0';
		symb_decoder(16#85#) <= '1' when (INPUT = X"85") else
                          '0';
		symb_decoder(16#82#) <= '1' when (INPUT = X"82") else
                          '0';
		symb_decoder(16#9f#) <= '1' when (INPUT = X"9f") else
                          '0';
		symb_decoder(16#09#) <= '1' when (INPUT = X"09") else
                          '0';
		symb_decoder(16#59#) <= '1' when (INPUT = X"59") else
                          '0';
		symb_decoder(16#c0#) <= '1' when (INPUT = X"c0") else
                          '0';
		symb_decoder(16#ee#) <= '1' when (INPUT = X"ee") else
                          '0';
		symb_decoder(16#51#) <= '1' when (INPUT = X"51") else
                          '0';
		symb_decoder(16#0e#) <= '1' when (INPUT = X"0e") else
                          '0';
		symb_decoder(16#c1#) <= '1' when (INPUT = X"c1") else
                          '0';
		symb_decoder(16#ea#) <= '1' when (INPUT = X"ea") else
                          '0';
		symb_decoder(16#3a#) <= '1' when (INPUT = X"3a") else
                          '0';
		symb_decoder(16#01#) <= '1' when (INPUT = X"01") else
                          '0';
		symb_decoder(16#2c#) <= '1' when (INPUT = X"2c") else
                          '0';
		symb_decoder(16#23#) <= '1' when (INPUT = X"23") else
                          '0';
		symb_decoder(16#f6#) <= '1' when (INPUT = X"f6") else
                          '0';
		symb_decoder(16#07#) <= '1' when (INPUT = X"07") else
                          '0';
		symb_decoder(16#d1#) <= '1' when (INPUT = X"d1") else
                          '0';
		symb_decoder(16#90#) <= '1' when (INPUT = X"90") else
                          '0';
		symb_decoder(16#32#) <= '1' when (INPUT = X"32") else
                          '0';
		symb_decoder(16#ec#) <= '1' when (INPUT = X"ec") else
                          '0';
		symb_decoder(16#73#) <= '1' when (INPUT = X"73") else
                          '0';
		symb_decoder(16#f8#) <= '1' when (INPUT = X"f8") else
                          '0';
		symb_decoder(16#61#) <= '1' when (INPUT = X"61") else
                          '0';
		symb_decoder(16#a3#) <= '1' when (INPUT = X"a3") else
                          '0';
		symb_decoder(16#99#) <= '1' when (INPUT = X"99") else
                          '0';
		symb_decoder(16#b2#) <= '1' when (INPUT = X"b2") else
                          '0';
		symb_decoder(16#f2#) <= '1' when (INPUT = X"f2") else
                          '0';
		symb_decoder(16#29#) <= '1' when (INPUT = X"29") else
                          '0';
		symb_decoder(16#5a#) <= '1' when (INPUT = X"5a") else
                          '0';
		symb_decoder(16#cc#) <= '1' when (INPUT = X"cc") else
                          '0';
		symb_decoder(16#8e#) <= '1' when (INPUT = X"8e") else
                          '0';
		symb_decoder(16#91#) <= '1' when (INPUT = X"91") else
                          '0';
		symb_decoder(16#ff#) <= '1' when (INPUT = X"ff") else
                          '0';
		symb_decoder(16#7c#) <= '1' when (INPUT = X"7c") else
                          '0';
		symb_decoder(16#aa#) <= '1' when (INPUT = X"aa") else
                          '0';
		symb_decoder(16#18#) <= '1' when (INPUT = X"18") else
                          '0';
		symb_decoder(16#02#) <= '1' when (INPUT = X"02") else
                          '0';
		symb_decoder(16#e6#) <= '1' when (INPUT = X"e6") else
                          '0';
		symb_decoder(16#0b#) <= '1' when (INPUT = X"0b") else
                          '0';
		symb_decoder(16#6b#) <= '1' when (INPUT = X"6b") else
                          '0';
		symb_decoder(16#cf#) <= '1' when (INPUT = X"cf") else
                          '0';
		symb_decoder(16#57#) <= '1' when (INPUT = X"57") else
                          '0';
		symb_decoder(16#a8#) <= '1' when (INPUT = X"a8") else
                          '0';
		symb_decoder(16#74#) <= '1' when (INPUT = X"74") else
                          '0';
		symb_decoder(16#7a#) <= '1' when (INPUT = X"7a") else
                          '0';
		symb_decoder(16#8b#) <= '1' when (INPUT = X"8b") else
                          '0';
		symb_decoder(16#04#) <= '1' when (INPUT = X"04") else
                          '0';
		symb_decoder(16#9e#) <= '1' when (INPUT = X"9e") else
                          '0';
		symb_decoder(16#79#) <= '1' when (INPUT = X"79") else
                          '0';
		symb_decoder(16#8a#) <= '1' when (INPUT = X"8a") else
                          '0';
		symb_decoder(16#03#) <= '1' when (INPUT = X"03") else
                          '0';
		symb_decoder(16#10#) <= '1' when (INPUT = X"10") else
                          '0';
		symb_decoder(16#bc#) <= '1' when (INPUT = X"bc") else
                          '0';
		symb_decoder(16#5f#) <= '1' when (INPUT = X"5f") else
                          '0';
		symb_decoder(16#f0#) <= '1' when (INPUT = X"f0") else
                          '0';
		symb_decoder(16#e7#) <= '1' when (INPUT = X"e7") else
                          '0';
		symb_decoder(16#4b#) <= '1' when (INPUT = X"4b") else
                          '0';
		symb_decoder(16#d0#) <= '1' when (INPUT = X"d0") else
                          '0';
		symb_decoder(16#a4#) <= '1' when (INPUT = X"a4") else
                          '0';
		symb_decoder(16#93#) <= '1' when (INPUT = X"93") else
                          '0';
		symb_decoder(16#dd#) <= '1' when (INPUT = X"dd") else
                          '0';
		symb_decoder(16#1d#) <= '1' when (INPUT = X"1d") else
                          '0';
		symb_decoder(16#c4#) <= '1' when (INPUT = X"c4") else
                          '0';
		symb_decoder(16#eb#) <= '1' when (INPUT = X"eb") else
                          '0';
		symb_decoder(16#6d#) <= '1' when (INPUT = X"6d") else
                          '0';
		symb_decoder(16#b7#) <= '1' when (INPUT = X"b7") else
                          '0';
		symb_decoder(16#6a#) <= '1' when (INPUT = X"6a") else
                          '0';
		symb_decoder(16#f7#) <= '1' when (INPUT = X"f7") else
                          '0';
		symb_decoder(16#13#) <= '1' when (INPUT = X"13") else
                          '0';
		symb_decoder(16#b4#) <= '1' when (INPUT = X"b4") else
                          '0';
		symb_decoder(16#12#) <= '1' when (INPUT = X"12") else
                          '0';
		symb_decoder(16#8f#) <= '1' when (INPUT = X"8f") else
                          '0';
		symb_decoder(16#bf#) <= '1' when (INPUT = X"bf") else
                          '0';
		symb_decoder(16#26#) <= '1' when (INPUT = X"26") else
                          '0';
		symb_decoder(16#4a#) <= '1' when (INPUT = X"4a") else
                          '0';
		symb_decoder(16#62#) <= '1' when (INPUT = X"62") else
                          '0';
		symb_decoder(16#e2#) <= '1' when (INPUT = X"e2") else
                          '0';
		symb_decoder(16#3e#) <= '1' when (INPUT = X"3e") else
                          '0';
		symb_decoder(16#56#) <= '1' when (INPUT = X"56") else
                          '0';
		symb_decoder(16#3d#) <= '1' when (INPUT = X"3d") else
                          '0';
		symb_decoder(16#7d#) <= '1' when (INPUT = X"7d") else
                          '0';
		symb_decoder(16#15#) <= '1' when (INPUT = X"15") else
                          '0';
		symb_decoder(16#1c#) <= '1' when (INPUT = X"1c") else
                          '0';
		symb_decoder(16#11#) <= '1' when (INPUT = X"11") else
                          '0';
		symb_decoder(16#71#) <= '1' when (INPUT = X"71") else
                          '0';
		symb_decoder(16#b3#) <= '1' when (INPUT = X"b3") else
                          '0';
		symb_decoder(16#ac#) <= '1' when (INPUT = X"ac") else
                          '0';
		symb_decoder(16#bb#) <= '1' when (INPUT = X"bb") else
                          '0';
		symb_decoder(16#d8#) <= '1' when (INPUT = X"d8") else
                          '0';
		symb_decoder(16#30#) <= '1' when (INPUT = X"30") else
                          '0';
		symb_decoder(16#33#) <= '1' when (INPUT = X"33") else
                          '0';
		symb_decoder(16#22#) <= '1' when (INPUT = X"22") else
                          '0';
		symb_decoder(16#0f#) <= '1' when (INPUT = X"0f") else
                          '0';
		symb_decoder(16#3c#) <= '1' when (INPUT = X"3c") else
                          '0';
		symb_decoder(16#83#) <= '1' when (INPUT = X"83") else
                          '0';
		symb_decoder(16#a5#) <= '1' when (INPUT = X"a5") else
                          '0';
		symb_decoder(16#97#) <= '1' when (INPUT = X"97") else
                          '0';
		symb_decoder(16#1b#) <= '1' when (INPUT = X"1b") else
                          '0';
		symb_decoder(16#ce#) <= '1' when (INPUT = X"ce") else
                          '0';
		symb_decoder(16#c7#) <= '1' when (INPUT = X"c7") else
                          '0';
		symb_decoder(16#b6#) <= '1' when (INPUT = X"b6") else
                          '0';
		symb_decoder(16#c3#) <= '1' when (INPUT = X"c3") else
                          '0';
		symb_decoder(16#53#) <= '1' when (INPUT = X"53") else
                          '0';
		symb_decoder(16#be#) <= '1' when (INPUT = X"be") else
                          '0';
		symb_decoder(16#94#) <= '1' when (INPUT = X"94") else
                          '0';
		symb_decoder(16#9c#) <= '1' when (INPUT = X"9c") else
                          '0';
		symb_decoder(16#ba#) <= '1' when (INPUT = X"ba") else
                          '0';
		symb_decoder(16#a6#) <= '1' when (INPUT = X"a6") else
                          '0';
		symb_decoder(16#b1#) <= '1' when (INPUT = X"b1") else
                          '0';
		symb_decoder(16#1a#) <= '1' when (INPUT = X"1a") else
                          '0';
		symb_decoder(16#31#) <= '1' when (INPUT = X"31") else
                          '0';
		symb_decoder(16#cb#) <= '1' when (INPUT = X"cb") else
                          '0';
		symb_decoder(16#ae#) <= '1' when (INPUT = X"ae") else
                          '0';
		symb_decoder(16#e5#) <= '1' when (INPUT = X"e5") else
                          '0';
		symb_decoder(16#6f#) <= '1' when (INPUT = X"6f") else
                          '0';
		symb_decoder(16#52#) <= '1' when (INPUT = X"52") else
                          '0';
		symb_decoder(16#40#) <= '1' when (INPUT = X"40") else
                          '0';
		symb_decoder(16#80#) <= '1' when (INPUT = X"80") else
                          '0';
		symb_decoder(16#c9#) <= '1' when (INPUT = X"c9") else
                          '0';
		symb_decoder(16#1f#) <= '1' when (INPUT = X"1f") else
                          '0';
		symb_decoder(16#de#) <= '1' when (INPUT = X"de") else
                          '0';
		symb_decoder(16#d6#) <= '1' when (INPUT = X"d6") else
                          '0';
		symb_decoder(16#46#) <= '1' when (INPUT = X"46") else
                          '0';
		symb_decoder(16#af#) <= '1' when (INPUT = X"af") else
                          '0';
		symb_decoder(16#58#) <= '1' when (INPUT = X"58") else
                          '0';
		symb_decoder(16#e0#) <= '1' when (INPUT = X"e0") else
                          '0';
		symb_decoder(16#e9#) <= '1' when (INPUT = X"e9") else
                          '0';
		symb_decoder(16#95#) <= '1' when (INPUT = X"95") else
                          '0';
		symb_decoder(16#81#) <= '1' when (INPUT = X"81") else
                          '0';
		symb_decoder(16#fe#) <= '1' when (INPUT = X"fe") else
                          '0';
		symb_decoder(16#84#) <= '1' when (INPUT = X"84") else
                          '0';
		symb_decoder(16#2f#) <= '1' when (INPUT = X"2f") else
                          '0';
		symb_decoder(16#df#) <= '1' when (INPUT = X"df") else
                          '0';
		symb_decoder(16#d7#) <= '1' when (INPUT = X"d7") else
                          '0';
		symb_decoder(16#25#) <= '1' when (INPUT = X"25") else
                          '0';
		symb_decoder(16#24#) <= '1' when (INPUT = X"24") else
                          '0';
		symb_decoder(16#0a#) <= '1' when (INPUT = X"0a") else
                          '0';
		symb_decoder(16#9d#) <= '1' when (INPUT = X"9d") else
                          '0';
		symb_decoder(16#d5#) <= '1' when (INPUT = X"d5") else
                          '0';
		symb_decoder(16#38#) <= '1' when (INPUT = X"38") else
                          '0';
		symb_decoder(16#44#) <= '1' when (INPUT = X"44") else
                          '0';
		symb_decoder(16#28#) <= '1' when (INPUT = X"28") else
                          '0';
		symb_decoder(16#89#) <= '1' when (INPUT = X"89") else
                          '0';
		symb_decoder(16#34#) <= '1' when (INPUT = X"34") else
                          '0';
		symb_decoder(16#d9#) <= '1' when (INPUT = X"d9") else
                          '0';
		symb_decoder(16#5b#) <= '1' when (INPUT = X"5b") else
                          '0';
		symb_decoder(16#3b#) <= '1' when (INPUT = X"3b") else
                          '0';
		symb_decoder(16#3f#) <= '1' when (INPUT = X"3f") else
                          '0';
		symb_decoder(16#54#) <= '1' when (INPUT = X"54") else
                          '0';
		symb_decoder(16#b9#) <= '1' when (INPUT = X"b9") else
                          '0';
		symb_decoder(16#d2#) <= '1' when (INPUT = X"d2") else
                          '0';
		symb_decoder(16#0c#) <= '1' when (INPUT = X"0c") else
                          '0';
		symb_decoder(16#17#) <= '1' when (INPUT = X"17") else
                          '0';
		symb_decoder(16#f3#) <= '1' when (INPUT = X"f3") else
                          '0';
		symb_decoder(16#36#) <= '1' when (INPUT = X"36") else
                          '0';
		symb_decoder(16#b0#) <= '1' when (INPUT = X"b0") else
                          '0';
		symb_decoder(16#2d#) <= '1' when (INPUT = X"2d") else
                          '0';
		symb_decoder(16#7f#) <= '1' when (INPUT = X"7f") else
                          '0';
		symb_decoder(16#b8#) <= '1' when (INPUT = X"b8") else
                          '0';
		symb_decoder(16#8c#) <= '1' when (INPUT = X"8c") else
                          '0';
		symb_decoder(16#4e#) <= '1' when (INPUT = X"4e") else
                          '0';
		symb_decoder(16#2a#) <= '1' when (INPUT = X"2a") else
                          '0';
		symb_decoder(16#76#) <= '1' when (INPUT = X"76") else
                          '0';
		symb_decoder(16#37#) <= '1' when (INPUT = X"37") else
                          '0';
		symb_decoder(16#87#) <= '1' when (INPUT = X"87") else
                          '0';
		symb_decoder(16#c2#) <= '1' when (INPUT = X"c2") else
                          '0';
		symb_decoder(16#50#) <= '1' when (INPUT = X"50") else
                          '0';
		symb_decoder(16#a9#) <= '1' when (INPUT = X"a9") else
                          '0';
		symb_decoder(16#72#) <= '1' when (INPUT = X"72") else
                          '0';
		symb_decoder(16#db#) <= '1' when (INPUT = X"db") else
                          '0';
		symb_decoder(16#39#) <= '1' when (INPUT = X"39") else
                          '0';
		symb_decoder(16#78#) <= '1' when (INPUT = X"78") else
                          '0';
		symb_decoder(16#4d#) <= '1' when (INPUT = X"4d") else
                          '0';
		symb_decoder(16#c5#) <= '1' when (INPUT = X"c5") else
                          '0';
		symb_decoder(16#19#) <= '1' when (INPUT = X"19") else
                          '0';
		symb_decoder(16#41#) <= '1' when (INPUT = X"41") else
                          '0';
		symb_decoder(16#c6#) <= '1' when (INPUT = X"c6") else
                          '0';
		symb_decoder(16#ab#) <= '1' when (INPUT = X"ab") else
                          '0';
		symb_decoder(16#bd#) <= '1' when (INPUT = X"bd") else
                          '0';
		symb_decoder(16#da#) <= '1' when (INPUT = X"da") else
                          '0';
		symb_decoder(16#a2#) <= '1' when (INPUT = X"a2") else
                          '0';
		symb_decoder(16#55#) <= '1' when (INPUT = X"55") else
                          '0';
		symb_decoder(16#64#) <= '1' when (INPUT = X"64") else
                          '0';
		symb_decoder(16#47#) <= '1' when (INPUT = X"47") else
                          '0';
		symb_decoder(16#5d#) <= '1' when (INPUT = X"5d") else
                          '0';
		symb_decoder(16#5e#) <= '1' when (INPUT = X"5e") else
                          '0';
		symb_decoder(16#1e#) <= '1' when (INPUT = X"1e") else
                          '0';
		symb_decoder(16#fc#) <= '1' when (INPUT = X"fc") else
                          '0';
		symb_decoder(16#ef#) <= '1' when (INPUT = X"ef") else
                          '0';
		symb_decoder(16#77#) <= '1' when (INPUT = X"77") else
                          '0';
		symb_decoder(16#5c#) <= '1' when (INPUT = X"5c") else
                          '0';
		symb_decoder(16#43#) <= '1' when (INPUT = X"43") else
                          '0';
		symb_decoder(16#2e#) <= '1' when (INPUT = X"2e") else
                          '0';
		symb_decoder(16#a7#) <= '1' when (INPUT = X"a7") else
                          '0';
		symb_decoder(16#e1#) <= '1' when (INPUT = X"e1") else
                          '0';
		symb_decoder(16#05#) <= '1' when (INPUT = X"05") else
                          '0';
		symb_decoder(16#e4#) <= '1' when (INPUT = X"e4") else
                          '0';
		symb_decoder(16#35#) <= '1' when (INPUT = X"35") else
                          '0';
		symb_decoder(16#e3#) <= '1' when (INPUT = X"e3") else
                          '0';
		symb_decoder(16#00#) <= '1' when (INPUT = X"00") else
                          '0';
		symb_decoder(16#d4#) <= '1' when (INPUT = X"d4") else
                          '0';
		symb_decoder(16#45#) <= '1' when (INPUT = X"45") else
                          '0';
		symb_decoder(16#66#) <= '1' when (INPUT = X"66") else
                          '0';
		symb_decoder(16#75#) <= '1' when (INPUT = X"75") else
                          '0';
		symb_decoder(16#ad#) <= '1' when (INPUT = X"ad") else
                          '0';
		symb_decoder(16#fb#) <= '1' when (INPUT = X"fb") else
                          '0';
		symb_decoder(16#f9#) <= '1' when (INPUT = X"f9") else
                          '0';
		symb_decoder(16#4c#) <= '1' when (INPUT = X"4c") else
                          '0';
		symb_decoder(16#70#) <= '1' when (INPUT = X"70") else
                          '0';
		symb_decoder(16#7b#) <= '1' when (INPUT = X"7b") else
                          '0';
		symb_decoder(16#68#) <= '1' when (INPUT = X"68") else
                          '0';
		symb_decoder(16#dc#) <= '1' when (INPUT = X"dc") else
                          '0';
		symb_decoder(16#92#) <= '1' when (INPUT = X"92") else
                          '0';
		symb_decoder(16#d3#) <= '1' when (INPUT = X"d3") else
                          '0';
		symb_decoder(16#42#) <= '1' when (INPUT = X"42") else
                          '0';
		symb_decoder(16#96#) <= '1' when (INPUT = X"96") else
                          '0';
		symb_decoder(16#e8#) <= '1' when (INPUT = X"e8") else
                          '0';
		symb_decoder(16#6c#) <= '1' when (INPUT = X"6c") else
                          '0';
		symb_decoder(16#c8#) <= '1' when (INPUT = X"c8") else
                          '0';
		symb_decoder(16#14#) <= '1' when (INPUT = X"14") else
                          '0';
		symb_decoder(16#06#) <= '1' when (INPUT = X"06") else
                          '0';
		symb_decoder(16#8d#) <= '1' when (INPUT = X"8d") else
                          '0';
		symb_decoder(16#69#) <= '1' when (INPUT = X"69") else
                          '0';
		symb_decoder(16#86#) <= '1' when (INPUT = X"86") else
                          '0';
		symb_decoder(16#f1#) <= '1' when (INPUT = X"f1") else
                          '0';
		symb_decoder(16#65#) <= '1' when (INPUT = X"65") else
                          '0';
		symb_decoder(16#67#) <= '1' when (INPUT = X"67") else
                          '0';
		symb_decoder(16#9b#) <= '1' when (INPUT = X"9b") else
                          '0';
		symb_decoder(16#ed#) <= '1' when (INPUT = X"ed") else
                          '0';
		symb_decoder(16#6e#) <= '1' when (INPUT = X"6e") else
                          '0';
		symb_decoder(16#88#) <= '1' when (INPUT = X"88") else
                          '0';
		symb_decoder(16#4f#) <= '1' when (INPUT = X"4f") else
                          '0';
		symb_decoder(16#21#) <= '1' when (INPUT = X"21") else
                          '0';
		symb_decoder(16#a1#) <= '1' when (INPUT = X"a1") else
                          '0';
		symb_decoder(16#2b#) <= '1' when (INPUT = X"2b") else
                          '0';
		symb_decoder(16#16#) <= '1' when (INPUT = X"16") else
                          '0';
		symb_decoder(16#63#) <= '1' when (INPUT = X"63") else
                          '0';
		symb_decoder(16#49#) <= '1' when (INPUT = X"49") else
                          '0';
		symb_decoder(16#b5#) <= '1' when (INPUT = X"b5") else
                          '0';

--######################################################
--fullgraph0

reg_q345_in <= (reg_q345 AND symb_decoder(16#ca#)) OR
 					(reg_q345 AND symb_decoder(16#f4#)) OR
 					(reg_q345 AND symb_decoder(16#fa#)) OR
 					(reg_q345 AND symb_decoder(16#a0#)) OR
 					(reg_q345 AND symb_decoder(16#60#)) OR
 					(reg_q345 AND symb_decoder(16#f5#)) OR
 					(reg_q345 AND symb_decoder(16#cd#)) OR
 					(reg_q345 AND symb_decoder(16#98#)) OR
 					(reg_q345 AND symb_decoder(16#27#)) OR
 					(reg_q345 AND symb_decoder(16#48#)) OR
 					(reg_q345 AND symb_decoder(16#7e#)) OR
 					(reg_q345 AND symb_decoder(16#20#)) OR
 					(reg_q345 AND symb_decoder(16#fd#)) OR
 					(reg_q345 AND symb_decoder(16#0d#)) OR
 					(reg_q345 AND symb_decoder(16#9a#)) OR
 					(reg_q345 AND symb_decoder(16#08#)) OR
 					(reg_q345 AND symb_decoder(16#85#)) OR
 					(reg_q345 AND symb_decoder(16#82#)) OR
 					(reg_q345 AND symb_decoder(16#9f#)) OR
 					(reg_q345 AND symb_decoder(16#09#)) OR
 					(reg_q345 AND symb_decoder(16#59#)) OR
 					(reg_q345 AND symb_decoder(16#c0#)) OR
 					(reg_q345 AND symb_decoder(16#ee#)) OR
 					(reg_q345 AND symb_decoder(16#51#)) OR
 					(reg_q345 AND symb_decoder(16#0e#)) OR
 					(reg_q345 AND symb_decoder(16#c1#)) OR
 					(reg_q345 AND symb_decoder(16#ea#)) OR
 					(reg_q345 AND symb_decoder(16#3a#)) OR
 					(reg_q345 AND symb_decoder(16#01#)) OR
 					(reg_q345 AND symb_decoder(16#2c#)) OR
 					(reg_q345 AND symb_decoder(16#23#)) OR
 					(reg_q345 AND symb_decoder(16#f6#)) OR
 					(reg_q345 AND symb_decoder(16#07#)) OR
 					(reg_q345 AND symb_decoder(16#d1#)) OR
 					(reg_q345 AND symb_decoder(16#90#)) OR
 					(reg_q345 AND symb_decoder(16#32#)) OR
 					(reg_q345 AND symb_decoder(16#ec#)) OR
 					(reg_q345 AND symb_decoder(16#73#)) OR
 					(reg_q345 AND symb_decoder(16#f8#)) OR
 					(reg_q345 AND symb_decoder(16#61#)) OR
 					(reg_q345 AND symb_decoder(16#a3#)) OR
 					(reg_q345 AND symb_decoder(16#99#)) OR
 					(reg_q345 AND symb_decoder(16#b2#)) OR
 					(reg_q345 AND symb_decoder(16#f2#)) OR
 					(reg_q345 AND symb_decoder(16#29#)) OR
 					(reg_q345 AND symb_decoder(16#5a#)) OR
 					(reg_q345 AND symb_decoder(16#cc#)) OR
 					(reg_q345 AND symb_decoder(16#8e#)) OR
 					(reg_q345 AND symb_decoder(16#91#)) OR
 					(reg_q345 AND symb_decoder(16#ff#)) OR
 					(reg_q345 AND symb_decoder(16#7c#)) OR
 					(reg_q345 AND symb_decoder(16#aa#)) OR
 					(reg_q345 AND symb_decoder(16#18#)) OR
 					(reg_q345 AND symb_decoder(16#02#)) OR
 					(reg_q345 AND symb_decoder(16#e6#)) OR
 					(reg_q345 AND symb_decoder(16#0b#)) OR
 					(reg_q345 AND symb_decoder(16#6b#)) OR
 					(reg_q345 AND symb_decoder(16#cf#)) OR
 					(reg_q345 AND symb_decoder(16#57#)) OR
 					(reg_q345 AND symb_decoder(16#a8#)) OR
 					(reg_q345 AND symb_decoder(16#74#)) OR
 					(reg_q345 AND symb_decoder(16#7a#)) OR
 					(reg_q345 AND symb_decoder(16#8b#)) OR
 					(reg_q345 AND symb_decoder(16#04#)) OR
 					(reg_q345 AND symb_decoder(16#9e#)) OR
 					(reg_q345 AND symb_decoder(16#79#)) OR
 					(reg_q345 AND symb_decoder(16#8a#)) OR
 					(reg_q345 AND symb_decoder(16#03#)) OR
 					(reg_q345 AND symb_decoder(16#10#)) OR
 					(reg_q345 AND symb_decoder(16#bc#)) OR
 					(reg_q345 AND symb_decoder(16#5f#)) OR
 					(reg_q345 AND symb_decoder(16#f0#)) OR
 					(reg_q345 AND symb_decoder(16#e7#)) OR
 					(reg_q345 AND symb_decoder(16#4b#)) OR
 					(reg_q345 AND symb_decoder(16#d0#)) OR
 					(reg_q345 AND symb_decoder(16#a4#)) OR
 					(reg_q345 AND symb_decoder(16#93#)) OR
 					(reg_q345 AND symb_decoder(16#dd#)) OR
 					(reg_q345 AND symb_decoder(16#1d#)) OR
 					(reg_q345 AND symb_decoder(16#c4#)) OR
 					(reg_q345 AND symb_decoder(16#eb#)) OR
 					(reg_q345 AND symb_decoder(16#6d#)) OR
 					(reg_q345 AND symb_decoder(16#b7#)) OR
 					(reg_q345 AND symb_decoder(16#6a#)) OR
 					(reg_q345 AND symb_decoder(16#f7#)) OR
 					(reg_q345 AND symb_decoder(16#13#)) OR
 					(reg_q345 AND symb_decoder(16#b4#)) OR
 					(reg_q345 AND symb_decoder(16#12#)) OR
 					(reg_q345 AND symb_decoder(16#8f#)) OR
 					(reg_q345 AND symb_decoder(16#bf#)) OR
 					(reg_q345 AND symb_decoder(16#26#)) OR
 					(reg_q345 AND symb_decoder(16#4a#)) OR
 					(reg_q345 AND symb_decoder(16#62#)) OR
 					(reg_q345 AND symb_decoder(16#e2#)) OR
 					(reg_q345 AND symb_decoder(16#3e#)) OR
 					(reg_q345 AND symb_decoder(16#56#)) OR
 					(reg_q345 AND symb_decoder(16#3d#)) OR
 					(reg_q345 AND symb_decoder(16#7d#)) OR
 					(reg_q345 AND symb_decoder(16#15#)) OR
 					(reg_q345 AND symb_decoder(16#1c#)) OR
 					(reg_q345 AND symb_decoder(16#11#)) OR
 					(reg_q345 AND symb_decoder(16#71#)) OR
 					(reg_q345 AND symb_decoder(16#b3#)) OR
 					(reg_q345 AND symb_decoder(16#ac#)) OR
 					(reg_q345 AND symb_decoder(16#bb#)) OR
 					(reg_q345 AND symb_decoder(16#d8#)) OR
 					(reg_q345 AND symb_decoder(16#30#)) OR
 					(reg_q345 AND symb_decoder(16#33#)) OR
 					(reg_q345 AND symb_decoder(16#22#)) OR
 					(reg_q345 AND symb_decoder(16#0f#)) OR
 					(reg_q345 AND symb_decoder(16#3c#)) OR
 					(reg_q345 AND symb_decoder(16#83#)) OR
 					(reg_q345 AND symb_decoder(16#a5#)) OR
 					(reg_q345 AND symb_decoder(16#97#)) OR
 					(reg_q345 AND symb_decoder(16#1b#)) OR
 					(reg_q345 AND symb_decoder(16#ce#)) OR
 					(reg_q345 AND symb_decoder(16#c7#)) OR
 					(reg_q345 AND symb_decoder(16#b6#)) OR
 					(reg_q345 AND symb_decoder(16#c3#)) OR
 					(reg_q345 AND symb_decoder(16#53#)) OR
 					(reg_q345 AND symb_decoder(16#be#)) OR
 					(reg_q345 AND symb_decoder(16#94#)) OR
 					(reg_q345 AND symb_decoder(16#9c#)) OR
 					(reg_q345 AND symb_decoder(16#ba#)) OR
 					(reg_q345 AND symb_decoder(16#a6#)) OR
 					(reg_q345 AND symb_decoder(16#b1#)) OR
 					(reg_q345 AND symb_decoder(16#1a#)) OR
 					(reg_q345 AND symb_decoder(16#31#)) OR
 					(reg_q345 AND symb_decoder(16#cb#)) OR
 					(reg_q345 AND symb_decoder(16#ae#)) OR
 					(reg_q345 AND symb_decoder(16#e5#)) OR
 					(reg_q345 AND symb_decoder(16#6f#)) OR
 					(reg_q345 AND symb_decoder(16#52#)) OR
 					(reg_q345 AND symb_decoder(16#40#)) OR
 					(reg_q345 AND symb_decoder(16#80#)) OR
 					(reg_q345 AND symb_decoder(16#c9#)) OR
 					(reg_q345 AND symb_decoder(16#1f#)) OR
 					(reg_q345 AND symb_decoder(16#de#)) OR
 					(reg_q345 AND symb_decoder(16#d6#)) OR
 					(reg_q345 AND symb_decoder(16#46#)) OR
 					(reg_q345 AND symb_decoder(16#af#)) OR
 					(reg_q345 AND symb_decoder(16#58#)) OR
 					(reg_q345 AND symb_decoder(16#e0#)) OR
 					(reg_q345 AND symb_decoder(16#e9#)) OR
 					(reg_q345 AND symb_decoder(16#95#)) OR
 					(reg_q345 AND symb_decoder(16#81#)) OR
 					(reg_q345 AND symb_decoder(16#fe#)) OR
 					(reg_q345 AND symb_decoder(16#84#)) OR
 					(reg_q345 AND symb_decoder(16#2f#)) OR
 					(reg_q345 AND symb_decoder(16#df#)) OR
 					(reg_q345 AND symb_decoder(16#d7#)) OR
 					(reg_q345 AND symb_decoder(16#25#)) OR
 					(reg_q345 AND symb_decoder(16#24#)) OR
 					(reg_q345 AND symb_decoder(16#0a#)) OR
 					(reg_q345 AND symb_decoder(16#9d#)) OR
 					(reg_q345 AND symb_decoder(16#d5#)) OR
 					(reg_q345 AND symb_decoder(16#38#)) OR
 					(reg_q345 AND symb_decoder(16#44#)) OR
 					(reg_q345 AND symb_decoder(16#28#)) OR
 					(reg_q345 AND symb_decoder(16#89#)) OR
 					(reg_q345 AND symb_decoder(16#34#)) OR
 					(reg_q345 AND symb_decoder(16#d9#)) OR
 					(reg_q345 AND symb_decoder(16#5b#)) OR
 					(reg_q345 AND symb_decoder(16#3b#)) OR
 					(reg_q345 AND symb_decoder(16#3f#)) OR
 					(reg_q345 AND symb_decoder(16#54#)) OR
 					(reg_q345 AND symb_decoder(16#b9#)) OR
 					(reg_q345 AND symb_decoder(16#d2#)) OR
 					(reg_q345 AND symb_decoder(16#0c#)) OR
 					(reg_q345 AND symb_decoder(16#17#)) OR
 					(reg_q345 AND symb_decoder(16#f3#)) OR
 					(reg_q345 AND symb_decoder(16#36#)) OR
 					(reg_q345 AND symb_decoder(16#b0#)) OR
 					(reg_q345 AND symb_decoder(16#2d#)) OR
 					(reg_q345 AND symb_decoder(16#7f#)) OR
 					(reg_q345 AND symb_decoder(16#b8#)) OR
 					(reg_q345 AND symb_decoder(16#8c#)) OR
 					(reg_q345 AND symb_decoder(16#4e#)) OR
 					(reg_q345 AND symb_decoder(16#2a#)) OR
 					(reg_q345 AND symb_decoder(16#76#)) OR
 					(reg_q345 AND symb_decoder(16#37#)) OR
 					(reg_q345 AND symb_decoder(16#87#)) OR
 					(reg_q345 AND symb_decoder(16#c2#)) OR
 					(reg_q345 AND symb_decoder(16#50#)) OR
 					(reg_q345 AND symb_decoder(16#a9#)) OR
 					(reg_q345 AND symb_decoder(16#72#)) OR
 					(reg_q345 AND symb_decoder(16#db#)) OR
 					(reg_q345 AND symb_decoder(16#39#)) OR
 					(reg_q345 AND symb_decoder(16#78#)) OR
 					(reg_q345 AND symb_decoder(16#4d#)) OR
 					(reg_q345 AND symb_decoder(16#c5#)) OR
 					(reg_q345 AND symb_decoder(16#19#)) OR
 					(reg_q345 AND symb_decoder(16#41#)) OR
 					(reg_q345 AND symb_decoder(16#c6#)) OR
 					(reg_q345 AND symb_decoder(16#ab#)) OR
 					(reg_q345 AND symb_decoder(16#bd#)) OR
 					(reg_q345 AND symb_decoder(16#da#)) OR
 					(reg_q345 AND symb_decoder(16#a2#)) OR
 					(reg_q345 AND symb_decoder(16#55#)) OR
 					(reg_q345 AND symb_decoder(16#64#)) OR
 					(reg_q345 AND symb_decoder(16#47#)) OR
 					(reg_q345 AND symb_decoder(16#5d#)) OR
 					(reg_q345 AND symb_decoder(16#5e#)) OR
 					(reg_q345 AND symb_decoder(16#1e#)) OR
 					(reg_q345 AND symb_decoder(16#fc#)) OR
 					(reg_q345 AND symb_decoder(16#ef#)) OR
 					(reg_q345 AND symb_decoder(16#77#)) OR
 					(reg_q345 AND symb_decoder(16#5c#)) OR
 					(reg_q345 AND symb_decoder(16#43#)) OR
 					(reg_q345 AND symb_decoder(16#2e#)) OR
 					(reg_q345 AND symb_decoder(16#a7#)) OR
 					(reg_q345 AND symb_decoder(16#e1#)) OR
 					(reg_q345 AND symb_decoder(16#05#)) OR
 					(reg_q345 AND symb_decoder(16#e4#)) OR
 					(reg_q345 AND symb_decoder(16#35#)) OR
 					(reg_q345 AND symb_decoder(16#e3#)) OR
 					(reg_q345 AND symb_decoder(16#00#)) OR
 					(reg_q345 AND symb_decoder(16#d4#)) OR
 					(reg_q345 AND symb_decoder(16#45#)) OR
 					(reg_q345 AND symb_decoder(16#66#)) OR
 					(reg_q345 AND symb_decoder(16#75#)) OR
 					(reg_q345 AND symb_decoder(16#ad#)) OR
 					(reg_q345 AND symb_decoder(16#fb#)) OR
 					(reg_q345 AND symb_decoder(16#f9#)) OR
 					(reg_q345 AND symb_decoder(16#4c#)) OR
 					(reg_q345 AND symb_decoder(16#70#)) OR
 					(reg_q345 AND symb_decoder(16#7b#)) OR
 					(reg_q345 AND symb_decoder(16#68#)) OR
 					(reg_q345 AND symb_decoder(16#dc#)) OR
 					(reg_q345 AND symb_decoder(16#92#)) OR
 					(reg_q345 AND symb_decoder(16#d3#)) OR
 					(reg_q345 AND symb_decoder(16#42#)) OR
 					(reg_q345 AND symb_decoder(16#96#)) OR
 					(reg_q345 AND symb_decoder(16#e8#)) OR
 					(reg_q345 AND symb_decoder(16#6c#)) OR
 					(reg_q345 AND symb_decoder(16#c8#)) OR
 					(reg_q345 AND symb_decoder(16#14#)) OR
 					(reg_q345 AND symb_decoder(16#06#)) OR
 					(reg_q345 AND symb_decoder(16#8d#)) OR
 					(reg_q345 AND symb_decoder(16#69#)) OR
 					(reg_q345 AND symb_decoder(16#86#)) OR
 					(reg_q345 AND symb_decoder(16#f1#)) OR
 					(reg_q345 AND symb_decoder(16#65#)) OR
 					(reg_q345 AND symb_decoder(16#67#)) OR
 					(reg_q345 AND symb_decoder(16#9b#)) OR
 					(reg_q345 AND symb_decoder(16#ed#)) OR
 					(reg_q345 AND symb_decoder(16#6e#)) OR
 					(reg_q345 AND symb_decoder(16#88#)) OR
 					(reg_q345 AND symb_decoder(16#4f#)) OR
 					(reg_q345 AND symb_decoder(16#21#)) OR
 					(reg_q345 AND symb_decoder(16#a1#)) OR
 					(reg_q345 AND symb_decoder(16#2b#)) OR
 					(reg_q345 AND symb_decoder(16#16#)) OR
 					(reg_q345 AND symb_decoder(16#63#)) OR
 					(reg_q345 AND symb_decoder(16#49#)) OR
 					(reg_q345 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#));
reg_q2757_in <= '0';
reg_fullgraph0_init <= "10";

reg_fullgraph0_sel <= "00" & reg_q2757_in & reg_q345_in;

	--coder fullgraph0
with reg_fullgraph0_sel select
reg_fullgraph0_in <=
	"01" when "0001",
	"10" when "0010",
	"00" when others;
 --end coder

	p_reg_fullgraph0: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph0 <= reg_fullgraph0_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph0 <= reg_fullgraph0_init;
        else
          reg_fullgraph0 <= reg_fullgraph0_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph0

		reg_q345 <= '1' when reg_fullgraph0 = "01" else '0'; 
		reg_q2757 <= '1' when reg_fullgraph0 = "10" else '0'; 
--end decoder 
--######################################################
--fullgraph1

reg_q565_in <= (reg_q563 AND symb_decoder(16#23#));
reg_q587_in <= (reg_q565 AND symb_decoder(16#33#)) OR
 					(reg_q565 AND symb_decoder(16#4b#)) OR
 					(reg_q565 AND symb_decoder(16#08#)) OR
 					(reg_q565 AND symb_decoder(16#4e#)) OR
 					(reg_q565 AND symb_decoder(16#6e#)) OR
 					(reg_q565 AND symb_decoder(16#62#)) OR
 					(reg_q565 AND symb_decoder(16#a4#)) OR
 					(reg_q565 AND symb_decoder(16#90#)) OR
 					(reg_q565 AND symb_decoder(16#20#)) OR
 					(reg_q565 AND symb_decoder(16#75#)) OR
 					(reg_q565 AND symb_decoder(16#71#)) OR
 					(reg_q565 AND symb_decoder(16#e4#)) OR
 					(reg_q565 AND symb_decoder(16#12#)) OR
 					(reg_q565 AND symb_decoder(16#01#)) OR
 					(reg_q565 AND symb_decoder(16#e1#)) OR
 					(reg_q565 AND symb_decoder(16#87#)) OR
 					(reg_q565 AND symb_decoder(16#7c#)) OR
 					(reg_q565 AND symb_decoder(16#88#)) OR
 					(reg_q565 AND symb_decoder(16#9f#)) OR
 					(reg_q565 AND symb_decoder(16#9c#)) OR
 					(reg_q565 AND symb_decoder(16#49#)) OR
 					(reg_q565 AND symb_decoder(16#ef#)) OR
 					(reg_q565 AND symb_decoder(16#7d#)) OR
 					(reg_q565 AND symb_decoder(16#b9#)) OR
 					(reg_q565 AND symb_decoder(16#70#)) OR
 					(reg_q565 AND symb_decoder(16#4c#)) OR
 					(reg_q565 AND symb_decoder(16#26#)) OR
 					(reg_q565 AND symb_decoder(16#6d#)) OR
 					(reg_q565 AND symb_decoder(16#02#)) OR
 					(reg_q565 AND symb_decoder(16#b6#)) OR
 					(reg_q565 AND symb_decoder(16#0b#)) OR
 					(reg_q565 AND symb_decoder(16#10#)) OR
 					(reg_q565 AND symb_decoder(16#a1#)) OR
 					(reg_q565 AND symb_decoder(16#92#)) OR
 					(reg_q565 AND symb_decoder(16#36#)) OR
 					(reg_q565 AND symb_decoder(16#30#)) OR
 					(reg_q565 AND symb_decoder(16#40#)) OR
 					(reg_q565 AND symb_decoder(16#41#)) OR
 					(reg_q565 AND symb_decoder(16#16#)) OR
 					(reg_q565 AND symb_decoder(16#fa#)) OR
 					(reg_q565 AND symb_decoder(16#5b#)) OR
 					(reg_q565 AND symb_decoder(16#c7#)) OR
 					(reg_q565 AND symb_decoder(16#5c#)) OR
 					(reg_q565 AND symb_decoder(16#42#)) OR
 					(reg_q565 AND symb_decoder(16#db#)) OR
 					(reg_q565 AND symb_decoder(16#23#)) OR
 					(reg_q565 AND symb_decoder(16#68#)) OR
 					(reg_q565 AND symb_decoder(16#00#)) OR
 					(reg_q565 AND symb_decoder(16#1d#)) OR
 					(reg_q565 AND symb_decoder(16#2a#)) OR
 					(reg_q565 AND symb_decoder(16#d1#)) OR
 					(reg_q565 AND symb_decoder(16#c0#)) OR
 					(reg_q565 AND symb_decoder(16#fd#)) OR
 					(reg_q565 AND symb_decoder(16#f3#)) OR
 					(reg_q565 AND symb_decoder(16#f5#)) OR
 					(reg_q565 AND symb_decoder(16#5e#)) OR
 					(reg_q565 AND symb_decoder(16#f2#)) OR
 					(reg_q565 AND symb_decoder(16#56#)) OR
 					(reg_q565 AND symb_decoder(16#4a#)) OR
 					(reg_q565 AND symb_decoder(16#6b#)) OR
 					(reg_q565 AND symb_decoder(16#f9#)) OR
 					(reg_q565 AND symb_decoder(16#3d#)) OR
 					(reg_q565 AND symb_decoder(16#7f#)) OR
 					(reg_q565 AND symb_decoder(16#b8#)) OR
 					(reg_q565 AND symb_decoder(16#bb#)) OR
 					(reg_q565 AND symb_decoder(16#91#)) OR
 					(reg_q565 AND symb_decoder(16#b0#)) OR
 					(reg_q565 AND symb_decoder(16#59#)) OR
 					(reg_q565 AND symb_decoder(16#96#)) OR
 					(reg_q565 AND symb_decoder(16#d6#)) OR
 					(reg_q565 AND symb_decoder(16#a0#)) OR
 					(reg_q565 AND symb_decoder(16#53#)) OR
 					(reg_q565 AND symb_decoder(16#ac#)) OR
 					(reg_q565 AND symb_decoder(16#0f#)) OR
 					(reg_q565 AND symb_decoder(16#67#)) OR
 					(reg_q565 AND symb_decoder(16#f6#)) OR
 					(reg_q565 AND symb_decoder(16#0c#)) OR
 					(reg_q565 AND symb_decoder(16#d3#)) OR
 					(reg_q565 AND symb_decoder(16#5f#)) OR
 					(reg_q565 AND symb_decoder(16#29#)) OR
 					(reg_q565 AND symb_decoder(16#3a#)) OR
 					(reg_q565 AND symb_decoder(16#17#)) OR
 					(reg_q565 AND symb_decoder(16#04#)) OR
 					(reg_q565 AND symb_decoder(16#51#)) OR
 					(reg_q565 AND symb_decoder(16#b3#)) OR
 					(reg_q565 AND symb_decoder(16#fc#)) OR
 					(reg_q565 AND symb_decoder(16#b4#)) OR
 					(reg_q565 AND symb_decoder(16#1f#)) OR
 					(reg_q565 AND symb_decoder(16#05#)) OR
 					(reg_q565 AND symb_decoder(16#f1#)) OR
 					(reg_q565 AND symb_decoder(16#9b#)) OR
 					(reg_q565 AND symb_decoder(16#39#)) OR
 					(reg_q565 AND symb_decoder(16#cd#)) OR
 					(reg_q565 AND symb_decoder(16#2f#)) OR
 					(reg_q565 AND symb_decoder(16#37#)) OR
 					(reg_q565 AND symb_decoder(16#2c#)) OR
 					(reg_q565 AND symb_decoder(16#ec#)) OR
 					(reg_q565 AND symb_decoder(16#52#)) OR
 					(reg_q565 AND symb_decoder(16#8a#)) OR
 					(reg_q565 AND symb_decoder(16#81#)) OR
 					(reg_q565 AND symb_decoder(16#a9#)) OR
 					(reg_q565 AND symb_decoder(16#9d#)) OR
 					(reg_q565 AND symb_decoder(16#21#)) OR
 					(reg_q565 AND symb_decoder(16#14#)) OR
 					(reg_q565 AND symb_decoder(16#73#)) OR
 					(reg_q565 AND symb_decoder(16#45#)) OR
 					(reg_q565 AND symb_decoder(16#f4#)) OR
 					(reg_q565 AND symb_decoder(16#c1#)) OR
 					(reg_q565 AND symb_decoder(16#a2#)) OR
 					(reg_q565 AND symb_decoder(16#5a#)) OR
 					(reg_q565 AND symb_decoder(16#ed#)) OR
 					(reg_q565 AND symb_decoder(16#e0#)) OR
 					(reg_q565 AND symb_decoder(16#35#)) OR
 					(reg_q565 AND symb_decoder(16#27#)) OR
 					(reg_q565 AND symb_decoder(16#78#)) OR
 					(reg_q565 AND symb_decoder(16#48#)) OR
 					(reg_q565 AND symb_decoder(16#77#)) OR
 					(reg_q565 AND symb_decoder(16#a8#)) OR
 					(reg_q565 AND symb_decoder(16#c4#)) OR
 					(reg_q565 AND symb_decoder(16#38#)) OR
 					(reg_q565 AND symb_decoder(16#25#)) OR
 					(reg_q565 AND symb_decoder(16#eb#)) OR
 					(reg_q565 AND symb_decoder(16#15#)) OR
 					(reg_q565 AND symb_decoder(16#c6#)) OR
 					(reg_q565 AND symb_decoder(16#cc#)) OR
 					(reg_q565 AND symb_decoder(16#79#)) OR
 					(reg_q565 AND symb_decoder(16#cb#)) OR
 					(reg_q565 AND symb_decoder(16#99#)) OR
 					(reg_q565 AND symb_decoder(16#8f#)) OR
 					(reg_q565 AND symb_decoder(16#bc#)) OR
 					(reg_q565 AND symb_decoder(16#86#)) OR
 					(reg_q565 AND symb_decoder(16#c8#)) OR
 					(reg_q565 AND symb_decoder(16#ee#)) OR
 					(reg_q565 AND symb_decoder(16#34#)) OR
 					(reg_q565 AND symb_decoder(16#24#)) OR
 					(reg_q565 AND symb_decoder(16#1c#)) OR
 					(reg_q565 AND symb_decoder(16#8c#)) OR
 					(reg_q565 AND symb_decoder(16#61#)) OR
 					(reg_q565 AND symb_decoder(16#13#)) OR
 					(reg_q565 AND symb_decoder(16#2e#)) OR
 					(reg_q565 AND symb_decoder(16#4f#)) OR
 					(reg_q565 AND symb_decoder(16#a6#)) OR
 					(reg_q565 AND symb_decoder(16#fb#)) OR
 					(reg_q565 AND symb_decoder(16#0e#)) OR
 					(reg_q565 AND symb_decoder(16#3b#)) OR
 					(reg_q565 AND symb_decoder(16#5d#)) OR
 					(reg_q565 AND symb_decoder(16#3f#)) OR
 					(reg_q565 AND symb_decoder(16#7e#)) OR
 					(reg_q565 AND symb_decoder(16#e8#)) OR
 					(reg_q565 AND symb_decoder(16#03#)) OR
 					(reg_q565 AND symb_decoder(16#d8#)) OR
 					(reg_q565 AND symb_decoder(16#a7#)) OR
 					(reg_q565 AND symb_decoder(16#aa#)) OR
 					(reg_q565 AND symb_decoder(16#64#)) OR
 					(reg_q565 AND symb_decoder(16#e6#)) OR
 					(reg_q565 AND symb_decoder(16#e7#)) OR
 					(reg_q565 AND symb_decoder(16#1b#)) OR
 					(reg_q565 AND symb_decoder(16#b5#)) OR
 					(reg_q565 AND symb_decoder(16#be#)) OR
 					(reg_q565 AND symb_decoder(16#c3#)) OR
 					(reg_q565 AND symb_decoder(16#e9#)) OR
 					(reg_q565 AND symb_decoder(16#bf#)) OR
 					(reg_q565 AND symb_decoder(16#82#)) OR
 					(reg_q565 AND symb_decoder(16#8e#)) OR
 					(reg_q565 AND symb_decoder(16#80#)) OR
 					(reg_q565 AND symb_decoder(16#46#)) OR
 					(reg_q565 AND symb_decoder(16#ca#)) OR
 					(reg_q565 AND symb_decoder(16#f8#)) OR
 					(reg_q565 AND symb_decoder(16#4d#)) OR
 					(reg_q565 AND symb_decoder(16#7b#)) OR
 					(reg_q565 AND symb_decoder(16#a3#)) OR
 					(reg_q565 AND symb_decoder(16#f7#)) OR
 					(reg_q565 AND symb_decoder(16#18#)) OR
 					(reg_q565 AND symb_decoder(16#72#)) OR
 					(reg_q565 AND symb_decoder(16#bd#)) OR
 					(reg_q565 AND symb_decoder(16#c5#)) OR
 					(reg_q565 AND symb_decoder(16#da#)) OR
 					(reg_q565 AND symb_decoder(16#8d#)) OR
 					(reg_q565 AND symb_decoder(16#94#)) OR
 					(reg_q565 AND symb_decoder(16#c2#)) OR
 					(reg_q565 AND symb_decoder(16#60#)) OR
 					(reg_q565 AND symb_decoder(16#3e#)) OR
 					(reg_q565 AND symb_decoder(16#06#)) OR
 					(reg_q565 AND symb_decoder(16#98#)) OR
 					(reg_q565 AND symb_decoder(16#1a#)) OR
 					(reg_q565 AND symb_decoder(16#de#)) OR
 					(reg_q565 AND symb_decoder(16#58#)) OR
 					(reg_q565 AND symb_decoder(16#50#)) OR
 					(reg_q565 AND symb_decoder(16#ce#)) OR
 					(reg_q565 AND symb_decoder(16#9a#)) OR
 					(reg_q565 AND symb_decoder(16#76#)) OR
 					(reg_q565 AND symb_decoder(16#d2#)) OR
 					(reg_q565 AND symb_decoder(16#ae#)) OR
 					(reg_q565 AND symb_decoder(16#2d#)) OR
 					(reg_q565 AND symb_decoder(16#cf#)) OR
 					(reg_q565 AND symb_decoder(16#54#)) OR
 					(reg_q565 AND symb_decoder(16#ad#)) OR
 					(reg_q565 AND symb_decoder(16#ea#)) OR
 					(reg_q565 AND symb_decoder(16#fe#)) OR
 					(reg_q565 AND symb_decoder(16#c9#)) OR
 					(reg_q565 AND symb_decoder(16#31#)) OR
 					(reg_q565 AND symb_decoder(16#2b#)) OR
 					(reg_q565 AND symb_decoder(16#6c#)) OR
 					(reg_q565 AND symb_decoder(16#19#)) OR
 					(reg_q565 AND symb_decoder(16#dd#)) OR
 					(reg_q565 AND symb_decoder(16#22#)) OR
 					(reg_q565 AND symb_decoder(16#44#)) OR
 					(reg_q565 AND symb_decoder(16#47#)) OR
 					(reg_q565 AND symb_decoder(16#b7#)) OR
 					(reg_q565 AND symb_decoder(16#3c#)) OR
 					(reg_q565 AND symb_decoder(16#ff#)) OR
 					(reg_q565 AND symb_decoder(16#93#)) OR
 					(reg_q565 AND symb_decoder(16#1e#)) OR
 					(reg_q565 AND symb_decoder(16#6f#)) OR
 					(reg_q565 AND symb_decoder(16#d4#)) OR
 					(reg_q565 AND symb_decoder(16#d7#)) OR
 					(reg_q565 AND symb_decoder(16#8b#)) OR
 					(reg_q565 AND symb_decoder(16#b1#)) OR
 					(reg_q565 AND symb_decoder(16#83#)) OR
 					(reg_q565 AND symb_decoder(16#74#)) OR
 					(reg_q565 AND symb_decoder(16#a5#)) OR
 					(reg_q565 AND symb_decoder(16#df#)) OR
 					(reg_q565 AND symb_decoder(16#11#)) OR
 					(reg_q565 AND symb_decoder(16#32#)) OR
 					(reg_q565 AND symb_decoder(16#e5#)) OR
 					(reg_q565 AND symb_decoder(16#85#)) OR
 					(reg_q565 AND symb_decoder(16#28#)) OR
 					(reg_q565 AND symb_decoder(16#65#)) OR
 					(reg_q565 AND symb_decoder(16#43#)) OR
 					(reg_q565 AND symb_decoder(16#63#)) OR
 					(reg_q565 AND symb_decoder(16#e2#)) OR
 					(reg_q565 AND symb_decoder(16#84#)) OR
 					(reg_q565 AND symb_decoder(16#55#)) OR
 					(reg_q565 AND symb_decoder(16#6a#)) OR
 					(reg_q565 AND symb_decoder(16#b2#)) OR
 					(reg_q565 AND symb_decoder(16#57#)) OR
 					(reg_q565 AND symb_decoder(16#7a#)) OR
 					(reg_q565 AND symb_decoder(16#9e#)) OR
 					(reg_q565 AND symb_decoder(16#07#)) OR
 					(reg_q565 AND symb_decoder(16#66#)) OR
 					(reg_q565 AND symb_decoder(16#af#)) OR
 					(reg_q565 AND symb_decoder(16#95#)) OR
 					(reg_q565 AND symb_decoder(16#dc#)) OR
 					(reg_q565 AND symb_decoder(16#ba#)) OR
 					(reg_q565 AND symb_decoder(16#ab#)) OR
 					(reg_q565 AND symb_decoder(16#89#)) OR
 					(reg_q565 AND symb_decoder(16#d0#)) OR
 					(reg_q565 AND symb_decoder(16#d5#)) OR
 					(reg_q565 AND symb_decoder(16#d9#)) OR
 					(reg_q565 AND symb_decoder(16#f0#)) OR
 					(reg_q565 AND symb_decoder(16#e3#)) OR
 					(reg_q565 AND symb_decoder(16#09#)) OR
 					(reg_q565 AND symb_decoder(16#69#)) OR
 					(reg_q565 AND symb_decoder(16#97#)) OR
 					(reg_q587 AND symb_decoder(16#33#)) OR
 					(reg_q587 AND symb_decoder(16#e8#)) OR
 					(reg_q587 AND symb_decoder(16#05#)) OR
 					(reg_q587 AND symb_decoder(16#d9#)) OR
 					(reg_q587 AND symb_decoder(16#8e#)) OR
 					(reg_q587 AND symb_decoder(16#be#)) OR
 					(reg_q587 AND symb_decoder(16#66#)) OR
 					(reg_q587 AND symb_decoder(16#01#)) OR
 					(reg_q587 AND symb_decoder(16#d8#)) OR
 					(reg_q587 AND symb_decoder(16#53#)) OR
 					(reg_q587 AND symb_decoder(16#7a#)) OR
 					(reg_q587 AND symb_decoder(16#1d#)) OR
 					(reg_q587 AND symb_decoder(16#2f#)) OR
 					(reg_q587 AND symb_decoder(16#5e#)) OR
 					(reg_q587 AND symb_decoder(16#7e#)) OR
 					(reg_q587 AND symb_decoder(16#9f#)) OR
 					(reg_q587 AND symb_decoder(16#06#)) OR
 					(reg_q587 AND symb_decoder(16#bc#)) OR
 					(reg_q587 AND symb_decoder(16#03#)) OR
 					(reg_q587 AND symb_decoder(16#3b#)) OR
 					(reg_q587 AND symb_decoder(16#24#)) OR
 					(reg_q587 AND symb_decoder(16#75#)) OR
 					(reg_q587 AND symb_decoder(16#7f#)) OR
 					(reg_q587 AND symb_decoder(16#91#)) OR
 					(reg_q587 AND symb_decoder(16#7b#)) OR
 					(reg_q587 AND symb_decoder(16#c7#)) OR
 					(reg_q587 AND symb_decoder(16#89#)) OR
 					(reg_q587 AND symb_decoder(16#7c#)) OR
 					(reg_q587 AND symb_decoder(16#5c#)) OR
 					(reg_q587 AND symb_decoder(16#eb#)) OR
 					(reg_q587 AND symb_decoder(16#a6#)) OR
 					(reg_q587 AND symb_decoder(16#6e#)) OR
 					(reg_q587 AND symb_decoder(16#84#)) OR
 					(reg_q587 AND symb_decoder(16#d0#)) OR
 					(reg_q587 AND symb_decoder(16#9c#)) OR
 					(reg_q587 AND symb_decoder(16#04#)) OR
 					(reg_q587 AND symb_decoder(16#1f#)) OR
 					(reg_q587 AND symb_decoder(16#de#)) OR
 					(reg_q587 AND symb_decoder(16#6f#)) OR
 					(reg_q587 AND symb_decoder(16#b1#)) OR
 					(reg_q587 AND symb_decoder(16#2a#)) OR
 					(reg_q587 AND symb_decoder(16#72#)) OR
 					(reg_q587 AND symb_decoder(16#21#)) OR
 					(reg_q587 AND symb_decoder(16#23#)) OR
 					(reg_q587 AND symb_decoder(16#62#)) OR
 					(reg_q587 AND symb_decoder(16#74#)) OR
 					(reg_q587 AND symb_decoder(16#48#)) OR
 					(reg_q587 AND symb_decoder(16#49#)) OR
 					(reg_q587 AND symb_decoder(16#13#)) OR
 					(reg_q587 AND symb_decoder(16#cf#)) OR
 					(reg_q587 AND symb_decoder(16#4e#)) OR
 					(reg_q587 AND symb_decoder(16#82#)) OR
 					(reg_q587 AND symb_decoder(16#16#)) OR
 					(reg_q587 AND symb_decoder(16#f7#)) OR
 					(reg_q587 AND symb_decoder(16#67#)) OR
 					(reg_q587 AND symb_decoder(16#00#)) OR
 					(reg_q587 AND symb_decoder(16#d1#)) OR
 					(reg_q587 AND symb_decoder(16#0c#)) OR
 					(reg_q587 AND symb_decoder(16#d6#)) OR
 					(reg_q587 AND symb_decoder(16#52#)) OR
 					(reg_q587 AND symb_decoder(16#57#)) OR
 					(reg_q587 AND symb_decoder(16#f6#)) OR
 					(reg_q587 AND symb_decoder(16#71#)) OR
 					(reg_q587 AND symb_decoder(16#bb#)) OR
 					(reg_q587 AND symb_decoder(16#ef#)) OR
 					(reg_q587 AND symb_decoder(16#4b#)) OR
 					(reg_q587 AND symb_decoder(16#e5#)) OR
 					(reg_q587 AND symb_decoder(16#96#)) OR
 					(reg_q587 AND symb_decoder(16#f8#)) OR
 					(reg_q587 AND symb_decoder(16#fa#)) OR
 					(reg_q587 AND symb_decoder(16#fd#)) OR
 					(reg_q587 AND symb_decoder(16#fc#)) OR
 					(reg_q587 AND symb_decoder(16#5d#)) OR
 					(reg_q587 AND symb_decoder(16#4f#)) OR
 					(reg_q587 AND symb_decoder(16#b4#)) OR
 					(reg_q587 AND symb_decoder(16#47#)) OR
 					(reg_q587 AND symb_decoder(16#02#)) OR
 					(reg_q587 AND symb_decoder(16#5a#)) OR
 					(reg_q587 AND symb_decoder(16#d4#)) OR
 					(reg_q587 AND symb_decoder(16#e3#)) OR
 					(reg_q587 AND symb_decoder(16#8c#)) OR
 					(reg_q587 AND symb_decoder(16#7d#)) OR
 					(reg_q587 AND symb_decoder(16#f2#)) OR
 					(reg_q587 AND symb_decoder(16#46#)) OR
 					(reg_q587 AND symb_decoder(16#29#)) OR
 					(reg_q587 AND symb_decoder(16#45#)) OR
 					(reg_q587 AND symb_decoder(16#97#)) OR
 					(reg_q587 AND symb_decoder(16#63#)) OR
 					(reg_q587 AND symb_decoder(16#37#)) OR
 					(reg_q587 AND symb_decoder(16#cd#)) OR
 					(reg_q587 AND symb_decoder(16#54#)) OR
 					(reg_q587 AND symb_decoder(16#f3#)) OR
 					(reg_q587 AND symb_decoder(16#36#)) OR
 					(reg_q587 AND symb_decoder(16#56#)) OR
 					(reg_q587 AND symb_decoder(16#ae#)) OR
 					(reg_q587 AND symb_decoder(16#b8#)) OR
 					(reg_q587 AND symb_decoder(16#f0#)) OR
 					(reg_q587 AND symb_decoder(16#77#)) OR
 					(reg_q587 AND symb_decoder(16#ba#)) OR
 					(reg_q587 AND symb_decoder(16#78#)) OR
 					(reg_q587 AND symb_decoder(16#e6#)) OR
 					(reg_q587 AND symb_decoder(16#e0#)) OR
 					(reg_q587 AND symb_decoder(16#ac#)) OR
 					(reg_q587 AND symb_decoder(16#ee#)) OR
 					(reg_q587 AND symb_decoder(16#ff#)) OR
 					(reg_q587 AND symb_decoder(16#e2#)) OR
 					(reg_q587 AND symb_decoder(16#4a#)) OR
 					(reg_q587 AND symb_decoder(16#e7#)) OR
 					(reg_q587 AND symb_decoder(16#a3#)) OR
 					(reg_q587 AND symb_decoder(16#10#)) OR
 					(reg_q587 AND symb_decoder(16#c6#)) OR
 					(reg_q587 AND symb_decoder(16#85#)) OR
 					(reg_q587 AND symb_decoder(16#88#)) OR
 					(reg_q587 AND symb_decoder(16#07#)) OR
 					(reg_q587 AND symb_decoder(16#80#)) OR
 					(reg_q587 AND symb_decoder(16#61#)) OR
 					(reg_q587 AND symb_decoder(16#ec#)) OR
 					(reg_q587 AND symb_decoder(16#c4#)) OR
 					(reg_q587 AND symb_decoder(16#fb#)) OR
 					(reg_q587 AND symb_decoder(16#ab#)) OR
 					(reg_q587 AND symb_decoder(16#76#)) OR
 					(reg_q587 AND symb_decoder(16#3f#)) OR
 					(reg_q587 AND symb_decoder(16#ed#)) OR
 					(reg_q587 AND symb_decoder(16#db#)) OR
 					(reg_q587 AND symb_decoder(16#14#)) OR
 					(reg_q587 AND symb_decoder(16#9e#)) OR
 					(reg_q587 AND symb_decoder(16#73#)) OR
 					(reg_q587 AND symb_decoder(16#50#)) OR
 					(reg_q587 AND symb_decoder(16#42#)) OR
 					(reg_q587 AND symb_decoder(16#3e#)) OR
 					(reg_q587 AND symb_decoder(16#79#)) OR
 					(reg_q587 AND symb_decoder(16#55#)) OR
 					(reg_q587 AND symb_decoder(16#41#)) OR
 					(reg_q587 AND symb_decoder(16#3d#)) OR
 					(reg_q587 AND symb_decoder(16#b6#)) OR
 					(reg_q587 AND symb_decoder(16#c1#)) OR
 					(reg_q587 AND symb_decoder(16#0e#)) OR
 					(reg_q587 AND symb_decoder(16#f4#)) OR
 					(reg_q587 AND symb_decoder(16#df#)) OR
 					(reg_q587 AND symb_decoder(16#a5#)) OR
 					(reg_q587 AND symb_decoder(16#3a#)) OR
 					(reg_q587 AND symb_decoder(16#60#)) OR
 					(reg_q587 AND symb_decoder(16#8f#)) OR
 					(reg_q587 AND symb_decoder(16#59#)) OR
 					(reg_q587 AND symb_decoder(16#30#)) OR
 					(reg_q587 AND symb_decoder(16#d5#)) OR
 					(reg_q587 AND symb_decoder(16#08#)) OR
 					(reg_q587 AND symb_decoder(16#99#)) OR
 					(reg_q587 AND symb_decoder(16#3c#)) OR
 					(reg_q587 AND symb_decoder(16#20#)) OR
 					(reg_q587 AND symb_decoder(16#ca#)) OR
 					(reg_q587 AND symb_decoder(16#e1#)) OR
 					(reg_q587 AND symb_decoder(16#d2#)) OR
 					(reg_q587 AND symb_decoder(16#e9#)) OR
 					(reg_q587 AND symb_decoder(16#6b#)) OR
 					(reg_q587 AND symb_decoder(16#86#)) OR
 					(reg_q587 AND symb_decoder(16#ad#)) OR
 					(reg_q587 AND symb_decoder(16#c0#)) OR
 					(reg_q587 AND symb_decoder(16#b5#)) OR
 					(reg_q587 AND symb_decoder(16#ea#)) OR
 					(reg_q587 AND symb_decoder(16#c2#)) OR
 					(reg_q587 AND symb_decoder(16#64#)) OR
 					(reg_q587 AND symb_decoder(16#32#)) OR
 					(reg_q587 AND symb_decoder(16#51#)) OR
 					(reg_q587 AND symb_decoder(16#ce#)) OR
 					(reg_q587 AND symb_decoder(16#bd#)) OR
 					(reg_q587 AND symb_decoder(16#68#)) OR
 					(reg_q587 AND symb_decoder(16#6d#)) OR
 					(reg_q587 AND symb_decoder(16#e4#)) OR
 					(reg_q587 AND symb_decoder(16#2c#)) OR
 					(reg_q587 AND symb_decoder(16#2b#)) OR
 					(reg_q587 AND symb_decoder(16#a7#)) OR
 					(reg_q587 AND symb_decoder(16#2d#)) OR
 					(reg_q587 AND symb_decoder(16#17#)) OR
 					(reg_q587 AND symb_decoder(16#70#)) OR
 					(reg_q587 AND symb_decoder(16#f9#)) OR
 					(reg_q587 AND symb_decoder(16#a8#)) OR
 					(reg_q587 AND symb_decoder(16#34#)) OR
 					(reg_q587 AND symb_decoder(16#27#)) OR
 					(reg_q587 AND symb_decoder(16#98#)) OR
 					(reg_q587 AND symb_decoder(16#15#)) OR
 					(reg_q587 AND symb_decoder(16#fe#)) OR
 					(reg_q587 AND symb_decoder(16#18#)) OR
 					(reg_q587 AND symb_decoder(16#8d#)) OR
 					(reg_q587 AND symb_decoder(16#81#)) OR
 					(reg_q587 AND symb_decoder(16#cb#)) OR
 					(reg_q587 AND symb_decoder(16#83#)) OR
 					(reg_q587 AND symb_decoder(16#af#)) OR
 					(reg_q587 AND symb_decoder(16#4d#)) OR
 					(reg_q587 AND symb_decoder(16#c9#)) OR
 					(reg_q587 AND symb_decoder(16#5f#)) OR
 					(reg_q587 AND symb_decoder(16#c5#)) OR
 					(reg_q587 AND symb_decoder(16#c8#)) OR
 					(reg_q587 AND symb_decoder(16#8a#)) OR
 					(reg_q587 AND symb_decoder(16#9b#)) OR
 					(reg_q587 AND symb_decoder(16#90#)) OR
 					(reg_q587 AND symb_decoder(16#a1#)) OR
 					(reg_q587 AND symb_decoder(16#da#)) OR
 					(reg_q587 AND symb_decoder(16#9a#)) OR
 					(reg_q587 AND symb_decoder(16#2e#)) OR
 					(reg_q587 AND symb_decoder(16#94#)) OR
 					(reg_q587 AND symb_decoder(16#a2#)) OR
 					(reg_q587 AND symb_decoder(16#44#)) OR
 					(reg_q587 AND symb_decoder(16#d7#)) OR
 					(reg_q587 AND symb_decoder(16#40#)) OR
 					(reg_q587 AND symb_decoder(16#0f#)) OR
 					(reg_q587 AND symb_decoder(16#1e#)) OR
 					(reg_q587 AND symb_decoder(16#92#)) OR
 					(reg_q587 AND symb_decoder(16#bf#)) OR
 					(reg_q587 AND symb_decoder(16#11#)) OR
 					(reg_q587 AND symb_decoder(16#4c#)) OR
 					(reg_q587 AND symb_decoder(16#cc#)) OR
 					(reg_q587 AND symb_decoder(16#19#)) OR
 					(reg_q587 AND symb_decoder(16#f1#)) OR
 					(reg_q587 AND symb_decoder(16#31#)) OR
 					(reg_q587 AND symb_decoder(16#b7#)) OR
 					(reg_q587 AND symb_decoder(16#6c#)) OR
 					(reg_q587 AND symb_decoder(16#93#)) OR
 					(reg_q587 AND symb_decoder(16#26#)) OR
 					(reg_q587 AND symb_decoder(16#69#)) OR
 					(reg_q587 AND symb_decoder(16#b3#)) OR
 					(reg_q587 AND symb_decoder(16#c3#)) OR
 					(reg_q587 AND symb_decoder(16#87#)) OR
 					(reg_q587 AND symb_decoder(16#25#)) OR
 					(reg_q587 AND symb_decoder(16#35#)) OR
 					(reg_q587 AND symb_decoder(16#43#)) OR
 					(reg_q587 AND symb_decoder(16#b0#)) OR
 					(reg_q587 AND symb_decoder(16#1c#)) OR
 					(reg_q587 AND symb_decoder(16#f5#)) OR
 					(reg_q587 AND symb_decoder(16#65#)) OR
 					(reg_q587 AND symb_decoder(16#8b#)) OR
 					(reg_q587 AND symb_decoder(16#5b#)) OR
 					(reg_q587 AND symb_decoder(16#b2#)) OR
 					(reg_q587 AND symb_decoder(16#38#)) OR
 					(reg_q587 AND symb_decoder(16#12#)) OR
 					(reg_q587 AND symb_decoder(16#28#)) OR
 					(reg_q587 AND symb_decoder(16#95#)) OR
 					(reg_q587 AND symb_decoder(16#1b#)) OR
 					(reg_q587 AND symb_decoder(16#b9#)) OR
 					(reg_q587 AND symb_decoder(16#dc#)) OR
 					(reg_q587 AND symb_decoder(16#dd#)) OR
 					(reg_q587 AND symb_decoder(16#9d#)) OR
 					(reg_q587 AND symb_decoder(16#1a#)) OR
 					(reg_q587 AND symb_decoder(16#58#)) OR
 					(reg_q587 AND symb_decoder(16#09#)) OR
 					(reg_q587 AND symb_decoder(16#0b#)) OR
 					(reg_q587 AND symb_decoder(16#22#)) OR
 					(reg_q587 AND symb_decoder(16#a4#)) OR
 					(reg_q587 AND symb_decoder(16#aa#)) OR
 					(reg_q587 AND symb_decoder(16#39#)) OR
 					(reg_q587 AND symb_decoder(16#a0#)) OR
 					(reg_q587 AND symb_decoder(16#6a#)) OR
 					(reg_q587 AND symb_decoder(16#a9#)) OR
 					(reg_q587 AND symb_decoder(16#d3#));
reg_q1323_in <= (reg_q1323 AND symb_decoder(16#0a#)) OR
 					(reg_q1323 AND symb_decoder(16#0c#)) OR
 					(reg_q1323 AND symb_decoder(16#09#)) OR
 					(reg_q1323 AND symb_decoder(16#0d#)) OR
 					(reg_q1323 AND symb_decoder(16#20#)) OR
 					(reg_q1321 AND symb_decoder(16#0a#)) OR
 					(reg_q1321 AND symb_decoder(16#0c#)) OR
 					(reg_q1321 AND symb_decoder(16#0d#)) OR
 					(reg_q1321 AND symb_decoder(16#09#)) OR
 					(reg_q1321 AND symb_decoder(16#20#));
reg_q494_in <= (reg_q494 AND symb_decoder(16#b1#)) OR
 					(reg_q494 AND symb_decoder(16#63#)) OR
 					(reg_q494 AND symb_decoder(16#93#)) OR
 					(reg_q494 AND symb_decoder(16#15#)) OR
 					(reg_q494 AND symb_decoder(16#d5#)) OR
 					(reg_q494 AND symb_decoder(16#9a#)) OR
 					(reg_q494 AND symb_decoder(16#ef#)) OR
 					(reg_q494 AND symb_decoder(16#4c#)) OR
 					(reg_q494 AND symb_decoder(16#aa#)) OR
 					(reg_q494 AND symb_decoder(16#50#)) OR
 					(reg_q494 AND symb_decoder(16#fc#)) OR
 					(reg_q494 AND symb_decoder(16#a5#)) OR
 					(reg_q494 AND symb_decoder(16#75#)) OR
 					(reg_q494 AND symb_decoder(16#24#)) OR
 					(reg_q494 AND symb_decoder(16#37#)) OR
 					(reg_q494 AND symb_decoder(16#06#)) OR
 					(reg_q494 AND symb_decoder(16#3e#)) OR
 					(reg_q494 AND symb_decoder(16#a4#)) OR
 					(reg_q494 AND symb_decoder(16#e7#)) OR
 					(reg_q494 AND symb_decoder(16#8b#)) OR
 					(reg_q494 AND symb_decoder(16#0e#)) OR
 					(reg_q494 AND symb_decoder(16#86#)) OR
 					(reg_q494 AND symb_decoder(16#04#)) OR
 					(reg_q494 AND symb_decoder(16#5d#)) OR
 					(reg_q494 AND symb_decoder(16#84#)) OR
 					(reg_q494 AND symb_decoder(16#a7#)) OR
 					(reg_q494 AND symb_decoder(16#30#)) OR
 					(reg_q494 AND symb_decoder(16#d4#)) OR
 					(reg_q494 AND symb_decoder(16#ee#)) OR
 					(reg_q494 AND symb_decoder(16#5b#)) OR
 					(reg_q494 AND symb_decoder(16#d6#)) OR
 					(reg_q494 AND symb_decoder(16#f5#)) OR
 					(reg_q494 AND symb_decoder(16#a6#)) OR
 					(reg_q494 AND symb_decoder(16#f7#)) OR
 					(reg_q494 AND symb_decoder(16#cc#)) OR
 					(reg_q494 AND symb_decoder(16#79#)) OR
 					(reg_q494 AND symb_decoder(16#23#)) OR
 					(reg_q494 AND symb_decoder(16#45#)) OR
 					(reg_q494 AND symb_decoder(16#5f#)) OR
 					(reg_q494 AND symb_decoder(16#7d#)) OR
 					(reg_q494 AND symb_decoder(16#02#)) OR
 					(reg_q494 AND symb_decoder(16#dd#)) OR
 					(reg_q494 AND symb_decoder(16#71#)) OR
 					(reg_q494 AND symb_decoder(16#19#)) OR
 					(reg_q494 AND symb_decoder(16#ab#)) OR
 					(reg_q494 AND symb_decoder(16#ac#)) OR
 					(reg_q494 AND symb_decoder(16#44#)) OR
 					(reg_q494 AND symb_decoder(16#08#)) OR
 					(reg_q494 AND symb_decoder(16#c9#)) OR
 					(reg_q494 AND symb_decoder(16#1b#)) OR
 					(reg_q494 AND symb_decoder(16#01#)) OR
 					(reg_q494 AND symb_decoder(16#33#)) OR
 					(reg_q494 AND symb_decoder(16#03#)) OR
 					(reg_q494 AND symb_decoder(16#d9#)) OR
 					(reg_q494 AND symb_decoder(16#0c#)) OR
 					(reg_q494 AND symb_decoder(16#e8#)) OR
 					(reg_q494 AND symb_decoder(16#95#)) OR
 					(reg_q494 AND symb_decoder(16#14#)) OR
 					(reg_q494 AND symb_decoder(16#12#)) OR
 					(reg_q494 AND symb_decoder(16#e3#)) OR
 					(reg_q494 AND symb_decoder(16#29#)) OR
 					(reg_q494 AND symb_decoder(16#cf#)) OR
 					(reg_q494 AND symb_decoder(16#16#)) OR
 					(reg_q494 AND symb_decoder(16#c4#)) OR
 					(reg_q494 AND symb_decoder(16#ca#)) OR
 					(reg_q494 AND symb_decoder(16#90#)) OR
 					(reg_q494 AND symb_decoder(16#f0#)) OR
 					(reg_q494 AND symb_decoder(16#9c#)) OR
 					(reg_q494 AND symb_decoder(16#76#)) OR
 					(reg_q494 AND symb_decoder(16#f8#)) OR
 					(reg_q494 AND symb_decoder(16#db#)) OR
 					(reg_q494 AND symb_decoder(16#da#)) OR
 					(reg_q494 AND symb_decoder(16#9e#)) OR
 					(reg_q494 AND symb_decoder(16#64#)) OR
 					(reg_q494 AND symb_decoder(16#59#)) OR
 					(reg_q494 AND symb_decoder(16#a9#)) OR
 					(reg_q494 AND symb_decoder(16#87#)) OR
 					(reg_q494 AND symb_decoder(16#ed#)) OR
 					(reg_q494 AND symb_decoder(16#e2#)) OR
 					(reg_q494 AND symb_decoder(16#09#)) OR
 					(reg_q494 AND symb_decoder(16#2f#)) OR
 					(reg_q494 AND symb_decoder(16#d3#)) OR
 					(reg_q494 AND symb_decoder(16#49#)) OR
 					(reg_q494 AND symb_decoder(16#ea#)) OR
 					(reg_q494 AND symb_decoder(16#47#)) OR
 					(reg_q494 AND symb_decoder(16#a3#)) OR
 					(reg_q494 AND symb_decoder(16#55#)) OR
 					(reg_q494 AND symb_decoder(16#af#)) OR
 					(reg_q494 AND symb_decoder(16#c0#)) OR
 					(reg_q494 AND symb_decoder(16#ce#)) OR
 					(reg_q494 AND symb_decoder(16#a0#)) OR
 					(reg_q494 AND symb_decoder(16#2c#)) OR
 					(reg_q494 AND symb_decoder(16#7f#)) OR
 					(reg_q494 AND symb_decoder(16#77#)) OR
 					(reg_q494 AND symb_decoder(16#74#)) OR
 					(reg_q494 AND symb_decoder(16#2a#)) OR
 					(reg_q494 AND symb_decoder(16#66#)) OR
 					(reg_q494 AND symb_decoder(16#70#)) OR
 					(reg_q494 AND symb_decoder(16#69#)) OR
 					(reg_q494 AND symb_decoder(16#9d#)) OR
 					(reg_q494 AND symb_decoder(16#32#)) OR
 					(reg_q494 AND symb_decoder(16#b5#)) OR
 					(reg_q494 AND symb_decoder(16#96#)) OR
 					(reg_q494 AND symb_decoder(16#f2#)) OR
 					(reg_q494 AND symb_decoder(16#10#)) OR
 					(reg_q494 AND symb_decoder(16#bf#)) OR
 					(reg_q494 AND symb_decoder(16#83#)) OR
 					(reg_q494 AND symb_decoder(16#e4#)) OR
 					(reg_q494 AND symb_decoder(16#3d#)) OR
 					(reg_q494 AND symb_decoder(16#17#)) OR
 					(reg_q494 AND symb_decoder(16#ff#)) OR
 					(reg_q494 AND symb_decoder(16#3b#)) OR
 					(reg_q494 AND symb_decoder(16#73#)) OR
 					(reg_q494 AND symb_decoder(16#f6#)) OR
 					(reg_q494 AND symb_decoder(16#7b#)) OR
 					(reg_q494 AND symb_decoder(16#4e#)) OR
 					(reg_q494 AND symb_decoder(16#3a#)) OR
 					(reg_q494 AND symb_decoder(16#9f#)) OR
 					(reg_q494 AND symb_decoder(16#e0#)) OR
 					(reg_q494 AND symb_decoder(16#1e#)) OR
 					(reg_q494 AND symb_decoder(16#c3#)) OR
 					(reg_q494 AND symb_decoder(16#57#)) OR
 					(reg_q494 AND symb_decoder(16#b6#)) OR
 					(reg_q494 AND symb_decoder(16#11#)) OR
 					(reg_q494 AND symb_decoder(16#c2#)) OR
 					(reg_q494 AND symb_decoder(16#d0#)) OR
 					(reg_q494 AND symb_decoder(16#3f#)) OR
 					(reg_q494 AND symb_decoder(16#67#)) OR
 					(reg_q494 AND symb_decoder(16#4d#)) OR
 					(reg_q494 AND symb_decoder(16#4b#)) OR
 					(reg_q494 AND symb_decoder(16#e5#)) OR
 					(reg_q494 AND symb_decoder(16#ad#)) OR
 					(reg_q494 AND symb_decoder(16#cd#)) OR
 					(reg_q494 AND symb_decoder(16#bd#)) OR
 					(reg_q494 AND symb_decoder(16#3c#)) OR
 					(reg_q494 AND symb_decoder(16#d2#)) OR
 					(reg_q494 AND symb_decoder(16#18#)) OR
 					(reg_q494 AND symb_decoder(16#42#)) OR
 					(reg_q494 AND symb_decoder(16#7a#)) OR
 					(reg_q494 AND symb_decoder(16#89#)) OR
 					(reg_q494 AND symb_decoder(16#a8#)) OR
 					(reg_q494 AND symb_decoder(16#38#)) OR
 					(reg_q494 AND symb_decoder(16#41#)) OR
 					(reg_q494 AND symb_decoder(16#35#)) OR
 					(reg_q494 AND symb_decoder(16#40#)) OR
 					(reg_q494 AND symb_decoder(16#e6#)) OR
 					(reg_q494 AND symb_decoder(16#eb#)) OR
 					(reg_q494 AND symb_decoder(16#88#)) OR
 					(reg_q494 AND symb_decoder(16#5e#)) OR
 					(reg_q494 AND symb_decoder(16#6d#)) OR
 					(reg_q494 AND symb_decoder(16#c6#)) OR
 					(reg_q494 AND symb_decoder(16#d1#)) OR
 					(reg_q494 AND symb_decoder(16#62#)) OR
 					(reg_q494 AND symb_decoder(16#b9#)) OR
 					(reg_q494 AND symb_decoder(16#1c#)) OR
 					(reg_q494 AND symb_decoder(16#0f#)) OR
 					(reg_q494 AND symb_decoder(16#58#)) OR
 					(reg_q494 AND symb_decoder(16#28#)) OR
 					(reg_q494 AND symb_decoder(16#80#)) OR
 					(reg_q494 AND symb_decoder(16#dc#)) OR
 					(reg_q494 AND symb_decoder(16#ae#)) OR
 					(reg_q494 AND symb_decoder(16#c5#)) OR
 					(reg_q494 AND symb_decoder(16#97#)) OR
 					(reg_q494 AND symb_decoder(16#e9#)) OR
 					(reg_q494 AND symb_decoder(16#22#)) OR
 					(reg_q494 AND symb_decoder(16#fb#)) OR
 					(reg_q494 AND symb_decoder(16#52#)) OR
 					(reg_q494 AND symb_decoder(16#b8#)) OR
 					(reg_q494 AND symb_decoder(16#de#)) OR
 					(reg_q494 AND symb_decoder(16#20#)) OR
 					(reg_q494 AND symb_decoder(16#fd#)) OR
 					(reg_q494 AND symb_decoder(16#99#)) OR
 					(reg_q494 AND symb_decoder(16#f3#)) OR
 					(reg_q494 AND symb_decoder(16#a1#)) OR
 					(reg_q494 AND symb_decoder(16#b7#)) OR
 					(reg_q494 AND symb_decoder(16#6e#)) OR
 					(reg_q494 AND symb_decoder(16#46#)) OR
 					(reg_q494 AND symb_decoder(16#60#)) OR
 					(reg_q494 AND symb_decoder(16#be#)) OR
 					(reg_q494 AND symb_decoder(16#07#)) OR
 					(reg_q494 AND symb_decoder(16#2b#)) OR
 					(reg_q494 AND symb_decoder(16#b2#)) OR
 					(reg_q494 AND symb_decoder(16#5a#)) OR
 					(reg_q494 AND symb_decoder(16#8a#)) OR
 					(reg_q494 AND symb_decoder(16#8e#)) OR
 					(reg_q494 AND symb_decoder(16#05#)) OR
 					(reg_q494 AND symb_decoder(16#d8#)) OR
 					(reg_q494 AND symb_decoder(16#bc#)) OR
 					(reg_q494 AND symb_decoder(16#98#)) OR
 					(reg_q494 AND symb_decoder(16#8f#)) OR
 					(reg_q494 AND symb_decoder(16#b3#)) OR
 					(reg_q494 AND symb_decoder(16#82#)) OR
 					(reg_q494 AND symb_decoder(16#c8#)) OR
 					(reg_q494 AND symb_decoder(16#25#)) OR
 					(reg_q494 AND symb_decoder(16#72#)) OR
 					(reg_q494 AND symb_decoder(16#d7#)) OR
 					(reg_q494 AND symb_decoder(16#6a#)) OR
 					(reg_q494 AND symb_decoder(16#61#)) OR
 					(reg_q494 AND symb_decoder(16#21#)) OR
 					(reg_q494 AND symb_decoder(16#df#)) OR
 					(reg_q494 AND symb_decoder(16#92#)) OR
 					(reg_q494 AND symb_decoder(16#e1#)) OR
 					(reg_q494 AND symb_decoder(16#27#)) OR
 					(reg_q494 AND symb_decoder(16#1d#)) OR
 					(reg_q494 AND symb_decoder(16#94#)) OR
 					(reg_q494 AND symb_decoder(16#7c#)) OR
 					(reg_q494 AND symb_decoder(16#f4#)) OR
 					(reg_q494 AND symb_decoder(16#b4#)) OR
 					(reg_q494 AND symb_decoder(16#85#)) OR
 					(reg_q494 AND symb_decoder(16#5c#)) OR
 					(reg_q494 AND symb_decoder(16#c7#)) OR
 					(reg_q494 AND symb_decoder(16#48#)) OR
 					(reg_q494 AND symb_decoder(16#53#)) OR
 					(reg_q494 AND symb_decoder(16#0b#)) OR
 					(reg_q494 AND symb_decoder(16#f9#)) OR
 					(reg_q494 AND symb_decoder(16#65#)) OR
 					(reg_q494 AND symb_decoder(16#1f#)) OR
 					(reg_q494 AND symb_decoder(16#fe#)) OR
 					(reg_q494 AND symb_decoder(16#81#)) OR
 					(reg_q494 AND symb_decoder(16#f1#)) OR
 					(reg_q494 AND symb_decoder(16#ba#)) OR
 					(reg_q494 AND symb_decoder(16#cb#)) OR
 					(reg_q494 AND symb_decoder(16#78#)) OR
 					(reg_q494 AND symb_decoder(16#8d#)) OR
 					(reg_q494 AND symb_decoder(16#2e#)) OR
 					(reg_q494 AND symb_decoder(16#c1#)) OR
 					(reg_q494 AND symb_decoder(16#6b#)) OR
 					(reg_q494 AND symb_decoder(16#4f#)) OR
 					(reg_q494 AND symb_decoder(16#fa#)) OR
 					(reg_q494 AND symb_decoder(16#8c#)) OR
 					(reg_q494 AND symb_decoder(16#43#)) OR
 					(reg_q494 AND symb_decoder(16#a2#)) OR
 					(reg_q494 AND symb_decoder(16#68#)) OR
 					(reg_q494 AND symb_decoder(16#34#)) OR
 					(reg_q494 AND symb_decoder(16#2d#)) OR
 					(reg_q494 AND symb_decoder(16#ec#)) OR
 					(reg_q494 AND symb_decoder(16#91#)) OR
 					(reg_q494 AND symb_decoder(16#13#)) OR
 					(reg_q494 AND symb_decoder(16#36#)) OR
 					(reg_q494 AND symb_decoder(16#4a#)) OR
 					(reg_q494 AND symb_decoder(16#31#)) OR
 					(reg_q494 AND symb_decoder(16#00#)) OR
 					(reg_q494 AND symb_decoder(16#54#)) OR
 					(reg_q494 AND symb_decoder(16#9b#)) OR
 					(reg_q494 AND symb_decoder(16#56#)) OR
 					(reg_q494 AND symb_decoder(16#1a#)) OR
 					(reg_q494 AND symb_decoder(16#26#)) OR
 					(reg_q494 AND symb_decoder(16#6c#)) OR
 					(reg_q494 AND symb_decoder(16#39#)) OR
 					(reg_q494 AND symb_decoder(16#7e#)) OR
 					(reg_q494 AND symb_decoder(16#bb#)) OR
 					(reg_q494 AND symb_decoder(16#6f#)) OR
 					(reg_q494 AND symb_decoder(16#51#)) OR
 					(reg_q494 AND symb_decoder(16#b0#)) OR
 					(reg_q480 AND symb_decoder(16#5e#)) OR
 					(reg_q480 AND symb_decoder(16#9d#)) OR
 					(reg_q480 AND symb_decoder(16#10#)) OR
 					(reg_q480 AND symb_decoder(16#ec#)) OR
 					(reg_q480 AND symb_decoder(16#f8#)) OR
 					(reg_q480 AND symb_decoder(16#94#)) OR
 					(reg_q480 AND symb_decoder(16#18#)) OR
 					(reg_q480 AND symb_decoder(16#ad#)) OR
 					(reg_q480 AND symb_decoder(16#2b#)) OR
 					(reg_q480 AND symb_decoder(16#ee#)) OR
 					(reg_q480 AND symb_decoder(16#66#)) OR
 					(reg_q480 AND symb_decoder(16#c0#)) OR
 					(reg_q480 AND symb_decoder(16#2d#)) OR
 					(reg_q480 AND symb_decoder(16#01#)) OR
 					(reg_q480 AND symb_decoder(16#8a#)) OR
 					(reg_q480 AND symb_decoder(16#8f#)) OR
 					(reg_q480 AND symb_decoder(16#6a#)) OR
 					(reg_q480 AND symb_decoder(16#eb#)) OR
 					(reg_q480 AND symb_decoder(16#73#)) OR
 					(reg_q480 AND symb_decoder(16#9b#)) OR
 					(reg_q480 AND symb_decoder(16#ff#)) OR
 					(reg_q480 AND symb_decoder(16#82#)) OR
 					(reg_q480 AND symb_decoder(16#6b#)) OR
 					(reg_q480 AND symb_decoder(16#55#)) OR
 					(reg_q480 AND symb_decoder(16#a6#)) OR
 					(reg_q480 AND symb_decoder(16#3a#)) OR
 					(reg_q480 AND symb_decoder(16#ea#)) OR
 					(reg_q480 AND symb_decoder(16#72#)) OR
 					(reg_q480 AND symb_decoder(16#44#)) OR
 					(reg_q480 AND symb_decoder(16#fa#)) OR
 					(reg_q480 AND symb_decoder(16#b4#)) OR
 					(reg_q480 AND symb_decoder(16#e6#)) OR
 					(reg_q480 AND symb_decoder(16#61#)) OR
 					(reg_q480 AND symb_decoder(16#ce#)) OR
 					(reg_q480 AND symb_decoder(16#42#)) OR
 					(reg_q480 AND symb_decoder(16#5c#)) OR
 					(reg_q480 AND symb_decoder(16#d8#)) OR
 					(reg_q480 AND symb_decoder(16#b1#)) OR
 					(reg_q480 AND symb_decoder(16#bc#)) OR
 					(reg_q480 AND symb_decoder(16#84#)) OR
 					(reg_q480 AND symb_decoder(16#d5#)) OR
 					(reg_q480 AND symb_decoder(16#d1#)) OR
 					(reg_q480 AND symb_decoder(16#60#)) OR
 					(reg_q480 AND symb_decoder(16#58#)) OR
 					(reg_q480 AND symb_decoder(16#2f#)) OR
 					(reg_q480 AND symb_decoder(16#c2#)) OR
 					(reg_q480 AND symb_decoder(16#c8#)) OR
 					(reg_q480 AND symb_decoder(16#6e#)) OR
 					(reg_q480 AND symb_decoder(16#76#)) OR
 					(reg_q480 AND symb_decoder(16#d2#)) OR
 					(reg_q480 AND symb_decoder(16#77#)) OR
 					(reg_q480 AND symb_decoder(16#4d#)) OR
 					(reg_q480 AND symb_decoder(16#51#)) OR
 					(reg_q480 AND symb_decoder(16#81#)) OR
 					(reg_q480 AND symb_decoder(16#e2#)) OR
 					(reg_q480 AND symb_decoder(16#da#)) OR
 					(reg_q480 AND symb_decoder(16#80#)) OR
 					(reg_q480 AND symb_decoder(16#e8#)) OR
 					(reg_q480 AND symb_decoder(16#33#)) OR
 					(reg_q480 AND symb_decoder(16#46#)) OR
 					(reg_q480 AND symb_decoder(16#6f#)) OR
 					(reg_q480 AND symb_decoder(16#27#)) OR
 					(reg_q480 AND symb_decoder(16#45#)) OR
 					(reg_q480 AND symb_decoder(16#dc#)) OR
 					(reg_q480 AND symb_decoder(16#59#)) OR
 					(reg_q480 AND symb_decoder(16#40#)) OR
 					(reg_q480 AND symb_decoder(16#d0#)) OR
 					(reg_q480 AND symb_decoder(16#39#)) OR
 					(reg_q480 AND symb_decoder(16#08#)) OR
 					(reg_q480 AND symb_decoder(16#4f#)) OR
 					(reg_q480 AND symb_decoder(16#86#)) OR
 					(reg_q480 AND symb_decoder(16#67#)) OR
 					(reg_q480 AND symb_decoder(16#ed#)) OR
 					(reg_q480 AND symb_decoder(16#8b#)) OR
 					(reg_q480 AND symb_decoder(16#65#)) OR
 					(reg_q480 AND symb_decoder(16#a5#)) OR
 					(reg_q480 AND symb_decoder(16#35#)) OR
 					(reg_q480 AND symb_decoder(16#69#)) OR
 					(reg_q480 AND symb_decoder(16#3f#)) OR
 					(reg_q480 AND symb_decoder(16#b3#)) OR
 					(reg_q480 AND symb_decoder(16#07#)) OR
 					(reg_q480 AND symb_decoder(16#24#)) OR
 					(reg_q480 AND symb_decoder(16#70#)) OR
 					(reg_q480 AND symb_decoder(16#dd#)) OR
 					(reg_q480 AND symb_decoder(16#16#)) OR
 					(reg_q480 AND symb_decoder(16#0f#)) OR
 					(reg_q480 AND symb_decoder(16#96#)) OR
 					(reg_q480 AND symb_decoder(16#d7#)) OR
 					(reg_q480 AND symb_decoder(16#63#)) OR
 					(reg_q480 AND symb_decoder(16#29#)) OR
 					(reg_q480 AND symb_decoder(16#fe#)) OR
 					(reg_q480 AND symb_decoder(16#ef#)) OR
 					(reg_q480 AND symb_decoder(16#e1#)) OR
 					(reg_q480 AND symb_decoder(16#9f#)) OR
 					(reg_q480 AND symb_decoder(16#17#)) OR
 					(reg_q480 AND symb_decoder(16#1e#)) OR
 					(reg_q480 AND symb_decoder(16#ac#)) OR
 					(reg_q480 AND symb_decoder(16#a2#)) OR
 					(reg_q480 AND symb_decoder(16#2c#)) OR
 					(reg_q480 AND symb_decoder(16#25#)) OR
 					(reg_q480 AND symb_decoder(16#31#)) OR
 					(reg_q480 AND symb_decoder(16#97#)) OR
 					(reg_q480 AND symb_decoder(16#f3#)) OR
 					(reg_q480 AND symb_decoder(16#26#)) OR
 					(reg_q480 AND symb_decoder(16#2e#)) OR
 					(reg_q480 AND symb_decoder(16#91#)) OR
 					(reg_q480 AND symb_decoder(16#c6#)) OR
 					(reg_q480 AND symb_decoder(16#c7#)) OR
 					(reg_q480 AND symb_decoder(16#23#)) OR
 					(reg_q480 AND symb_decoder(16#1f#)) OR
 					(reg_q480 AND symb_decoder(16#e3#)) OR
 					(reg_q480 AND symb_decoder(16#bb#)) OR
 					(reg_q480 AND symb_decoder(16#75#)) OR
 					(reg_q480 AND symb_decoder(16#56#)) OR
 					(reg_q480 AND symb_decoder(16#02#)) OR
 					(reg_q480 AND symb_decoder(16#df#)) OR
 					(reg_q480 AND symb_decoder(16#54#)) OR
 					(reg_q480 AND symb_decoder(16#6d#)) OR
 					(reg_q480 AND symb_decoder(16#50#)) OR
 					(reg_q480 AND symb_decoder(16#1b#)) OR
 					(reg_q480 AND symb_decoder(16#a0#)) OR
 					(reg_q480 AND symb_decoder(16#bd#)) OR
 					(reg_q480 AND symb_decoder(16#62#)) OR
 					(reg_q480 AND symb_decoder(16#0e#)) OR
 					(reg_q480 AND symb_decoder(16#c9#)) OR
 					(reg_q480 AND symb_decoder(16#bf#)) OR
 					(reg_q480 AND symb_decoder(16#d9#)) OR
 					(reg_q480 AND symb_decoder(16#7d#)) OR
 					(reg_q480 AND symb_decoder(16#49#)) OR
 					(reg_q480 AND symb_decoder(16#c4#)) OR
 					(reg_q480 AND symb_decoder(16#37#)) OR
 					(reg_q480 AND symb_decoder(16#4a#)) OR
 					(reg_q480 AND symb_decoder(16#b8#)) OR
 					(reg_q480 AND symb_decoder(16#1d#)) OR
 					(reg_q480 AND symb_decoder(16#e4#)) OR
 					(reg_q480 AND symb_decoder(16#9e#)) OR
 					(reg_q480 AND symb_decoder(16#f2#)) OR
 					(reg_q480 AND symb_decoder(16#5d#)) OR
 					(reg_q480 AND symb_decoder(16#34#)) OR
 					(reg_q480 AND symb_decoder(16#d3#)) OR
 					(reg_q480 AND symb_decoder(16#52#)) OR
 					(reg_q480 AND symb_decoder(16#7c#)) OR
 					(reg_q480 AND symb_decoder(16#a4#)) OR
 					(reg_q480 AND symb_decoder(16#92#)) OR
 					(reg_q480 AND symb_decoder(16#68#)) OR
 					(reg_q480 AND symb_decoder(16#cd#)) OR
 					(reg_q480 AND symb_decoder(16#14#)) OR
 					(reg_q480 AND symb_decoder(16#0b#)) OR
 					(reg_q480 AND symb_decoder(16#f5#)) OR
 					(reg_q480 AND symb_decoder(16#13#)) OR
 					(reg_q480 AND symb_decoder(16#79#)) OR
 					(reg_q480 AND symb_decoder(16#03#)) OR
 					(reg_q480 AND symb_decoder(16#36#)) OR
 					(reg_q480 AND symb_decoder(16#4b#)) OR
 					(reg_q480 AND symb_decoder(16#15#)) OR
 					(reg_q480 AND symb_decoder(16#f7#)) OR
 					(reg_q480 AND symb_decoder(16#ba#)) OR
 					(reg_q480 AND symb_decoder(16#f6#)) OR
 					(reg_q480 AND symb_decoder(16#38#)) OR
 					(reg_q480 AND symb_decoder(16#f4#)) OR
 					(reg_q480 AND symb_decoder(16#3c#)) OR
 					(reg_q480 AND symb_decoder(16#89#)) OR
 					(reg_q480 AND symb_decoder(16#aa#)) OR
 					(reg_q480 AND symb_decoder(16#9c#)) OR
 					(reg_q480 AND symb_decoder(16#64#)) OR
 					(reg_q480 AND symb_decoder(16#b5#)) OR
 					(reg_q480 AND symb_decoder(16#fc#)) OR
 					(reg_q480 AND symb_decoder(16#9a#)) OR
 					(reg_q480 AND symb_decoder(16#8c#)) OR
 					(reg_q480 AND symb_decoder(16#53#)) OR
 					(reg_q480 AND symb_decoder(16#28#)) OR
 					(reg_q480 AND symb_decoder(16#b2#)) OR
 					(reg_q480 AND symb_decoder(16#4e#)) OR
 					(reg_q480 AND symb_decoder(16#30#)) OR
 					(reg_q480 AND symb_decoder(16#85#)) OR
 					(reg_q480 AND symb_decoder(16#5b#)) OR
 					(reg_q480 AND symb_decoder(16#05#)) OR
 					(reg_q480 AND symb_decoder(16#f0#)) OR
 					(reg_q480 AND symb_decoder(16#cf#)) OR
 					(reg_q480 AND symb_decoder(16#20#)) OR
 					(reg_q480 AND symb_decoder(16#09#)) OR
 					(reg_q480 AND symb_decoder(16#32#)) OR
 					(reg_q480 AND symb_decoder(16#90#)) OR
 					(reg_q480 AND symb_decoder(16#e5#)) OR
 					(reg_q480 AND symb_decoder(16#2a#)) OR
 					(reg_q480 AND symb_decoder(16#00#)) OR
 					(reg_q480 AND symb_decoder(16#93#)) OR
 					(reg_q480 AND symb_decoder(16#e0#)) OR
 					(reg_q480 AND symb_decoder(16#c1#)) OR
 					(reg_q480 AND symb_decoder(16#d6#)) OR
 					(reg_q480 AND symb_decoder(16#12#)) OR
 					(reg_q480 AND symb_decoder(16#af#)) OR
 					(reg_q480 AND symb_decoder(16#78#)) OR
 					(reg_q480 AND symb_decoder(16#83#)) OR
 					(reg_q480 AND symb_decoder(16#cb#)) OR
 					(reg_q480 AND symb_decoder(16#3b#)) OR
 					(reg_q480 AND symb_decoder(16#99#)) OR
 					(reg_q480 AND symb_decoder(16#ab#)) OR
 					(reg_q480 AND symb_decoder(16#88#)) OR
 					(reg_q480 AND symb_decoder(16#87#)) OR
 					(reg_q480 AND symb_decoder(16#43#)) OR
 					(reg_q480 AND symb_decoder(16#21#)) OR
 					(reg_q480 AND symb_decoder(16#4c#)) OR
 					(reg_q480 AND symb_decoder(16#be#)) OR
 					(reg_q480 AND symb_decoder(16#7e#)) OR
 					(reg_q480 AND symb_decoder(16#5f#)) OR
 					(reg_q480 AND symb_decoder(16#cc#)) OR
 					(reg_q480 AND symb_decoder(16#71#)) OR
 					(reg_q480 AND symb_decoder(16#8d#)) OR
 					(reg_q480 AND symb_decoder(16#ae#)) OR
 					(reg_q480 AND symb_decoder(16#b0#)) OR
 					(reg_q480 AND symb_decoder(16#1c#)) OR
 					(reg_q480 AND symb_decoder(16#a3#)) OR
 					(reg_q480 AND symb_decoder(16#a1#)) OR
 					(reg_q480 AND symb_decoder(16#3e#)) OR
 					(reg_q480 AND symb_decoder(16#c3#)) OR
 					(reg_q480 AND symb_decoder(16#7f#)) OR
 					(reg_q480 AND symb_decoder(16#47#)) OR
 					(reg_q480 AND symb_decoder(16#fb#)) OR
 					(reg_q480 AND symb_decoder(16#98#)) OR
 					(reg_q480 AND symb_decoder(16#d4#)) OR
 					(reg_q480 AND symb_decoder(16#74#)) OR
 					(reg_q480 AND symb_decoder(16#b6#)) OR
 					(reg_q480 AND symb_decoder(16#7a#)) OR
 					(reg_q480 AND symb_decoder(16#e9#)) OR
 					(reg_q480 AND symb_decoder(16#06#)) OR
 					(reg_q480 AND symb_decoder(16#b7#)) OR
 					(reg_q480 AND symb_decoder(16#fd#)) OR
 					(reg_q480 AND symb_decoder(16#3d#)) OR
 					(reg_q480 AND symb_decoder(16#0c#)) OR
 					(reg_q480 AND symb_decoder(16#11#)) OR
 					(reg_q480 AND symb_decoder(16#8e#)) OR
 					(reg_q480 AND symb_decoder(16#a8#)) OR
 					(reg_q480 AND symb_decoder(16#1a#)) OR
 					(reg_q480 AND symb_decoder(16#f9#)) OR
 					(reg_q480 AND symb_decoder(16#db#)) OR
 					(reg_q480 AND symb_decoder(16#57#)) OR
 					(reg_q480 AND symb_decoder(16#ca#)) OR
 					(reg_q480 AND symb_decoder(16#6c#)) OR
 					(reg_q480 AND symb_decoder(16#95#)) OR
 					(reg_q480 AND symb_decoder(16#b9#)) OR
 					(reg_q480 AND symb_decoder(16#5a#)) OR
 					(reg_q480 AND symb_decoder(16#19#)) OR
 					(reg_q480 AND symb_decoder(16#7b#)) OR
 					(reg_q480 AND symb_decoder(16#48#)) OR
 					(reg_q480 AND symb_decoder(16#a7#)) OR
 					(reg_q480 AND symb_decoder(16#41#)) OR
 					(reg_q480 AND symb_decoder(16#e7#)) OR
 					(reg_q480 AND symb_decoder(16#f1#)) OR
 					(reg_q480 AND symb_decoder(16#a9#)) OR
 					(reg_q480 AND symb_decoder(16#de#)) OR
 					(reg_q480 AND symb_decoder(16#c5#)) OR
 					(reg_q480 AND symb_decoder(16#22#)) OR
 					(reg_q480 AND symb_decoder(16#04#));
reg_q2526_in <= (reg_q2524 AND symb_decoder(16#20#));
reg_q377_in <= (reg_q375 AND symb_decoder(16#54#)) OR
 					(reg_q375 AND symb_decoder(16#74#));
reg_q185_in <= (reg_q185 AND symb_decoder(16#3c#)) OR
 					(reg_q185 AND symb_decoder(16#3b#)) OR
 					(reg_q185 AND symb_decoder(16#51#)) OR
 					(reg_q185 AND symb_decoder(16#c7#)) OR
 					(reg_q185 AND symb_decoder(16#7c#)) OR
 					(reg_q185 AND symb_decoder(16#7d#)) OR
 					(reg_q185 AND symb_decoder(16#ef#)) OR
 					(reg_q185 AND symb_decoder(16#34#)) OR
 					(reg_q185 AND symb_decoder(16#bd#)) OR
 					(reg_q185 AND symb_decoder(16#7f#)) OR
 					(reg_q185 AND symb_decoder(16#96#)) OR
 					(reg_q185 AND symb_decoder(16#fa#)) OR
 					(reg_q185 AND symb_decoder(16#9f#)) OR
 					(reg_q185 AND symb_decoder(16#fe#)) OR
 					(reg_q185 AND symb_decoder(16#f9#)) OR
 					(reg_q185 AND symb_decoder(16#5b#)) OR
 					(reg_q185 AND symb_decoder(16#69#)) OR
 					(reg_q185 AND symb_decoder(16#bf#)) OR
 					(reg_q185 AND symb_decoder(16#83#)) OR
 					(reg_q185 AND symb_decoder(16#22#)) OR
 					(reg_q185 AND symb_decoder(16#26#)) OR
 					(reg_q185 AND symb_decoder(16#c6#)) OR
 					(reg_q185 AND symb_decoder(16#b6#)) OR
 					(reg_q185 AND symb_decoder(16#8e#)) OR
 					(reg_q185 AND symb_decoder(16#f0#)) OR
 					(reg_q185 AND symb_decoder(16#fc#)) OR
 					(reg_q185 AND symb_decoder(16#86#)) OR
 					(reg_q185 AND symb_decoder(16#e0#)) OR
 					(reg_q185 AND symb_decoder(16#d4#)) OR
 					(reg_q185 AND symb_decoder(16#ee#)) OR
 					(reg_q185 AND symb_decoder(16#1a#)) OR
 					(reg_q185 AND symb_decoder(16#4e#)) OR
 					(reg_q185 AND symb_decoder(16#be#)) OR
 					(reg_q185 AND symb_decoder(16#e5#)) OR
 					(reg_q185 AND symb_decoder(16#6f#)) OR
 					(reg_q185 AND symb_decoder(16#91#)) OR
 					(reg_q185 AND symb_decoder(16#24#)) OR
 					(reg_q185 AND symb_decoder(16#1e#)) OR
 					(reg_q185 AND symb_decoder(16#a7#)) OR
 					(reg_q185 AND symb_decoder(16#f2#)) OR
 					(reg_q185 AND symb_decoder(16#ac#)) OR
 					(reg_q185 AND symb_decoder(16#02#)) OR
 					(reg_q185 AND symb_decoder(16#13#)) OR
 					(reg_q185 AND symb_decoder(16#28#)) OR
 					(reg_q185 AND symb_decoder(16#d6#)) OR
 					(reg_q185 AND symb_decoder(16#0c#)) OR
 					(reg_q185 AND symb_decoder(16#85#)) OR
 					(reg_q185 AND symb_decoder(16#67#)) OR
 					(reg_q185 AND symb_decoder(16#ce#)) OR
 					(reg_q185 AND symb_decoder(16#a6#)) OR
 					(reg_q185 AND symb_decoder(16#ae#)) OR
 					(reg_q185 AND symb_decoder(16#55#)) OR
 					(reg_q185 AND symb_decoder(16#de#)) OR
 					(reg_q185 AND symb_decoder(16#b5#)) OR
 					(reg_q185 AND symb_decoder(16#d9#)) OR
 					(reg_q185 AND symb_decoder(16#57#)) OR
 					(reg_q185 AND symb_decoder(16#89#)) OR
 					(reg_q185 AND symb_decoder(16#cc#)) OR
 					(reg_q185 AND symb_decoder(16#50#)) OR
 					(reg_q185 AND symb_decoder(16#a3#)) OR
 					(reg_q185 AND symb_decoder(16#99#)) OR
 					(reg_q185 AND symb_decoder(16#9d#)) OR
 					(reg_q185 AND symb_decoder(16#10#)) OR
 					(reg_q185 AND symb_decoder(16#e9#)) OR
 					(reg_q185 AND symb_decoder(16#cf#)) OR
 					(reg_q185 AND symb_decoder(16#e4#)) OR
 					(reg_q185 AND symb_decoder(16#d5#)) OR
 					(reg_q185 AND symb_decoder(16#95#)) OR
 					(reg_q185 AND symb_decoder(16#06#)) OR
 					(reg_q185 AND symb_decoder(16#70#)) OR
 					(reg_q185 AND symb_decoder(16#60#)) OR
 					(reg_q185 AND symb_decoder(16#53#)) OR
 					(reg_q185 AND symb_decoder(16#16#)) OR
 					(reg_q185 AND symb_decoder(16#0b#)) OR
 					(reg_q185 AND symb_decoder(16#2f#)) OR
 					(reg_q185 AND symb_decoder(16#b2#)) OR
 					(reg_q185 AND symb_decoder(16#e2#)) OR
 					(reg_q185 AND symb_decoder(16#1b#)) OR
 					(reg_q185 AND symb_decoder(16#df#)) OR
 					(reg_q185 AND symb_decoder(16#d1#)) OR
 					(reg_q185 AND symb_decoder(16#e3#)) OR
 					(reg_q185 AND symb_decoder(16#f8#)) OR
 					(reg_q185 AND symb_decoder(16#2a#)) OR
 					(reg_q185 AND symb_decoder(16#6d#)) OR
 					(reg_q185 AND symb_decoder(16#c9#)) OR
 					(reg_q185 AND symb_decoder(16#6a#)) OR
 					(reg_q185 AND symb_decoder(16#a8#)) OR
 					(reg_q185 AND symb_decoder(16#b9#)) OR
 					(reg_q185 AND symb_decoder(16#29#)) OR
 					(reg_q185 AND symb_decoder(16#b4#)) OR
 					(reg_q185 AND symb_decoder(16#f4#)) OR
 					(reg_q185 AND symb_decoder(16#54#)) OR
 					(reg_q185 AND symb_decoder(16#42#)) OR
 					(reg_q185 AND symb_decoder(16#d0#)) OR
 					(reg_q185 AND symb_decoder(16#33#)) OR
 					(reg_q185 AND symb_decoder(16#90#)) OR
 					(reg_q185 AND symb_decoder(16#58#)) OR
 					(reg_q185 AND symb_decoder(16#d2#)) OR
 					(reg_q185 AND symb_decoder(16#88#)) OR
 					(reg_q185 AND symb_decoder(16#d3#)) OR
 					(reg_q185 AND symb_decoder(16#97#)) OR
 					(reg_q185 AND symb_decoder(16#5e#)) OR
 					(reg_q185 AND symb_decoder(16#12#)) OR
 					(reg_q185 AND symb_decoder(16#47#)) OR
 					(reg_q185 AND symb_decoder(16#a0#)) OR
 					(reg_q185 AND symb_decoder(16#5d#)) OR
 					(reg_q185 AND symb_decoder(16#76#)) OR
 					(reg_q185 AND symb_decoder(16#f3#)) OR
 					(reg_q185 AND symb_decoder(16#ea#)) OR
 					(reg_q185 AND symb_decoder(16#73#)) OR
 					(reg_q185 AND symb_decoder(16#62#)) OR
 					(reg_q185 AND symb_decoder(16#15#)) OR
 					(reg_q185 AND symb_decoder(16#17#)) OR
 					(reg_q185 AND symb_decoder(16#44#)) OR
 					(reg_q185 AND symb_decoder(16#52#)) OR
 					(reg_q185 AND symb_decoder(16#3f#)) OR
 					(reg_q185 AND symb_decoder(16#7a#)) OR
 					(reg_q185 AND symb_decoder(16#8d#)) OR
 					(reg_q185 AND symb_decoder(16#3e#)) OR
 					(reg_q185 AND symb_decoder(16#87#)) OR
 					(reg_q185 AND symb_decoder(16#f6#)) OR
 					(reg_q185 AND symb_decoder(16#f5#)) OR
 					(reg_q185 AND symb_decoder(16#81#)) OR
 					(reg_q185 AND symb_decoder(16#5f#)) OR
 					(reg_q185 AND symb_decoder(16#0e#)) OR
 					(reg_q185 AND symb_decoder(16#65#)) OR
 					(reg_q185 AND symb_decoder(16#b8#)) OR
 					(reg_q185 AND symb_decoder(16#5c#)) OR
 					(reg_q185 AND symb_decoder(16#cd#)) OR
 					(reg_q185 AND symb_decoder(16#01#)) OR
 					(reg_q185 AND symb_decoder(16#cb#)) OR
 					(reg_q185 AND symb_decoder(16#8b#)) OR
 					(reg_q185 AND symb_decoder(16#e1#)) OR
 					(reg_q185 AND symb_decoder(16#04#)) OR
 					(reg_q185 AND symb_decoder(16#c0#)) OR
 					(reg_q185 AND symb_decoder(16#00#)) OR
 					(reg_q185 AND symb_decoder(16#75#)) OR
 					(reg_q185 AND symb_decoder(16#fb#)) OR
 					(reg_q185 AND symb_decoder(16#37#)) OR
 					(reg_q185 AND symb_decoder(16#94#)) OR
 					(reg_q185 AND symb_decoder(16#6c#)) OR
 					(reg_q185 AND symb_decoder(16#82#)) OR
 					(reg_q185 AND symb_decoder(16#ed#)) OR
 					(reg_q185 AND symb_decoder(16#6e#)) OR
 					(reg_q185 AND symb_decoder(16#eb#)) OR
 					(reg_q185 AND symb_decoder(16#2e#)) OR
 					(reg_q185 AND symb_decoder(16#74#)) OR
 					(reg_q185 AND symb_decoder(16#3d#)) OR
 					(reg_q185 AND symb_decoder(16#5a#)) OR
 					(reg_q185 AND symb_decoder(16#d7#)) OR
 					(reg_q185 AND symb_decoder(16#27#)) OR
 					(reg_q185 AND symb_decoder(16#63#)) OR
 					(reg_q185 AND symb_decoder(16#c8#)) OR
 					(reg_q185 AND symb_decoder(16#61#)) OR
 					(reg_q185 AND symb_decoder(16#66#)) OR
 					(reg_q185 AND symb_decoder(16#4b#)) OR
 					(reg_q185 AND symb_decoder(16#72#)) OR
 					(reg_q185 AND symb_decoder(16#ad#)) OR
 					(reg_q185 AND symb_decoder(16#31#)) OR
 					(reg_q185 AND symb_decoder(16#45#)) OR
 					(reg_q185 AND symb_decoder(16#3a#)) OR
 					(reg_q185 AND symb_decoder(16#41#)) OR
 					(reg_q185 AND symb_decoder(16#4f#)) OR
 					(reg_q185 AND symb_decoder(16#ba#)) OR
 					(reg_q185 AND symb_decoder(16#f7#)) OR
 					(reg_q185 AND symb_decoder(16#32#)) OR
 					(reg_q185 AND symb_decoder(16#bc#)) OR
 					(reg_q185 AND symb_decoder(16#1d#)) OR
 					(reg_q185 AND symb_decoder(16#2c#)) OR
 					(reg_q185 AND symb_decoder(16#db#)) OR
 					(reg_q185 AND symb_decoder(16#59#)) OR
 					(reg_q185 AND symb_decoder(16#23#)) OR
 					(reg_q185 AND symb_decoder(16#2d#)) OR
 					(reg_q185 AND symb_decoder(16#4c#)) OR
 					(reg_q185 AND symb_decoder(16#dc#)) OR
 					(reg_q185 AND symb_decoder(16#08#)) OR
 					(reg_q185 AND symb_decoder(16#48#)) OR
 					(reg_q185 AND symb_decoder(16#bb#)) OR
 					(reg_q185 AND symb_decoder(16#8f#)) OR
 					(reg_q185 AND symb_decoder(16#a9#)) OR
 					(reg_q185 AND symb_decoder(16#e6#)) OR
 					(reg_q185 AND symb_decoder(16#da#)) OR
 					(reg_q185 AND symb_decoder(16#4d#)) OR
 					(reg_q185 AND symb_decoder(16#71#)) OR
 					(reg_q185 AND symb_decoder(16#ff#)) OR
 					(reg_q185 AND symb_decoder(16#af#)) OR
 					(reg_q185 AND symb_decoder(16#a2#)) OR
 					(reg_q185 AND symb_decoder(16#9a#)) OR
 					(reg_q185 AND symb_decoder(16#c4#)) OR
 					(reg_q185 AND symb_decoder(16#05#)) OR
 					(reg_q185 AND symb_decoder(16#c5#)) OR
 					(reg_q185 AND symb_decoder(16#78#)) OR
 					(reg_q185 AND symb_decoder(16#39#)) OR
 					(reg_q185 AND symb_decoder(16#21#)) OR
 					(reg_q185 AND symb_decoder(16#46#)) OR
 					(reg_q185 AND symb_decoder(16#35#)) OR
 					(reg_q185 AND symb_decoder(16#6b#)) OR
 					(reg_q185 AND symb_decoder(16#36#)) OR
 					(reg_q185 AND symb_decoder(16#aa#)) OR
 					(reg_q185 AND symb_decoder(16#ec#)) OR
 					(reg_q185 AND symb_decoder(16#14#)) OR
 					(reg_q185 AND symb_decoder(16#b0#)) OR
 					(reg_q185 AND symb_decoder(16#a5#)) OR
 					(reg_q185 AND symb_decoder(16#18#)) OR
 					(reg_q185 AND symb_decoder(16#a1#)) OR
 					(reg_q185 AND symb_decoder(16#9b#)) OR
 					(reg_q185 AND symb_decoder(16#77#)) OR
 					(reg_q185 AND symb_decoder(16#30#)) OR
 					(reg_q185 AND symb_decoder(16#43#)) OR
 					(reg_q185 AND symb_decoder(16#4a#)) OR
 					(reg_q185 AND symb_decoder(16#b1#)) OR
 					(reg_q185 AND symb_decoder(16#11#)) OR
 					(reg_q185 AND symb_decoder(16#56#)) OR
 					(reg_q185 AND symb_decoder(16#1f#)) OR
 					(reg_q185 AND symb_decoder(16#03#)) OR
 					(reg_q185 AND symb_decoder(16#ca#)) OR
 					(reg_q185 AND symb_decoder(16#dd#)) OR
 					(reg_q185 AND symb_decoder(16#7b#)) OR
 					(reg_q185 AND symb_decoder(16#07#)) OR
 					(reg_q185 AND symb_decoder(16#38#)) OR
 					(reg_q185 AND symb_decoder(16#80#)) OR
 					(reg_q185 AND symb_decoder(16#40#)) OR
 					(reg_q185 AND symb_decoder(16#d8#)) OR
 					(reg_q185 AND symb_decoder(16#1c#)) OR
 					(reg_q185 AND symb_decoder(16#93#)) OR
 					(reg_q185 AND symb_decoder(16#68#)) OR
 					(reg_q185 AND symb_decoder(16#9c#)) OR
 					(reg_q185 AND symb_decoder(16#25#)) OR
 					(reg_q185 AND symb_decoder(16#8c#)) OR
 					(reg_q185 AND symb_decoder(16#b7#)) OR
 					(reg_q185 AND symb_decoder(16#92#)) OR
 					(reg_q185 AND symb_decoder(16#98#)) OR
 					(reg_q185 AND symb_decoder(16#2b#)) OR
 					(reg_q185 AND symb_decoder(16#09#)) OR
 					(reg_q185 AND symb_decoder(16#7e#)) OR
 					(reg_q185 AND symb_decoder(16#8a#)) OR
 					(reg_q185 AND symb_decoder(16#79#)) OR
 					(reg_q185 AND symb_decoder(16#e8#)) OR
 					(reg_q185 AND symb_decoder(16#49#)) OR
 					(reg_q185 AND symb_decoder(16#19#)) OR
 					(reg_q185 AND symb_decoder(16#0f#)) OR
 					(reg_q185 AND symb_decoder(16#c3#)) OR
 					(reg_q185 AND symb_decoder(16#64#)) OR
 					(reg_q185 AND symb_decoder(16#20#)) OR
 					(reg_q185 AND symb_decoder(16#f1#)) OR
 					(reg_q185 AND symb_decoder(16#9e#)) OR
 					(reg_q185 AND symb_decoder(16#ab#)) OR
 					(reg_q185 AND symb_decoder(16#c2#)) OR
 					(reg_q185 AND symb_decoder(16#fd#)) OR
 					(reg_q185 AND symb_decoder(16#84#)) OR
 					(reg_q185 AND symb_decoder(16#a4#)) OR
 					(reg_q185 AND symb_decoder(16#c1#)) OR
 					(reg_q185 AND symb_decoder(16#e7#)) OR
 					(reg_q185 AND symb_decoder(16#b3#)) OR
 					(reg_q173 AND symb_decoder(16#13#)) OR
 					(reg_q173 AND symb_decoder(16#87#)) OR
 					(reg_q173 AND symb_decoder(16#14#)) OR
 					(reg_q173 AND symb_decoder(16#d2#)) OR
 					(reg_q173 AND symb_decoder(16#63#)) OR
 					(reg_q173 AND symb_decoder(16#59#)) OR
 					(reg_q173 AND symb_decoder(16#f9#)) OR
 					(reg_q173 AND symb_decoder(16#28#)) OR
 					(reg_q173 AND symb_decoder(16#d1#)) OR
 					(reg_q173 AND symb_decoder(16#4b#)) OR
 					(reg_q173 AND symb_decoder(16#52#)) OR
 					(reg_q173 AND symb_decoder(16#de#)) OR
 					(reg_q173 AND symb_decoder(16#43#)) OR
 					(reg_q173 AND symb_decoder(16#44#)) OR
 					(reg_q173 AND symb_decoder(16#c1#)) OR
 					(reg_q173 AND symb_decoder(16#a9#)) OR
 					(reg_q173 AND symb_decoder(16#f4#)) OR
 					(reg_q173 AND symb_decoder(16#af#)) OR
 					(reg_q173 AND symb_decoder(16#d3#)) OR
 					(reg_q173 AND symb_decoder(16#ce#)) OR
 					(reg_q173 AND symb_decoder(16#f5#)) OR
 					(reg_q173 AND symb_decoder(16#a6#)) OR
 					(reg_q173 AND symb_decoder(16#5e#)) OR
 					(reg_q173 AND symb_decoder(16#e7#)) OR
 					(reg_q173 AND symb_decoder(16#aa#)) OR
 					(reg_q173 AND symb_decoder(16#6a#)) OR
 					(reg_q173 AND symb_decoder(16#b0#)) OR
 					(reg_q173 AND symb_decoder(16#8f#)) OR
 					(reg_q173 AND symb_decoder(16#9d#)) OR
 					(reg_q173 AND symb_decoder(16#2e#)) OR
 					(reg_q173 AND symb_decoder(16#81#)) OR
 					(reg_q173 AND symb_decoder(16#48#)) OR
 					(reg_q173 AND symb_decoder(16#3c#)) OR
 					(reg_q173 AND symb_decoder(16#41#)) OR
 					(reg_q173 AND symb_decoder(16#ee#)) OR
 					(reg_q173 AND symb_decoder(16#2c#)) OR
 					(reg_q173 AND symb_decoder(16#a8#)) OR
 					(reg_q173 AND symb_decoder(16#45#)) OR
 					(reg_q173 AND symb_decoder(16#26#)) OR
 					(reg_q173 AND symb_decoder(16#ff#)) OR
 					(reg_q173 AND symb_decoder(16#9b#)) OR
 					(reg_q173 AND symb_decoder(16#d6#)) OR
 					(reg_q173 AND symb_decoder(16#01#)) OR
 					(reg_q173 AND symb_decoder(16#ca#)) OR
 					(reg_q173 AND symb_decoder(16#39#)) OR
 					(reg_q173 AND symb_decoder(16#0b#)) OR
 					(reg_q173 AND symb_decoder(16#10#)) OR
 					(reg_q173 AND symb_decoder(16#c0#)) OR
 					(reg_q173 AND symb_decoder(16#7f#)) OR
 					(reg_q173 AND symb_decoder(16#e6#)) OR
 					(reg_q173 AND symb_decoder(16#eb#)) OR
 					(reg_q173 AND symb_decoder(16#36#)) OR
 					(reg_q173 AND symb_decoder(16#33#)) OR
 					(reg_q173 AND symb_decoder(16#61#)) OR
 					(reg_q173 AND symb_decoder(16#73#)) OR
 					(reg_q173 AND symb_decoder(16#82#)) OR
 					(reg_q173 AND symb_decoder(16#cb#)) OR
 					(reg_q173 AND symb_decoder(16#83#)) OR
 					(reg_q173 AND symb_decoder(16#86#)) OR
 					(reg_q173 AND symb_decoder(16#12#)) OR
 					(reg_q173 AND symb_decoder(16#b1#)) OR
 					(reg_q173 AND symb_decoder(16#be#)) OR
 					(reg_q173 AND symb_decoder(16#bd#)) OR
 					(reg_q173 AND symb_decoder(16#db#)) OR
 					(reg_q173 AND symb_decoder(16#32#)) OR
 					(reg_q173 AND symb_decoder(16#30#)) OR
 					(reg_q173 AND symb_decoder(16#c2#)) OR
 					(reg_q173 AND symb_decoder(16#8d#)) OR
 					(reg_q173 AND symb_decoder(16#e3#)) OR
 					(reg_q173 AND symb_decoder(16#d0#)) OR
 					(reg_q173 AND symb_decoder(16#ac#)) OR
 					(reg_q173 AND symb_decoder(16#9c#)) OR
 					(reg_q173 AND symb_decoder(16#04#)) OR
 					(reg_q173 AND symb_decoder(16#d8#)) OR
 					(reg_q173 AND symb_decoder(16#3e#)) OR
 					(reg_q173 AND symb_decoder(16#88#)) OR
 					(reg_q173 AND symb_decoder(16#0c#)) OR
 					(reg_q173 AND symb_decoder(16#3b#)) OR
 					(reg_q173 AND symb_decoder(16#6e#)) OR
 					(reg_q173 AND symb_decoder(16#11#)) OR
 					(reg_q173 AND symb_decoder(16#a0#)) OR
 					(reg_q173 AND symb_decoder(16#35#)) OR
 					(reg_q173 AND symb_decoder(16#7d#)) OR
 					(reg_q173 AND symb_decoder(16#75#)) OR
 					(reg_q173 AND symb_decoder(16#f3#)) OR
 					(reg_q173 AND symb_decoder(16#90#)) OR
 					(reg_q173 AND symb_decoder(16#7a#)) OR
 					(reg_q173 AND symb_decoder(16#b2#)) OR
 					(reg_q173 AND symb_decoder(16#3d#)) OR
 					(reg_q173 AND symb_decoder(16#ba#)) OR
 					(reg_q173 AND symb_decoder(16#93#)) OR
 					(reg_q173 AND symb_decoder(16#62#)) OR
 					(reg_q173 AND symb_decoder(16#8c#)) OR
 					(reg_q173 AND symb_decoder(16#72#)) OR
 					(reg_q173 AND symb_decoder(16#c6#)) OR
 					(reg_q173 AND symb_decoder(16#c4#)) OR
 					(reg_q173 AND symb_decoder(16#1e#)) OR
 					(reg_q173 AND symb_decoder(16#27#)) OR
 					(reg_q173 AND symb_decoder(16#00#)) OR
 					(reg_q173 AND symb_decoder(16#84#)) OR
 					(reg_q173 AND symb_decoder(16#23#)) OR
 					(reg_q173 AND symb_decoder(16#8b#)) OR
 					(reg_q173 AND symb_decoder(16#4f#)) OR
 					(reg_q173 AND symb_decoder(16#79#)) OR
 					(reg_q173 AND symb_decoder(16#4a#)) OR
 					(reg_q173 AND symb_decoder(16#31#)) OR
 					(reg_q173 AND symb_decoder(16#b4#)) OR
 					(reg_q173 AND symb_decoder(16#c7#)) OR
 					(reg_q173 AND symb_decoder(16#1c#)) OR
 					(reg_q173 AND symb_decoder(16#dc#)) OR
 					(reg_q173 AND symb_decoder(16#20#)) OR
 					(reg_q173 AND symb_decoder(16#47#)) OR
 					(reg_q173 AND symb_decoder(16#24#)) OR
 					(reg_q173 AND symb_decoder(16#67#)) OR
 					(reg_q173 AND symb_decoder(16#55#)) OR
 					(reg_q173 AND symb_decoder(16#60#)) OR
 					(reg_q173 AND symb_decoder(16#e2#)) OR
 					(reg_q173 AND symb_decoder(16#37#)) OR
 					(reg_q173 AND symb_decoder(16#74#)) OR
 					(reg_q173 AND symb_decoder(16#0f#)) OR
 					(reg_q173 AND symb_decoder(16#5b#)) OR
 					(reg_q173 AND symb_decoder(16#5d#)) OR
 					(reg_q173 AND symb_decoder(16#09#)) OR
 					(reg_q173 AND symb_decoder(16#e5#)) OR
 					(reg_q173 AND symb_decoder(16#4e#)) OR
 					(reg_q173 AND symb_decoder(16#99#)) OR
 					(reg_q173 AND symb_decoder(16#21#)) OR
 					(reg_q173 AND symb_decoder(16#9f#)) OR
 					(reg_q173 AND symb_decoder(16#6b#)) OR
 					(reg_q173 AND symb_decoder(16#15#)) OR
 					(reg_q173 AND symb_decoder(16#ef#)) OR
 					(reg_q173 AND symb_decoder(16#fe#)) OR
 					(reg_q173 AND symb_decoder(16#1f#)) OR
 					(reg_q173 AND symb_decoder(16#f2#)) OR
 					(reg_q173 AND symb_decoder(16#d9#)) OR
 					(reg_q173 AND symb_decoder(16#53#)) OR
 					(reg_q173 AND symb_decoder(16#a3#)) OR
 					(reg_q173 AND symb_decoder(16#64#)) OR
 					(reg_q173 AND symb_decoder(16#e4#)) OR
 					(reg_q173 AND symb_decoder(16#7c#)) OR
 					(reg_q173 AND symb_decoder(16#5f#)) OR
 					(reg_q173 AND symb_decoder(16#6f#)) OR
 					(reg_q173 AND symb_decoder(16#ab#)) OR
 					(reg_q173 AND symb_decoder(16#78#)) OR
 					(reg_q173 AND symb_decoder(16#2a#)) OR
 					(reg_q173 AND symb_decoder(16#51#)) OR
 					(reg_q173 AND symb_decoder(16#c3#)) OR
 					(reg_q173 AND symb_decoder(16#6c#)) OR
 					(reg_q173 AND symb_decoder(16#8e#)) OR
 					(reg_q173 AND symb_decoder(16#9e#)) OR
 					(reg_q173 AND symb_decoder(16#3a#)) OR
 					(reg_q173 AND symb_decoder(16#2d#)) OR
 					(reg_q173 AND symb_decoder(16#06#)) OR
 					(reg_q173 AND symb_decoder(16#a7#)) OR
 					(reg_q173 AND symb_decoder(16#08#)) OR
 					(reg_q173 AND symb_decoder(16#42#)) OR
 					(reg_q173 AND symb_decoder(16#dd#)) OR
 					(reg_q173 AND symb_decoder(16#71#)) OR
 					(reg_q173 AND symb_decoder(16#fb#)) OR
 					(reg_q173 AND symb_decoder(16#e8#)) OR
 					(reg_q173 AND symb_decoder(16#85#)) OR
 					(reg_q173 AND symb_decoder(16#38#)) OR
 					(reg_q173 AND symb_decoder(16#f7#)) OR
 					(reg_q173 AND symb_decoder(16#b7#)) OR
 					(reg_q173 AND symb_decoder(16#2b#)) OR
 					(reg_q173 AND symb_decoder(16#7e#)) OR
 					(reg_q173 AND symb_decoder(16#66#)) OR
 					(reg_q173 AND symb_decoder(16#18#)) OR
 					(reg_q173 AND symb_decoder(16#89#)) OR
 					(reg_q173 AND symb_decoder(16#cd#)) OR
 					(reg_q173 AND symb_decoder(16#69#)) OR
 					(reg_q173 AND symb_decoder(16#17#)) OR
 					(reg_q173 AND symb_decoder(16#03#)) OR
 					(reg_q173 AND symb_decoder(16#6d#)) OR
 					(reg_q173 AND symb_decoder(16#98#)) OR
 					(reg_q173 AND symb_decoder(16#16#)) OR
 					(reg_q173 AND symb_decoder(16#58#)) OR
 					(reg_q173 AND symb_decoder(16#02#)) OR
 					(reg_q173 AND symb_decoder(16#d4#)) OR
 					(reg_q173 AND symb_decoder(16#da#)) OR
 					(reg_q173 AND symb_decoder(16#ea#)) OR
 					(reg_q173 AND symb_decoder(16#56#)) OR
 					(reg_q173 AND symb_decoder(16#fd#)) OR
 					(reg_q173 AND symb_decoder(16#5a#)) OR
 					(reg_q173 AND symb_decoder(16#8a#)) OR
 					(reg_q173 AND symb_decoder(16#a2#)) OR
 					(reg_q173 AND symb_decoder(16#65#)) OR
 					(reg_q173 AND symb_decoder(16#05#)) OR
 					(reg_q173 AND symb_decoder(16#1d#)) OR
 					(reg_q173 AND symb_decoder(16#b5#)) OR
 					(reg_q173 AND symb_decoder(16#70#)) OR
 					(reg_q173 AND symb_decoder(16#e0#)) OR
 					(reg_q173 AND symb_decoder(16#cc#)) OR
 					(reg_q173 AND symb_decoder(16#94#)) OR
 					(reg_q173 AND symb_decoder(16#9a#)) OR
 					(reg_q173 AND symb_decoder(16#b3#)) OR
 					(reg_q173 AND symb_decoder(16#fa#)) OR
 					(reg_q173 AND symb_decoder(16#97#)) OR
 					(reg_q173 AND symb_decoder(16#1a#)) OR
 					(reg_q173 AND symb_decoder(16#b8#)) OR
 					(reg_q173 AND symb_decoder(16#77#)) OR
 					(reg_q173 AND symb_decoder(16#d7#)) OR
 					(reg_q173 AND symb_decoder(16#a4#)) OR
 					(reg_q173 AND symb_decoder(16#c5#)) OR
 					(reg_q173 AND symb_decoder(16#7b#)) OR
 					(reg_q173 AND symb_decoder(16#bc#)) OR
 					(reg_q173 AND symb_decoder(16#f1#)) OR
 					(reg_q173 AND symb_decoder(16#d5#)) OR
 					(reg_q173 AND symb_decoder(16#e9#)) OR
 					(reg_q173 AND symb_decoder(16#e1#)) OR
 					(reg_q173 AND symb_decoder(16#bb#)) OR
 					(reg_q173 AND symb_decoder(16#80#)) OR
 					(reg_q173 AND symb_decoder(16#1b#)) OR
 					(reg_q173 AND symb_decoder(16#50#)) OR
 					(reg_q173 AND symb_decoder(16#a1#)) OR
 					(reg_q173 AND symb_decoder(16#07#)) OR
 					(reg_q173 AND symb_decoder(16#91#)) OR
 					(reg_q173 AND symb_decoder(16#f0#)) OR
 					(reg_q173 AND symb_decoder(16#96#)) OR
 					(reg_q173 AND symb_decoder(16#ad#)) OR
 					(reg_q173 AND symb_decoder(16#b9#)) OR
 					(reg_q173 AND symb_decoder(16#46#)) OR
 					(reg_q173 AND symb_decoder(16#bf#)) OR
 					(reg_q173 AND symb_decoder(16#49#)) OR
 					(reg_q173 AND symb_decoder(16#25#)) OR
 					(reg_q173 AND symb_decoder(16#29#)) OR
 					(reg_q173 AND symb_decoder(16#22#)) OR
 					(reg_q173 AND symb_decoder(16#0e#)) OR
 					(reg_q173 AND symb_decoder(16#54#)) OR
 					(reg_q173 AND symb_decoder(16#34#)) OR
 					(reg_q173 AND symb_decoder(16#57#)) OR
 					(reg_q173 AND symb_decoder(16#df#)) OR
 					(reg_q173 AND symb_decoder(16#5c#)) OR
 					(reg_q173 AND symb_decoder(16#c9#)) OR
 					(reg_q173 AND symb_decoder(16#f8#)) OR
 					(reg_q173 AND symb_decoder(16#4d#)) OR
 					(reg_q173 AND symb_decoder(16#fc#)) OR
 					(reg_q173 AND symb_decoder(16#ae#)) OR
 					(reg_q173 AND symb_decoder(16#a5#)) OR
 					(reg_q173 AND symb_decoder(16#3f#)) OR
 					(reg_q173 AND symb_decoder(16#2f#)) OR
 					(reg_q173 AND symb_decoder(16#f6#)) OR
 					(reg_q173 AND symb_decoder(16#b6#)) OR
 					(reg_q173 AND symb_decoder(16#ec#)) OR
 					(reg_q173 AND symb_decoder(16#68#)) OR
 					(reg_q173 AND symb_decoder(16#4c#)) OR
 					(reg_q173 AND symb_decoder(16#92#)) OR
 					(reg_q173 AND symb_decoder(16#c8#)) OR
 					(reg_q173 AND symb_decoder(16#76#)) OR
 					(reg_q173 AND symb_decoder(16#ed#)) OR
 					(reg_q173 AND symb_decoder(16#19#)) OR
 					(reg_q173 AND symb_decoder(16#40#)) OR
 					(reg_q173 AND symb_decoder(16#95#)) OR
 					(reg_q173 AND symb_decoder(16#cf#));
reg_q522_in <= (reg_q520 AND symb_decoder(16#6e#)) OR
 					(reg_q520 AND symb_decoder(16#4e#));
reg_q1719_in <= (reg_q1719 AND symb_decoder(16#32#)) OR
 					(reg_q1719 AND symb_decoder(16#37#)) OR
 					(reg_q1719 AND symb_decoder(16#39#)) OR
 					(reg_q1719 AND symb_decoder(16#35#)) OR
 					(reg_q1719 AND symb_decoder(16#38#)) OR
 					(reg_q1719 AND symb_decoder(16#31#)) OR
 					(reg_q1719 AND symb_decoder(16#36#)) OR
 					(reg_q1719 AND symb_decoder(16#34#)) OR
 					(reg_q1719 AND symb_decoder(16#33#)) OR
 					(reg_q1719 AND symb_decoder(16#30#)) OR
 					(reg_q1717 AND symb_decoder(16#34#)) OR
 					(reg_q1717 AND symb_decoder(16#33#)) OR
 					(reg_q1717 AND symb_decoder(16#30#)) OR
 					(reg_q1717 AND symb_decoder(16#36#)) OR
 					(reg_q1717 AND symb_decoder(16#31#)) OR
 					(reg_q1717 AND symb_decoder(16#35#)) OR
 					(reg_q1717 AND symb_decoder(16#39#)) OR
 					(reg_q1717 AND symb_decoder(16#38#)) OR
 					(reg_q1717 AND symb_decoder(16#32#)) OR
 					(reg_q1717 AND symb_decoder(16#37#));
reg_q2736_in <= (reg_q2734 AND symb_decoder(16#0c#)) OR
 					(reg_q2734 AND symb_decoder(16#0a#)) OR
 					(reg_q2734 AND symb_decoder(16#09#)) OR
 					(reg_q2734 AND symb_decoder(16#0d#)) OR
 					(reg_q2734 AND symb_decoder(16#20#));
reg_q2738_in <= (reg_q2736 AND symb_decoder(16#73#)) OR
 					(reg_q2736 AND symb_decoder(16#53#));
reg_q876_in <= (reg_q874 AND symb_decoder(16#3a#));
reg_q942_in <= (reg_q876 AND symb_decoder(16#d9#)) OR
 					(reg_q876 AND symb_decoder(16#77#)) OR
 					(reg_q876 AND symb_decoder(16#8d#)) OR
 					(reg_q876 AND symb_decoder(16#f7#)) OR
 					(reg_q876 AND symb_decoder(16#a4#)) OR
 					(reg_q876 AND symb_decoder(16#35#)) OR
 					(reg_q876 AND symb_decoder(16#cb#)) OR
 					(reg_q876 AND symb_decoder(16#58#)) OR
 					(reg_q876 AND symb_decoder(16#c7#)) OR
 					(reg_q876 AND symb_decoder(16#9c#)) OR
 					(reg_q876 AND symb_decoder(16#27#)) OR
 					(reg_q876 AND symb_decoder(16#d3#)) OR
 					(reg_q876 AND symb_decoder(16#37#)) OR
 					(reg_q876 AND symb_decoder(16#a0#)) OR
 					(reg_q876 AND symb_decoder(16#7a#)) OR
 					(reg_q876 AND symb_decoder(16#e1#)) OR
 					(reg_q876 AND symb_decoder(16#c9#)) OR
 					(reg_q876 AND symb_decoder(16#75#)) OR
 					(reg_q876 AND symb_decoder(16#17#)) OR
 					(reg_q876 AND symb_decoder(16#2a#)) OR
 					(reg_q876 AND symb_decoder(16#12#)) OR
 					(reg_q876 AND symb_decoder(16#41#)) OR
 					(reg_q876 AND symb_decoder(16#c1#)) OR
 					(reg_q876 AND symb_decoder(16#a5#)) OR
 					(reg_q876 AND symb_decoder(16#5a#)) OR
 					(reg_q876 AND symb_decoder(16#1e#)) OR
 					(reg_q876 AND symb_decoder(16#c3#)) OR
 					(reg_q876 AND symb_decoder(16#95#)) OR
 					(reg_q876 AND symb_decoder(16#84#)) OR
 					(reg_q876 AND symb_decoder(16#d2#)) OR
 					(reg_q876 AND symb_decoder(16#26#)) OR
 					(reg_q876 AND symb_decoder(16#01#)) OR
 					(reg_q876 AND symb_decoder(16#4a#)) OR
 					(reg_q876 AND symb_decoder(16#21#)) OR
 					(reg_q876 AND symb_decoder(16#9a#)) OR
 					(reg_q876 AND symb_decoder(16#16#)) OR
 					(reg_q876 AND symb_decoder(16#00#)) OR
 					(reg_q876 AND symb_decoder(16#8f#)) OR
 					(reg_q876 AND symb_decoder(16#76#)) OR
 					(reg_q876 AND symb_decoder(16#29#)) OR
 					(reg_q876 AND symb_decoder(16#71#)) OR
 					(reg_q876 AND symb_decoder(16#da#)) OR
 					(reg_q876 AND symb_decoder(16#f9#)) OR
 					(reg_q876 AND symb_decoder(16#92#)) OR
 					(reg_q876 AND symb_decoder(16#8b#)) OR
 					(reg_q876 AND symb_decoder(16#bb#)) OR
 					(reg_q876 AND symb_decoder(16#d7#)) OR
 					(reg_q876 AND symb_decoder(16#c4#)) OR
 					(reg_q876 AND symb_decoder(16#b5#)) OR
 					(reg_q876 AND symb_decoder(16#e4#)) OR
 					(reg_q876 AND symb_decoder(16#1a#)) OR
 					(reg_q876 AND symb_decoder(16#66#)) OR
 					(reg_q876 AND symb_decoder(16#b3#)) OR
 					(reg_q876 AND symb_decoder(16#6e#)) OR
 					(reg_q876 AND symb_decoder(16#90#)) OR
 					(reg_q876 AND symb_decoder(16#96#)) OR
 					(reg_q876 AND symb_decoder(16#94#)) OR
 					(reg_q876 AND symb_decoder(16#d8#)) OR
 					(reg_q876 AND symb_decoder(16#46#)) OR
 					(reg_q876 AND symb_decoder(16#c2#)) OR
 					(reg_q876 AND symb_decoder(16#9b#)) OR
 					(reg_q876 AND symb_decoder(16#1b#)) OR
 					(reg_q876 AND symb_decoder(16#04#)) OR
 					(reg_q876 AND symb_decoder(16#30#)) OR
 					(reg_q876 AND symb_decoder(16#19#)) OR
 					(reg_q876 AND symb_decoder(16#0e#)) OR
 					(reg_q876 AND symb_decoder(16#73#)) OR
 					(reg_q876 AND symb_decoder(16#c8#)) OR
 					(reg_q876 AND symb_decoder(16#b6#)) OR
 					(reg_q876 AND symb_decoder(16#bf#)) OR
 					(reg_q876 AND symb_decoder(16#1d#)) OR
 					(reg_q876 AND symb_decoder(16#10#)) OR
 					(reg_q876 AND symb_decoder(16#b9#)) OR
 					(reg_q876 AND symb_decoder(16#d4#)) OR
 					(reg_q876 AND symb_decoder(16#eb#)) OR
 					(reg_q876 AND symb_decoder(16#ff#)) OR
 					(reg_q876 AND symb_decoder(16#50#)) OR
 					(reg_q876 AND symb_decoder(16#e6#)) OR
 					(reg_q876 AND symb_decoder(16#b8#)) OR
 					(reg_q876 AND symb_decoder(16#68#)) OR
 					(reg_q876 AND symb_decoder(16#be#)) OR
 					(reg_q876 AND symb_decoder(16#32#)) OR
 					(reg_q876 AND symb_decoder(16#d6#)) OR
 					(reg_q876 AND symb_decoder(16#2b#)) OR
 					(reg_q876 AND symb_decoder(16#a3#)) OR
 					(reg_q876 AND symb_decoder(16#91#)) OR
 					(reg_q876 AND symb_decoder(16#ba#)) OR
 					(reg_q876 AND symb_decoder(16#23#)) OR
 					(reg_q876 AND symb_decoder(16#85#)) OR
 					(reg_q876 AND symb_decoder(16#63#)) OR
 					(reg_q876 AND symb_decoder(16#5f#)) OR
 					(reg_q876 AND symb_decoder(16#25#)) OR
 					(reg_q876 AND symb_decoder(16#3d#)) OR
 					(reg_q876 AND symb_decoder(16#03#)) OR
 					(reg_q876 AND symb_decoder(16#20#)) OR
 					(reg_q876 AND symb_decoder(16#81#)) OR
 					(reg_q876 AND symb_decoder(16#02#)) OR
 					(reg_q876 AND symb_decoder(16#dd#)) OR
 					(reg_q876 AND symb_decoder(16#4f#)) OR
 					(reg_q876 AND symb_decoder(16#4d#)) OR
 					(reg_q876 AND symb_decoder(16#c6#)) OR
 					(reg_q876 AND symb_decoder(16#9d#)) OR
 					(reg_q876 AND symb_decoder(16#b7#)) OR
 					(reg_q876 AND symb_decoder(16#d1#)) OR
 					(reg_q876 AND symb_decoder(16#fe#)) OR
 					(reg_q876 AND symb_decoder(16#7e#)) OR
 					(reg_q876 AND symb_decoder(16#b2#)) OR
 					(reg_q876 AND symb_decoder(16#87#)) OR
 					(reg_q876 AND symb_decoder(16#3f#)) OR
 					(reg_q876 AND symb_decoder(16#05#)) OR
 					(reg_q876 AND symb_decoder(16#e8#)) OR
 					(reg_q876 AND symb_decoder(16#bc#)) OR
 					(reg_q876 AND symb_decoder(16#ec#)) OR
 					(reg_q876 AND symb_decoder(16#13#)) OR
 					(reg_q876 AND symb_decoder(16#51#)) OR
 					(reg_q876 AND symb_decoder(16#2c#)) OR
 					(reg_q876 AND symb_decoder(16#39#)) OR
 					(reg_q876 AND symb_decoder(16#08#)) OR
 					(reg_q876 AND symb_decoder(16#86#)) OR
 					(reg_q876 AND symb_decoder(16#a6#)) OR
 					(reg_q876 AND symb_decoder(16#74#)) OR
 					(reg_q876 AND symb_decoder(16#ea#)) OR
 					(reg_q876 AND symb_decoder(16#83#)) OR
 					(reg_q876 AND symb_decoder(16#97#)) OR
 					(reg_q876 AND symb_decoder(16#40#)) OR
 					(reg_q876 AND symb_decoder(16#ed#)) OR
 					(reg_q876 AND symb_decoder(16#d5#)) OR
 					(reg_q876 AND symb_decoder(16#5e#)) OR
 					(reg_q876 AND symb_decoder(16#6d#)) OR
 					(reg_q876 AND symb_decoder(16#49#)) OR
 					(reg_q876 AND symb_decoder(16#4e#)) OR
 					(reg_q876 AND symb_decoder(16#72#)) OR
 					(reg_q876 AND symb_decoder(16#22#)) OR
 					(reg_q876 AND symb_decoder(16#14#)) OR
 					(reg_q876 AND symb_decoder(16#34#)) OR
 					(reg_q876 AND symb_decoder(16#a9#)) OR
 					(reg_q876 AND symb_decoder(16#93#)) OR
 					(reg_q876 AND symb_decoder(16#f1#)) OR
 					(reg_q876 AND symb_decoder(16#f4#)) OR
 					(reg_q876 AND symb_decoder(16#3c#)) OR
 					(reg_q876 AND symb_decoder(16#e2#)) OR
 					(reg_q876 AND symb_decoder(16#38#)) OR
 					(reg_q876 AND symb_decoder(16#98#)) OR
 					(reg_q876 AND symb_decoder(16#e5#)) OR
 					(reg_q876 AND symb_decoder(16#82#)) OR
 					(reg_q876 AND symb_decoder(16#78#)) OR
 					(reg_q876 AND symb_decoder(16#b0#)) OR
 					(reg_q876 AND symb_decoder(16#cc#)) OR
 					(reg_q876 AND symb_decoder(16#bd#)) OR
 					(reg_q876 AND symb_decoder(16#0c#)) OR
 					(reg_q876 AND symb_decoder(16#79#)) OR
 					(reg_q876 AND symb_decoder(16#fb#)) OR
 					(reg_q876 AND symb_decoder(16#80#)) OR
 					(reg_q876 AND symb_decoder(16#6b#)) OR
 					(reg_q876 AND symb_decoder(16#6f#)) OR
 					(reg_q876 AND symb_decoder(16#ee#)) OR
 					(reg_q876 AND symb_decoder(16#4b#)) OR
 					(reg_q876 AND symb_decoder(16#ad#)) OR
 					(reg_q876 AND symb_decoder(16#f5#)) OR
 					(reg_q876 AND symb_decoder(16#15#)) OR
 					(reg_q876 AND symb_decoder(16#ef#)) OR
 					(reg_q876 AND symb_decoder(16#0b#)) OR
 					(reg_q876 AND symb_decoder(16#69#)) OR
 					(reg_q876 AND symb_decoder(16#cf#)) OR
 					(reg_q876 AND symb_decoder(16#fd#)) OR
 					(reg_q876 AND symb_decoder(16#ae#)) OR
 					(reg_q876 AND symb_decoder(16#56#)) OR
 					(reg_q876 AND symb_decoder(16#f2#)) OR
 					(reg_q876 AND symb_decoder(16#88#)) OR
 					(reg_q876 AND symb_decoder(16#d0#)) OR
 					(reg_q876 AND symb_decoder(16#36#)) OR
 					(reg_q876 AND symb_decoder(16#3e#)) OR
 					(reg_q876 AND symb_decoder(16#6c#)) OR
 					(reg_q876 AND symb_decoder(16#11#)) OR
 					(reg_q876 AND symb_decoder(16#31#)) OR
 					(reg_q876 AND symb_decoder(16#f6#)) OR
 					(reg_q876 AND symb_decoder(16#61#)) OR
 					(reg_q876 AND symb_decoder(16#89#)) OR
 					(reg_q876 AND symb_decoder(16#e3#)) OR
 					(reg_q876 AND symb_decoder(16#4c#)) OR
 					(reg_q876 AND symb_decoder(16#1c#)) OR
 					(reg_q876 AND symb_decoder(16#70#)) OR
 					(reg_q876 AND symb_decoder(16#2e#)) OR
 					(reg_q876 AND symb_decoder(16#dc#)) OR
 					(reg_q876 AND symb_decoder(16#ce#)) OR
 					(reg_q876 AND symb_decoder(16#c0#)) OR
 					(reg_q876 AND symb_decoder(16#09#)) OR
 					(reg_q876 AND symb_decoder(16#07#)) OR
 					(reg_q876 AND symb_decoder(16#2d#)) OR
 					(reg_q876 AND symb_decoder(16#7f#)) OR
 					(reg_q876 AND symb_decoder(16#47#)) OR
 					(reg_q876 AND symb_decoder(16#aa#)) OR
 					(reg_q876 AND symb_decoder(16#53#)) OR
 					(reg_q876 AND symb_decoder(16#ac#)) OR
 					(reg_q876 AND symb_decoder(16#43#)) OR
 					(reg_q876 AND symb_decoder(16#3b#)) OR
 					(reg_q876 AND symb_decoder(16#cd#)) OR
 					(reg_q876 AND symb_decoder(16#c5#)) OR
 					(reg_q876 AND symb_decoder(16#60#)) OR
 					(reg_q876 AND symb_decoder(16#3a#)) OR
 					(reg_q876 AND symb_decoder(16#db#)) OR
 					(reg_q876 AND symb_decoder(16#57#)) OR
 					(reg_q876 AND symb_decoder(16#9f#)) OR
 					(reg_q876 AND symb_decoder(16#fc#)) OR
 					(reg_q876 AND symb_decoder(16#55#)) OR
 					(reg_q876 AND symb_decoder(16#6a#)) OR
 					(reg_q876 AND symb_decoder(16#f8#)) OR
 					(reg_q876 AND symb_decoder(16#06#)) OR
 					(reg_q876 AND symb_decoder(16#48#)) OR
 					(reg_q876 AND symb_decoder(16#df#)) OR
 					(reg_q876 AND symb_decoder(16#59#)) OR
 					(reg_q876 AND symb_decoder(16#44#)) OR
 					(reg_q876 AND symb_decoder(16#67#)) OR
 					(reg_q876 AND symb_decoder(16#52#)) OR
 					(reg_q876 AND symb_decoder(16#af#)) OR
 					(reg_q876 AND symb_decoder(16#42#)) OR
 					(reg_q876 AND symb_decoder(16#de#)) OR
 					(reg_q876 AND symb_decoder(16#1f#)) OR
 					(reg_q876 AND symb_decoder(16#e7#)) OR
 					(reg_q876 AND symb_decoder(16#54#)) OR
 					(reg_q876 AND symb_decoder(16#f3#)) OR
 					(reg_q876 AND symb_decoder(16#fa#)) OR
 					(reg_q876 AND symb_decoder(16#ab#)) OR
 					(reg_q876 AND symb_decoder(16#7c#)) OR
 					(reg_q876 AND symb_decoder(16#f0#)) OR
 					(reg_q876 AND symb_decoder(16#64#)) OR
 					(reg_q876 AND symb_decoder(16#5d#)) OR
 					(reg_q876 AND symb_decoder(16#e9#)) OR
 					(reg_q876 AND symb_decoder(16#a7#)) OR
 					(reg_q876 AND symb_decoder(16#18#)) OR
 					(reg_q876 AND symb_decoder(16#a1#)) OR
 					(reg_q876 AND symb_decoder(16#ca#)) OR
 					(reg_q876 AND symb_decoder(16#45#)) OR
 					(reg_q876 AND symb_decoder(16#65#)) OR
 					(reg_q876 AND symb_decoder(16#8c#)) OR
 					(reg_q876 AND symb_decoder(16#28#)) OR
 					(reg_q876 AND symb_decoder(16#5c#)) OR
 					(reg_q876 AND symb_decoder(16#2f#)) OR
 					(reg_q876 AND symb_decoder(16#8a#)) OR
 					(reg_q876 AND symb_decoder(16#7b#)) OR
 					(reg_q876 AND symb_decoder(16#8e#)) OR
 					(reg_q876 AND symb_decoder(16#7d#)) OR
 					(reg_q876 AND symb_decoder(16#99#)) OR
 					(reg_q876 AND symb_decoder(16#62#)) OR
 					(reg_q876 AND symb_decoder(16#b4#)) OR
 					(reg_q876 AND symb_decoder(16#e0#)) OR
 					(reg_q876 AND symb_decoder(16#0f#)) OR
 					(reg_q876 AND symb_decoder(16#33#)) OR
 					(reg_q876 AND symb_decoder(16#24#)) OR
 					(reg_q876 AND symb_decoder(16#9e#)) OR
 					(reg_q876 AND symb_decoder(16#b1#)) OR
 					(reg_q876 AND symb_decoder(16#a2#)) OR
 					(reg_q876 AND symb_decoder(16#5b#)) OR
 					(reg_q876 AND symb_decoder(16#a8#)) OR
 					(reg_q942 AND symb_decoder(16#a0#)) OR
 					(reg_q942 AND symb_decoder(16#f5#)) OR
 					(reg_q942 AND symb_decoder(16#60#)) OR
 					(reg_q942 AND symb_decoder(16#8f#)) OR
 					(reg_q942 AND symb_decoder(16#1f#)) OR
 					(reg_q942 AND symb_decoder(16#7b#)) OR
 					(reg_q942 AND symb_decoder(16#18#)) OR
 					(reg_q942 AND symb_decoder(16#ef#)) OR
 					(reg_q942 AND symb_decoder(16#f2#)) OR
 					(reg_q942 AND symb_decoder(16#6d#)) OR
 					(reg_q942 AND symb_decoder(16#36#)) OR
 					(reg_q942 AND symb_decoder(16#24#)) OR
 					(reg_q942 AND symb_decoder(16#a3#)) OR
 					(reg_q942 AND symb_decoder(16#5d#)) OR
 					(reg_q942 AND symb_decoder(16#34#)) OR
 					(reg_q942 AND symb_decoder(16#cb#)) OR
 					(reg_q942 AND symb_decoder(16#c8#)) OR
 					(reg_q942 AND symb_decoder(16#e3#)) OR
 					(reg_q942 AND symb_decoder(16#8a#)) OR
 					(reg_q942 AND symb_decoder(16#cc#)) OR
 					(reg_q942 AND symb_decoder(16#d2#)) OR
 					(reg_q942 AND symb_decoder(16#4a#)) OR
 					(reg_q942 AND symb_decoder(16#6e#)) OR
 					(reg_q942 AND symb_decoder(16#ed#)) OR
 					(reg_q942 AND symb_decoder(16#01#)) OR
 					(reg_q942 AND symb_decoder(16#d8#)) OR
 					(reg_q942 AND symb_decoder(16#e5#)) OR
 					(reg_q942 AND symb_decoder(16#47#)) OR
 					(reg_q942 AND symb_decoder(16#98#)) OR
 					(reg_q942 AND symb_decoder(16#2d#)) OR
 					(reg_q942 AND symb_decoder(16#6a#)) OR
 					(reg_q942 AND symb_decoder(16#17#)) OR
 					(reg_q942 AND symb_decoder(16#fd#)) OR
 					(reg_q942 AND symb_decoder(16#d9#)) OR
 					(reg_q942 AND symb_decoder(16#d5#)) OR
 					(reg_q942 AND symb_decoder(16#8d#)) OR
 					(reg_q942 AND symb_decoder(16#c2#)) OR
 					(reg_q942 AND symb_decoder(16#12#)) OR
 					(reg_q942 AND symb_decoder(16#67#)) OR
 					(reg_q942 AND symb_decoder(16#c7#)) OR
 					(reg_q942 AND symb_decoder(16#b6#)) OR
 					(reg_q942 AND symb_decoder(16#ce#)) OR
 					(reg_q942 AND symb_decoder(16#04#)) OR
 					(reg_q942 AND symb_decoder(16#f4#)) OR
 					(reg_q942 AND symb_decoder(16#84#)) OR
 					(reg_q942 AND symb_decoder(16#1d#)) OR
 					(reg_q942 AND symb_decoder(16#26#)) OR
 					(reg_q942 AND symb_decoder(16#29#)) OR
 					(reg_q942 AND symb_decoder(16#21#)) OR
 					(reg_q942 AND symb_decoder(16#fc#)) OR
 					(reg_q942 AND symb_decoder(16#2e#)) OR
 					(reg_q942 AND symb_decoder(16#37#)) OR
 					(reg_q942 AND symb_decoder(16#bd#)) OR
 					(reg_q942 AND symb_decoder(16#10#)) OR
 					(reg_q942 AND symb_decoder(16#ca#)) OR
 					(reg_q942 AND symb_decoder(16#bc#)) OR
 					(reg_q942 AND symb_decoder(16#da#)) OR
 					(reg_q942 AND symb_decoder(16#73#)) OR
 					(reg_q942 AND symb_decoder(16#a9#)) OR
 					(reg_q942 AND symb_decoder(16#d6#)) OR
 					(reg_q942 AND symb_decoder(16#b1#)) OR
 					(reg_q942 AND symb_decoder(16#2a#)) OR
 					(reg_q942 AND symb_decoder(16#e2#)) OR
 					(reg_q942 AND symb_decoder(16#4e#)) OR
 					(reg_q942 AND symb_decoder(16#02#)) OR
 					(reg_q942 AND symb_decoder(16#3e#)) OR
 					(reg_q942 AND symb_decoder(16#6b#)) OR
 					(reg_q942 AND symb_decoder(16#2c#)) OR
 					(reg_q942 AND symb_decoder(16#fe#)) OR
 					(reg_q942 AND symb_decoder(16#6c#)) OR
 					(reg_q942 AND symb_decoder(16#97#)) OR
 					(reg_q942 AND symb_decoder(16#ae#)) OR
 					(reg_q942 AND symb_decoder(16#aa#)) OR
 					(reg_q942 AND symb_decoder(16#55#)) OR
 					(reg_q942 AND symb_decoder(16#bb#)) OR
 					(reg_q942 AND symb_decoder(16#c9#)) OR
 					(reg_q942 AND symb_decoder(16#c3#)) OR
 					(reg_q942 AND symb_decoder(16#a5#)) OR
 					(reg_q942 AND symb_decoder(16#15#)) OR
 					(reg_q942 AND symb_decoder(16#58#)) OR
 					(reg_q942 AND symb_decoder(16#c0#)) OR
 					(reg_q942 AND symb_decoder(16#7f#)) OR
 					(reg_q942 AND symb_decoder(16#7a#)) OR
 					(reg_q942 AND symb_decoder(16#89#)) OR
 					(reg_q942 AND symb_decoder(16#b8#)) OR
 					(reg_q942 AND symb_decoder(16#ba#)) OR
 					(reg_q942 AND symb_decoder(16#43#)) OR
 					(reg_q942 AND symb_decoder(16#dc#)) OR
 					(reg_q942 AND symb_decoder(16#54#)) OR
 					(reg_q942 AND symb_decoder(16#72#)) OR
 					(reg_q942 AND symb_decoder(16#61#)) OR
 					(reg_q942 AND symb_decoder(16#9a#)) OR
 					(reg_q942 AND symb_decoder(16#45#)) OR
 					(reg_q942 AND symb_decoder(16#82#)) OR
 					(reg_q942 AND symb_decoder(16#0c#)) OR
 					(reg_q942 AND symb_decoder(16#80#)) OR
 					(reg_q942 AND symb_decoder(16#b4#)) OR
 					(reg_q942 AND symb_decoder(16#f3#)) OR
 					(reg_q942 AND symb_decoder(16#32#)) OR
 					(reg_q942 AND symb_decoder(16#dd#)) OR
 					(reg_q942 AND symb_decoder(16#e9#)) OR
 					(reg_q942 AND symb_decoder(16#ad#)) OR
 					(reg_q942 AND symb_decoder(16#f9#)) OR
 					(reg_q942 AND symb_decoder(16#06#)) OR
 					(reg_q942 AND symb_decoder(16#d4#)) OR
 					(reg_q942 AND symb_decoder(16#d7#)) OR
 					(reg_q942 AND symb_decoder(16#38#)) OR
 					(reg_q942 AND symb_decoder(16#91#)) OR
 					(reg_q942 AND symb_decoder(16#42#)) OR
 					(reg_q942 AND symb_decoder(16#9f#)) OR
 					(reg_q942 AND symb_decoder(16#08#)) OR
 					(reg_q942 AND symb_decoder(16#77#)) OR
 					(reg_q942 AND symb_decoder(16#05#)) OR
 					(reg_q942 AND symb_decoder(16#b9#)) OR
 					(reg_q942 AND symb_decoder(16#40#)) OR
 					(reg_q942 AND symb_decoder(16#50#)) OR
 					(reg_q942 AND symb_decoder(16#78#)) OR
 					(reg_q942 AND symb_decoder(16#1a#)) OR
 					(reg_q942 AND symb_decoder(16#71#)) OR
 					(reg_q942 AND symb_decoder(16#e0#)) OR
 					(reg_q942 AND symb_decoder(16#11#)) OR
 					(reg_q942 AND symb_decoder(16#2b#)) OR
 					(reg_q942 AND symb_decoder(16#86#)) OR
 					(reg_q942 AND symb_decoder(16#62#)) OR
 					(reg_q942 AND symb_decoder(16#9d#)) OR
 					(reg_q942 AND symb_decoder(16#a7#)) OR
 					(reg_q942 AND symb_decoder(16#63#)) OR
 					(reg_q942 AND symb_decoder(16#76#)) OR
 					(reg_q942 AND symb_decoder(16#b3#)) OR
 					(reg_q942 AND symb_decoder(16#81#)) OR
 					(reg_q942 AND symb_decoder(16#c4#)) OR
 					(reg_q942 AND symb_decoder(16#4c#)) OR
 					(reg_q942 AND symb_decoder(16#3a#)) OR
 					(reg_q942 AND symb_decoder(16#ec#)) OR
 					(reg_q942 AND symb_decoder(16#7e#)) OR
 					(reg_q942 AND symb_decoder(16#13#)) OR
 					(reg_q942 AND symb_decoder(16#ab#)) OR
 					(reg_q942 AND symb_decoder(16#3f#)) OR
 					(reg_q942 AND symb_decoder(16#23#)) OR
 					(reg_q942 AND symb_decoder(16#1e#)) OR
 					(reg_q942 AND symb_decoder(16#fb#)) OR
 					(reg_q942 AND symb_decoder(16#f6#)) OR
 					(reg_q942 AND symb_decoder(16#20#)) OR
 					(reg_q942 AND symb_decoder(16#c5#)) OR
 					(reg_q942 AND symb_decoder(16#6f#)) OR
 					(reg_q942 AND symb_decoder(16#5f#)) OR
 					(reg_q942 AND symb_decoder(16#96#)) OR
 					(reg_q942 AND symb_decoder(16#b2#)) OR
 					(reg_q942 AND symb_decoder(16#c6#)) OR
 					(reg_q942 AND symb_decoder(16#de#)) OR
 					(reg_q942 AND symb_decoder(16#16#)) OR
 					(reg_q942 AND symb_decoder(16#2f#)) OR
 					(reg_q942 AND symb_decoder(16#a1#)) OR
 					(reg_q942 AND symb_decoder(16#79#)) OR
 					(reg_q942 AND symb_decoder(16#8c#)) OR
 					(reg_q942 AND symb_decoder(16#5b#)) OR
 					(reg_q942 AND symb_decoder(16#53#)) OR
 					(reg_q942 AND symb_decoder(16#df#)) OR
 					(reg_q942 AND symb_decoder(16#4b#)) OR
 					(reg_q942 AND symb_decoder(16#00#)) OR
 					(reg_q942 AND symb_decoder(16#14#)) OR
 					(reg_q942 AND symb_decoder(16#5a#)) OR
 					(reg_q942 AND symb_decoder(16#3c#)) OR
 					(reg_q942 AND symb_decoder(16#ea#)) OR
 					(reg_q942 AND symb_decoder(16#25#)) OR
 					(reg_q942 AND symb_decoder(16#3d#)) OR
 					(reg_q942 AND symb_decoder(16#03#)) OR
 					(reg_q942 AND symb_decoder(16#66#)) OR
 					(reg_q942 AND symb_decoder(16#88#)) OR
 					(reg_q942 AND symb_decoder(16#56#)) OR
 					(reg_q942 AND symb_decoder(16#0b#)) OR
 					(reg_q942 AND symb_decoder(16#eb#)) OR
 					(reg_q942 AND symb_decoder(16#27#)) OR
 					(reg_q942 AND symb_decoder(16#f0#)) OR
 					(reg_q942 AND symb_decoder(16#09#)) OR
 					(reg_q942 AND symb_decoder(16#83#)) OR
 					(reg_q942 AND symb_decoder(16#d1#)) OR
 					(reg_q942 AND symb_decoder(16#93#)) OR
 					(reg_q942 AND symb_decoder(16#f8#)) OR
 					(reg_q942 AND symb_decoder(16#1c#)) OR
 					(reg_q942 AND symb_decoder(16#95#)) OR
 					(reg_q942 AND symb_decoder(16#ff#)) OR
 					(reg_q942 AND symb_decoder(16#a6#)) OR
 					(reg_q942 AND symb_decoder(16#90#)) OR
 					(reg_q942 AND symb_decoder(16#b7#)) OR
 					(reg_q942 AND symb_decoder(16#4d#)) OR
 					(reg_q942 AND symb_decoder(16#68#)) OR
 					(reg_q942 AND symb_decoder(16#8e#)) OR
 					(reg_q942 AND symb_decoder(16#d0#)) OR
 					(reg_q942 AND symb_decoder(16#a2#)) OR
 					(reg_q942 AND symb_decoder(16#4f#)) OR
 					(reg_q942 AND symb_decoder(16#41#)) OR
 					(reg_q942 AND symb_decoder(16#64#)) OR
 					(reg_q942 AND symb_decoder(16#28#)) OR
 					(reg_q942 AND symb_decoder(16#bf#)) OR
 					(reg_q942 AND symb_decoder(16#69#)) OR
 					(reg_q942 AND symb_decoder(16#7c#)) OR
 					(reg_q942 AND symb_decoder(16#5e#)) OR
 					(reg_q942 AND symb_decoder(16#0e#)) OR
 					(reg_q942 AND symb_decoder(16#7d#)) OR
 					(reg_q942 AND symb_decoder(16#b0#)) OR
 					(reg_q942 AND symb_decoder(16#94#)) OR
 					(reg_q942 AND symb_decoder(16#51#)) OR
 					(reg_q942 AND symb_decoder(16#a8#)) OR
 					(reg_q942 AND symb_decoder(16#af#)) OR
 					(reg_q942 AND symb_decoder(16#92#)) OR
 					(reg_q942 AND symb_decoder(16#35#)) OR
 					(reg_q942 AND symb_decoder(16#f7#)) OR
 					(reg_q942 AND symb_decoder(16#44#)) OR
 					(reg_q942 AND symb_decoder(16#ac#)) OR
 					(reg_q942 AND symb_decoder(16#1b#)) OR
 					(reg_q942 AND symb_decoder(16#87#)) OR
 					(reg_q942 AND symb_decoder(16#46#)) OR
 					(reg_q942 AND symb_decoder(16#5c#)) OR
 					(reg_q942 AND symb_decoder(16#85#)) OR
 					(reg_q942 AND symb_decoder(16#e1#)) OR
 					(reg_q942 AND symb_decoder(16#33#)) OR
 					(reg_q942 AND symb_decoder(16#cf#)) OR
 					(reg_q942 AND symb_decoder(16#39#)) OR
 					(reg_q942 AND symb_decoder(16#49#)) OR
 					(reg_q942 AND symb_decoder(16#30#)) OR
 					(reg_q942 AND symb_decoder(16#fa#)) OR
 					(reg_q942 AND symb_decoder(16#57#)) OR
 					(reg_q942 AND symb_decoder(16#9c#)) OR
 					(reg_q942 AND symb_decoder(16#c1#)) OR
 					(reg_q942 AND symb_decoder(16#e8#)) OR
 					(reg_q942 AND symb_decoder(16#e7#)) OR
 					(reg_q942 AND symb_decoder(16#ee#)) OR
 					(reg_q942 AND symb_decoder(16#9e#)) OR
 					(reg_q942 AND symb_decoder(16#db#)) OR
 					(reg_q942 AND symb_decoder(16#19#)) OR
 					(reg_q942 AND symb_decoder(16#75#)) OR
 					(reg_q942 AND symb_decoder(16#8b#)) OR
 					(reg_q942 AND symb_decoder(16#cd#)) OR
 					(reg_q942 AND symb_decoder(16#74#)) OR
 					(reg_q942 AND symb_decoder(16#52#)) OR
 					(reg_q942 AND symb_decoder(16#70#)) OR
 					(reg_q942 AND symb_decoder(16#0f#)) OR
 					(reg_q942 AND symb_decoder(16#31#)) OR
 					(reg_q942 AND symb_decoder(16#a4#)) OR
 					(reg_q942 AND symb_decoder(16#e6#)) OR
 					(reg_q942 AND symb_decoder(16#be#)) OR
 					(reg_q942 AND symb_decoder(16#9b#)) OR
 					(reg_q942 AND symb_decoder(16#e4#)) OR
 					(reg_q942 AND symb_decoder(16#65#)) OR
 					(reg_q942 AND symb_decoder(16#d3#)) OR
 					(reg_q942 AND symb_decoder(16#22#)) OR
 					(reg_q942 AND symb_decoder(16#3b#)) OR
 					(reg_q942 AND symb_decoder(16#48#)) OR
 					(reg_q942 AND symb_decoder(16#f1#)) OR
 					(reg_q942 AND symb_decoder(16#07#)) OR
 					(reg_q942 AND symb_decoder(16#99#)) OR
 					(reg_q942 AND symb_decoder(16#b5#)) OR
 					(reg_q942 AND symb_decoder(16#59#));
reg_q2524_in <= (reg_q2522 AND symb_decoder(16#41#)) OR
 					(reg_q2522 AND symb_decoder(16#61#));
reg_q359_in <= (reg_q357 AND symb_decoder(16#3a#));
reg_q2034_in <= (reg_q2032 AND symb_decoder(16#61#)) OR
 					(reg_q2032 AND symb_decoder(16#35#)) OR
 					(reg_q2032 AND symb_decoder(16#44#)) OR
 					(reg_q2032 AND symb_decoder(16#38#)) OR
 					(reg_q2032 AND symb_decoder(16#46#)) OR
 					(reg_q2032 AND symb_decoder(16#32#)) OR
 					(reg_q2032 AND symb_decoder(16#30#)) OR
 					(reg_q2032 AND symb_decoder(16#36#)) OR
 					(reg_q2032 AND symb_decoder(16#63#)) OR
 					(reg_q2032 AND symb_decoder(16#42#)) OR
 					(reg_q2032 AND symb_decoder(16#62#)) OR
 					(reg_q2032 AND symb_decoder(16#43#)) OR
 					(reg_q2032 AND symb_decoder(16#65#)) OR
 					(reg_q2032 AND symb_decoder(16#34#)) OR
 					(reg_q2032 AND symb_decoder(16#37#)) OR
 					(reg_q2032 AND symb_decoder(16#64#)) OR
 					(reg_q2032 AND symb_decoder(16#41#)) OR
 					(reg_q2032 AND symb_decoder(16#39#)) OR
 					(reg_q2032 AND symb_decoder(16#33#)) OR
 					(reg_q2032 AND symb_decoder(16#66#)) OR
 					(reg_q2032 AND symb_decoder(16#45#)) OR
 					(reg_q2032 AND symb_decoder(16#31#));
reg_q2036_in <= (reg_q2034 AND symb_decoder(16#33#)) OR
 					(reg_q2034 AND symb_decoder(16#30#)) OR
 					(reg_q2034 AND symb_decoder(16#39#)) OR
 					(reg_q2034 AND symb_decoder(16#46#)) OR
 					(reg_q2034 AND symb_decoder(16#36#)) OR
 					(reg_q2034 AND symb_decoder(16#34#)) OR
 					(reg_q2034 AND symb_decoder(16#64#)) OR
 					(reg_q2034 AND symb_decoder(16#32#)) OR
 					(reg_q2034 AND symb_decoder(16#61#)) OR
 					(reg_q2034 AND symb_decoder(16#43#)) OR
 					(reg_q2034 AND symb_decoder(16#31#)) OR
 					(reg_q2034 AND symb_decoder(16#41#)) OR
 					(reg_q2034 AND symb_decoder(16#44#)) OR
 					(reg_q2034 AND symb_decoder(16#62#)) OR
 					(reg_q2034 AND symb_decoder(16#38#)) OR
 					(reg_q2034 AND symb_decoder(16#66#)) OR
 					(reg_q2034 AND symb_decoder(16#35#)) OR
 					(reg_q2034 AND symb_decoder(16#37#)) OR
 					(reg_q2034 AND symb_decoder(16#45#)) OR
 					(reg_q2034 AND symb_decoder(16#65#)) OR
 					(reg_q2034 AND symb_decoder(16#63#)) OR
 					(reg_q2034 AND symb_decoder(16#42#));
reg_q2623_in <= (reg_q2623 AND symb_decoder(16#33#)) OR
 					(reg_q2623 AND symb_decoder(16#37#)) OR
 					(reg_q2623 AND symb_decoder(16#31#)) OR
 					(reg_q2623 AND symb_decoder(16#36#)) OR
 					(reg_q2623 AND symb_decoder(16#34#)) OR
 					(reg_q2623 AND symb_decoder(16#35#)) OR
 					(reg_q2623 AND symb_decoder(16#32#)) OR
 					(reg_q2623 AND symb_decoder(16#30#)) OR
 					(reg_q2623 AND symb_decoder(16#39#)) OR
 					(reg_q2623 AND symb_decoder(16#38#)) OR
 					(reg_q2621 AND symb_decoder(16#36#)) OR
 					(reg_q2621 AND symb_decoder(16#35#)) OR
 					(reg_q2621 AND symb_decoder(16#32#)) OR
 					(reg_q2621 AND symb_decoder(16#30#)) OR
 					(reg_q2621 AND symb_decoder(16#37#)) OR
 					(reg_q2621 AND symb_decoder(16#39#)) OR
 					(reg_q2621 AND symb_decoder(16#33#)) OR
 					(reg_q2621 AND symb_decoder(16#34#)) OR
 					(reg_q2621 AND symb_decoder(16#38#)) OR
 					(reg_q2621 AND symb_decoder(16#31#));
reg_q675_in <= (reg_q675 AND symb_decoder(16#33#)) OR
 					(reg_q675 AND symb_decoder(16#30#)) OR
 					(reg_q675 AND symb_decoder(16#37#)) OR
 					(reg_q675 AND symb_decoder(16#34#)) OR
 					(reg_q675 AND symb_decoder(16#35#)) OR
 					(reg_q675 AND symb_decoder(16#31#)) OR
 					(reg_q675 AND symb_decoder(16#32#)) OR
 					(reg_q675 AND symb_decoder(16#39#)) OR
 					(reg_q675 AND symb_decoder(16#38#)) OR
 					(reg_q675 AND symb_decoder(16#36#)) OR
 					(reg_q673 AND symb_decoder(16#35#)) OR
 					(reg_q673 AND symb_decoder(16#34#)) OR
 					(reg_q673 AND symb_decoder(16#30#)) OR
 					(reg_q673 AND symb_decoder(16#38#)) OR
 					(reg_q673 AND symb_decoder(16#37#)) OR
 					(reg_q673 AND symb_decoder(16#36#)) OR
 					(reg_q673 AND symb_decoder(16#33#)) OR
 					(reg_q673 AND symb_decoder(16#39#)) OR
 					(reg_q673 AND symb_decoder(16#32#)) OR
 					(reg_q673 AND symb_decoder(16#31#));
reg_q149_in <= (reg_q147 AND symb_decoder(16#72#)) OR
 					(reg_q147 AND symb_decoder(16#52#));
reg_q151_in <= (reg_q149 AND symb_decoder(16#0c#)) OR
 					(reg_q149 AND symb_decoder(16#20#)) OR
 					(reg_q149 AND symb_decoder(16#09#)) OR
 					(reg_q149 AND symb_decoder(16#0a#)) OR
 					(reg_q149 AND symb_decoder(16#0d#)) OR
 					(reg_q151 AND symb_decoder(16#0a#)) OR
 					(reg_q151 AND symb_decoder(16#0c#)) OR
 					(reg_q151 AND symb_decoder(16#09#)) OR
 					(reg_q151 AND symb_decoder(16#0d#)) OR
 					(reg_q151 AND symb_decoder(16#20#));
reg_q480_in <= (reg_q478 AND symb_decoder(16#3a#));
reg_q40_in <= (reg_q40 AND symb_decoder(16#0d#)) OR
 					(reg_q40 AND symb_decoder(16#09#)) OR
 					(reg_q40 AND symb_decoder(16#0a#)) OR
 					(reg_q40 AND symb_decoder(16#0c#)) OR
 					(reg_q40 AND symb_decoder(16#20#)) OR
 					(reg_q38 AND symb_decoder(16#0a#)) OR
 					(reg_q38 AND symb_decoder(16#20#)) OR
 					(reg_q38 AND symb_decoder(16#09#)) OR
 					(reg_q38 AND symb_decoder(16#0c#)) OR
 					(reg_q38 AND symb_decoder(16#0d#));
reg_q732_in <= (reg_q732 AND symb_decoder(16#20#)) OR
 					(reg_q732 AND symb_decoder(16#0c#)) OR
 					(reg_q732 AND symb_decoder(16#0a#)) OR
 					(reg_q732 AND symb_decoder(16#0d#)) OR
 					(reg_q732 AND symb_decoder(16#09#)) OR
 					(reg_q730 AND symb_decoder(16#09#)) OR
 					(reg_q730 AND symb_decoder(16#0a#)) OR
 					(reg_q730 AND symb_decoder(16#0d#)) OR
 					(reg_q730 AND symb_decoder(16#20#)) OR
 					(reg_q730 AND symb_decoder(16#0c#));
reg_q1357_in <= (reg_q1355 AND symb_decoder(16#4e#)) OR
 					(reg_q1355 AND symb_decoder(16#6e#));
reg_q107_in <= (reg_q107 AND symb_decoder(16#0c#)) OR
 					(reg_q107 AND symb_decoder(16#0d#)) OR
 					(reg_q107 AND symb_decoder(16#20#)) OR
 					(reg_q107 AND symb_decoder(16#09#)) OR
 					(reg_q107 AND symb_decoder(16#0a#)) OR
 					(reg_q105 AND symb_decoder(16#0a#)) OR
 					(reg_q105 AND symb_decoder(16#0d#)) OR
 					(reg_q105 AND symb_decoder(16#20#)) OR
 					(reg_q105 AND symb_decoder(16#09#)) OR
 					(reg_q105 AND symb_decoder(16#0c#));
reg_q2290_in <= (reg_q2290 AND symb_decoder(16#0d#)) OR
 					(reg_q2290 AND symb_decoder(16#0a#)) OR
 					(reg_q2290 AND symb_decoder(16#0c#)) OR
 					(reg_q2290 AND symb_decoder(16#20#)) OR
 					(reg_q2290 AND symb_decoder(16#09#)) OR
 					(reg_q2288 AND symb_decoder(16#0a#)) OR
 					(reg_q2288 AND symb_decoder(16#09#)) OR
 					(reg_q2288 AND symb_decoder(16#20#)) OR
 					(reg_q2288 AND symb_decoder(16#0d#)) OR
 					(reg_q2288 AND symb_decoder(16#0c#));
reg_q2312_in <= (reg_q2312 AND symb_decoder(16#09#)) OR
 					(reg_q2312 AND symb_decoder(16#0c#)) OR
 					(reg_q2312 AND symb_decoder(16#0d#)) OR
 					(reg_q2312 AND symb_decoder(16#0a#)) OR
 					(reg_q2312 AND symb_decoder(16#20#)) OR
 					(reg_q2310 AND symb_decoder(16#09#)) OR
 					(reg_q2310 AND symb_decoder(16#0d#)) OR
 					(reg_q2310 AND symb_decoder(16#20#)) OR
 					(reg_q2310 AND symb_decoder(16#0a#)) OR
 					(reg_q2310 AND symb_decoder(16#0c#));
reg_q2314_in <= (reg_q2312 AND symb_decoder(16#55#)) OR
 					(reg_q2312 AND symb_decoder(16#75#));
reg_q2038_in <= (reg_q2036 AND symb_decoder(16#66#)) OR
 					(reg_q2036 AND symb_decoder(16#45#)) OR
 					(reg_q2036 AND symb_decoder(16#62#)) OR
 					(reg_q2036 AND symb_decoder(16#64#)) OR
 					(reg_q2036 AND symb_decoder(16#30#)) OR
 					(reg_q2036 AND symb_decoder(16#35#)) OR
 					(reg_q2036 AND symb_decoder(16#42#)) OR
 					(reg_q2036 AND symb_decoder(16#31#)) OR
 					(reg_q2036 AND symb_decoder(16#34#)) OR
 					(reg_q2036 AND symb_decoder(16#37#)) OR
 					(reg_q2036 AND symb_decoder(16#44#)) OR
 					(reg_q2036 AND symb_decoder(16#65#)) OR
 					(reg_q2036 AND symb_decoder(16#32#)) OR
 					(reg_q2036 AND symb_decoder(16#63#)) OR
 					(reg_q2036 AND symb_decoder(16#43#)) OR
 					(reg_q2036 AND symb_decoder(16#36#)) OR
 					(reg_q2036 AND symb_decoder(16#61#)) OR
 					(reg_q2036 AND symb_decoder(16#46#)) OR
 					(reg_q2036 AND symb_decoder(16#38#)) OR
 					(reg_q2036 AND symb_decoder(16#39#)) OR
 					(reg_q2036 AND symb_decoder(16#33#)) OR
 					(reg_q2036 AND symb_decoder(16#41#));
reg_q1502_in <= (reg_q1500 AND symb_decoder(16#73#)) OR
 					(reg_q1500 AND symb_decoder(16#53#));
reg_q1504_in <= (reg_q1502 AND symb_decoder(16#45#)) OR
 					(reg_q1502 AND symb_decoder(16#65#));
reg_q1996_in <= (reg_q1994 AND symb_decoder(16#30#)) OR
 					(reg_q1994 AND symb_decoder(16#61#)) OR
 					(reg_q1994 AND symb_decoder(16#32#)) OR
 					(reg_q1994 AND symb_decoder(16#66#)) OR
 					(reg_q1994 AND symb_decoder(16#34#)) OR
 					(reg_q1994 AND symb_decoder(16#62#)) OR
 					(reg_q1994 AND symb_decoder(16#36#)) OR
 					(reg_q1994 AND symb_decoder(16#38#)) OR
 					(reg_q1994 AND symb_decoder(16#65#)) OR
 					(reg_q1994 AND symb_decoder(16#41#)) OR
 					(reg_q1994 AND symb_decoder(16#64#)) OR
 					(reg_q1994 AND symb_decoder(16#45#)) OR
 					(reg_q1994 AND symb_decoder(16#43#)) OR
 					(reg_q1994 AND symb_decoder(16#37#)) OR
 					(reg_q1994 AND symb_decoder(16#63#)) OR
 					(reg_q1994 AND symb_decoder(16#31#)) OR
 					(reg_q1994 AND symb_decoder(16#44#)) OR
 					(reg_q1994 AND symb_decoder(16#46#)) OR
 					(reg_q1994 AND symb_decoder(16#42#)) OR
 					(reg_q1994 AND symb_decoder(16#39#)) OR
 					(reg_q1994 AND symb_decoder(16#35#)) OR
 					(reg_q1994 AND symb_decoder(16#33#));
reg_q1998_in <= (reg_q1996 AND symb_decoder(16#33#)) OR
 					(reg_q1996 AND symb_decoder(16#35#)) OR
 					(reg_q1996 AND symb_decoder(16#46#)) OR
 					(reg_q1996 AND symb_decoder(16#65#)) OR
 					(reg_q1996 AND symb_decoder(16#37#)) OR
 					(reg_q1996 AND symb_decoder(16#62#)) OR
 					(reg_q1996 AND symb_decoder(16#61#)) OR
 					(reg_q1996 AND symb_decoder(16#36#)) OR
 					(reg_q1996 AND symb_decoder(16#30#)) OR
 					(reg_q1996 AND symb_decoder(16#39#)) OR
 					(reg_q1996 AND symb_decoder(16#63#)) OR
 					(reg_q1996 AND symb_decoder(16#38#)) OR
 					(reg_q1996 AND symb_decoder(16#31#)) OR
 					(reg_q1996 AND symb_decoder(16#32#)) OR
 					(reg_q1996 AND symb_decoder(16#41#)) OR
 					(reg_q1996 AND symb_decoder(16#64#)) OR
 					(reg_q1996 AND symb_decoder(16#44#)) OR
 					(reg_q1996 AND symb_decoder(16#43#)) OR
 					(reg_q1996 AND symb_decoder(16#42#)) OR
 					(reg_q1996 AND symb_decoder(16#45#)) OR
 					(reg_q1996 AND symb_decoder(16#66#)) OR
 					(reg_q1996 AND symb_decoder(16#34#));
reg_q2006_in <= (reg_q2004 AND symb_decoder(16#65#)) OR
 					(reg_q2004 AND symb_decoder(16#63#)) OR
 					(reg_q2004 AND symb_decoder(16#33#)) OR
 					(reg_q2004 AND symb_decoder(16#42#)) OR
 					(reg_q2004 AND symb_decoder(16#41#)) OR
 					(reg_q2004 AND symb_decoder(16#45#)) OR
 					(reg_q2004 AND symb_decoder(16#30#)) OR
 					(reg_q2004 AND symb_decoder(16#35#)) OR
 					(reg_q2004 AND symb_decoder(16#61#)) OR
 					(reg_q2004 AND symb_decoder(16#66#)) OR
 					(reg_q2004 AND symb_decoder(16#34#)) OR
 					(reg_q2004 AND symb_decoder(16#44#)) OR
 					(reg_q2004 AND symb_decoder(16#38#)) OR
 					(reg_q2004 AND symb_decoder(16#43#)) OR
 					(reg_q2004 AND symb_decoder(16#62#)) OR
 					(reg_q2004 AND symb_decoder(16#32#)) OR
 					(reg_q2004 AND symb_decoder(16#31#)) OR
 					(reg_q2004 AND symb_decoder(16#39#)) OR
 					(reg_q2004 AND symb_decoder(16#37#)) OR
 					(reg_q2004 AND symb_decoder(16#46#)) OR
 					(reg_q2004 AND symb_decoder(16#64#)) OR
 					(reg_q2004 AND symb_decoder(16#36#));
reg_q2008_in <= (reg_q2006 AND symb_decoder(16#43#)) OR
 					(reg_q2006 AND symb_decoder(16#63#)) OR
 					(reg_q2006 AND symb_decoder(16#38#)) OR
 					(reg_q2006 AND symb_decoder(16#33#)) OR
 					(reg_q2006 AND symb_decoder(16#36#)) OR
 					(reg_q2006 AND symb_decoder(16#31#)) OR
 					(reg_q2006 AND symb_decoder(16#66#)) OR
 					(reg_q2006 AND symb_decoder(16#39#)) OR
 					(reg_q2006 AND symb_decoder(16#62#)) OR
 					(reg_q2006 AND symb_decoder(16#32#)) OR
 					(reg_q2006 AND symb_decoder(16#65#)) OR
 					(reg_q2006 AND symb_decoder(16#61#)) OR
 					(reg_q2006 AND symb_decoder(16#37#)) OR
 					(reg_q2006 AND symb_decoder(16#44#)) OR
 					(reg_q2006 AND symb_decoder(16#34#)) OR
 					(reg_q2006 AND symb_decoder(16#64#)) OR
 					(reg_q2006 AND symb_decoder(16#30#)) OR
 					(reg_q2006 AND symb_decoder(16#41#)) OR
 					(reg_q2006 AND symb_decoder(16#35#)) OR
 					(reg_q2006 AND symb_decoder(16#46#)) OR
 					(reg_q2006 AND symb_decoder(16#42#)) OR
 					(reg_q2006 AND symb_decoder(16#45#));
reg_q817_in <= (reg_q815 AND symb_decoder(16#74#)) OR
 					(reg_q815 AND symb_decoder(16#54#));
reg_q1128_in <= (reg_q1126 AND symb_decoder(16#66#)) OR
 					(reg_q1126 AND symb_decoder(16#46#));
reg_q1130_in <= (reg_q1128 AND symb_decoder(16#69#)) OR
 					(reg_q1128 AND symb_decoder(16#49#));
reg_q2050_in <= (reg_q2048 AND symb_decoder(16#39#)) OR
 					(reg_q2048 AND symb_decoder(16#33#)) OR
 					(reg_q2048 AND symb_decoder(16#64#)) OR
 					(reg_q2048 AND symb_decoder(16#34#)) OR
 					(reg_q2048 AND symb_decoder(16#46#)) OR
 					(reg_q2048 AND symb_decoder(16#42#)) OR
 					(reg_q2048 AND symb_decoder(16#30#)) OR
 					(reg_q2048 AND symb_decoder(16#41#)) OR
 					(reg_q2048 AND symb_decoder(16#38#)) OR
 					(reg_q2048 AND symb_decoder(16#31#)) OR
 					(reg_q2048 AND symb_decoder(16#63#)) OR
 					(reg_q2048 AND symb_decoder(16#36#)) OR
 					(reg_q2048 AND symb_decoder(16#65#)) OR
 					(reg_q2048 AND symb_decoder(16#32#)) OR
 					(reg_q2048 AND symb_decoder(16#61#)) OR
 					(reg_q2048 AND symb_decoder(16#62#)) OR
 					(reg_q2048 AND symb_decoder(16#44#)) OR
 					(reg_q2048 AND symb_decoder(16#35#)) OR
 					(reg_q2048 AND symb_decoder(16#43#)) OR
 					(reg_q2048 AND symb_decoder(16#37#)) OR
 					(reg_q2048 AND symb_decoder(16#66#)) OR
 					(reg_q2048 AND symb_decoder(16#45#));
reg_q2054_in <= (reg_q2050 AND symb_decoder(16#64#)) OR
 					(reg_q2050 AND symb_decoder(16#37#)) OR
 					(reg_q2050 AND symb_decoder(16#44#)) OR
 					(reg_q2050 AND symb_decoder(16#61#)) OR
 					(reg_q2050 AND symb_decoder(16#35#)) OR
 					(reg_q2050 AND symb_decoder(16#39#)) OR
 					(reg_q2050 AND symb_decoder(16#38#)) OR
 					(reg_q2050 AND symb_decoder(16#30#)) OR
 					(reg_q2050 AND symb_decoder(16#32#)) OR
 					(reg_q2050 AND symb_decoder(16#46#)) OR
 					(reg_q2050 AND symb_decoder(16#45#)) OR
 					(reg_q2050 AND symb_decoder(16#33#)) OR
 					(reg_q2050 AND symb_decoder(16#65#)) OR
 					(reg_q2050 AND symb_decoder(16#42#)) OR
 					(reg_q2050 AND symb_decoder(16#63#)) OR
 					(reg_q2050 AND symb_decoder(16#34#)) OR
 					(reg_q2050 AND symb_decoder(16#36#)) OR
 					(reg_q2050 AND symb_decoder(16#41#)) OR
 					(reg_q2050 AND symb_decoder(16#66#)) OR
 					(reg_q2050 AND symb_decoder(16#31#)) OR
 					(reg_q2050 AND symb_decoder(16#62#)) OR
 					(reg_q2050 AND symb_decoder(16#43#)) OR
 					(reg_q2054 AND symb_decoder(16#43#)) OR
 					(reg_q2054 AND symb_decoder(16#35#)) OR
 					(reg_q2054 AND symb_decoder(16#64#)) OR
 					(reg_q2054 AND symb_decoder(16#63#)) OR
 					(reg_q2054 AND symb_decoder(16#62#)) OR
 					(reg_q2054 AND symb_decoder(16#34#)) OR
 					(reg_q2054 AND symb_decoder(16#32#)) OR
 					(reg_q2054 AND symb_decoder(16#66#)) OR
 					(reg_q2054 AND symb_decoder(16#44#)) OR
 					(reg_q2054 AND symb_decoder(16#38#)) OR
 					(reg_q2054 AND symb_decoder(16#42#)) OR
 					(reg_q2054 AND symb_decoder(16#39#)) OR
 					(reg_q2054 AND symb_decoder(16#46#)) OR
 					(reg_q2054 AND symb_decoder(16#30#)) OR
 					(reg_q2054 AND symb_decoder(16#33#)) OR
 					(reg_q2054 AND symb_decoder(16#41#)) OR
 					(reg_q2054 AND symb_decoder(16#36#)) OR
 					(reg_q2054 AND symb_decoder(16#45#)) OR
 					(reg_q2054 AND symb_decoder(16#61#)) OR
 					(reg_q2054 AND symb_decoder(16#37#)) OR
 					(reg_q2054 AND symb_decoder(16#31#)) OR
 					(reg_q2054 AND symb_decoder(16#65#));
reg_q210_in <= (reg_q210 AND symb_decoder(16#38#)) OR
 					(reg_q210 AND symb_decoder(16#34#)) OR
 					(reg_q210 AND symb_decoder(16#39#)) OR
 					(reg_q210 AND symb_decoder(16#35#)) OR
 					(reg_q210 AND symb_decoder(16#36#)) OR
 					(reg_q210 AND symb_decoder(16#31#)) OR
 					(reg_q210 AND symb_decoder(16#30#)) OR
 					(reg_q210 AND symb_decoder(16#37#)) OR
 					(reg_q210 AND symb_decoder(16#33#)) OR
 					(reg_q210 AND symb_decoder(16#32#)) OR
 					(reg_q208 AND symb_decoder(16#31#)) OR
 					(reg_q208 AND symb_decoder(16#33#)) OR
 					(reg_q208 AND symb_decoder(16#36#)) OR
 					(reg_q208 AND symb_decoder(16#35#)) OR
 					(reg_q208 AND symb_decoder(16#38#)) OR
 					(reg_q208 AND symb_decoder(16#34#)) OR
 					(reg_q208 AND symb_decoder(16#30#)) OR
 					(reg_q208 AND symb_decoder(16#37#)) OR
 					(reg_q208 AND symb_decoder(16#32#)) OR
 					(reg_q208 AND symb_decoder(16#39#));
reg_q369_in <= (reg_q367 AND symb_decoder(16#54#)) OR
 					(reg_q367 AND symb_decoder(16#74#));
reg_q712_in <= (reg_q710 AND symb_decoder(16#5c#));
reg_q714_in <= (reg_q712 AND symb_decoder(16#27#));
reg_q1924_in <= (reg_q1922 AND symb_decoder(16#52#));
reg_q1926_in <= (reg_q1924 AND symb_decoder(16#54#));
reg_q1709_in <= (reg_q1707 AND symb_decoder(16#6f#)) OR
 					(reg_q1707 AND symb_decoder(16#4f#));
reg_q1711_in <= (reg_q1709 AND symb_decoder(16#20#)) OR
 					(reg_q1709 AND symb_decoder(16#0d#)) OR
 					(reg_q1709 AND symb_decoder(16#0a#)) OR
 					(reg_q1709 AND symb_decoder(16#0c#)) OR
 					(reg_q1709 AND symb_decoder(16#09#)) OR
 					(reg_q1711 AND symb_decoder(16#0c#)) OR
 					(reg_q1711 AND symb_decoder(16#0a#)) OR
 					(reg_q1711 AND symb_decoder(16#20#)) OR
 					(reg_q1711 AND symb_decoder(16#09#)) OR
 					(reg_q1711 AND symb_decoder(16#0d#));
reg_q2280_in <= (reg_q2278 AND symb_decoder(16#77#)) OR
 					(reg_q2278 AND symb_decoder(16#57#));
reg_q2282_in <= (reg_q2280 AND symb_decoder(16#6e#)) OR
 					(reg_q2280 AND symb_decoder(16#4e#));
reg_q282_in <= (reg_q280 AND symb_decoder(16#69#)) OR
 					(reg_q280 AND symb_decoder(16#49#));
reg_q284_in <= (reg_q282 AND symb_decoder(16#53#)) OR
 					(reg_q282 AND symb_decoder(16#73#));
reg_q2387_in <= (reg_q2385 AND symb_decoder(16#72#)) OR
 					(reg_q2385 AND symb_decoder(16#52#));
reg_q2389_in <= (reg_q2387 AND symb_decoder(16#76#)) OR
 					(reg_q2387 AND symb_decoder(16#56#));
reg_q1500_in <= (reg_q1500 AND symb_decoder(16#0d#)) OR
 					(reg_q1500 AND symb_decoder(16#09#)) OR
 					(reg_q1500 AND symb_decoder(16#0a#)) OR
 					(reg_q1500 AND symb_decoder(16#20#)) OR
 					(reg_q1500 AND symb_decoder(16#0c#)) OR
 					(reg_q1498 AND symb_decoder(16#0d#)) OR
 					(reg_q1498 AND symb_decoder(16#09#)) OR
 					(reg_q1498 AND symb_decoder(16#0c#)) OR
 					(reg_q1498 AND symb_decoder(16#0a#)) OR
 					(reg_q1498 AND symb_decoder(16#20#));
reg_q2744_in <= (reg_q2742 AND symb_decoder(16#52#)) OR
 					(reg_q2742 AND symb_decoder(16#72#));
reg_q2746_in <= (reg_q2744 AND symb_decoder(16#54#)) OR
 					(reg_q2744 AND symb_decoder(16#74#));
reg_q1915_in <= (reg_q1915 AND symb_decoder(16#32#)) OR
 					(reg_q1915 AND symb_decoder(16#36#)) OR
 					(reg_q1915 AND symb_decoder(16#38#)) OR
 					(reg_q1915 AND symb_decoder(16#39#)) OR
 					(reg_q1915 AND symb_decoder(16#35#)) OR
 					(reg_q1915 AND symb_decoder(16#33#)) OR
 					(reg_q1915 AND symb_decoder(16#31#)) OR
 					(reg_q1915 AND symb_decoder(16#37#)) OR
 					(reg_q1915 AND symb_decoder(16#30#)) OR
 					(reg_q1915 AND symb_decoder(16#34#)) OR
 					(reg_q1913 AND symb_decoder(16#31#)) OR
 					(reg_q1913 AND symb_decoder(16#30#)) OR
 					(reg_q1913 AND symb_decoder(16#36#)) OR
 					(reg_q1913 AND symb_decoder(16#39#)) OR
 					(reg_q1913 AND symb_decoder(16#35#)) OR
 					(reg_q1913 AND symb_decoder(16#32#)) OR
 					(reg_q1913 AND symb_decoder(16#38#)) OR
 					(reg_q1913 AND symb_decoder(16#37#)) OR
 					(reg_q1913 AND symb_decoder(16#34#)) OR
 					(reg_q1913 AND symb_decoder(16#33#));
reg_q1498_in <= (reg_q1496 AND symb_decoder(16#68#)) OR
 					(reg_q1496 AND symb_decoder(16#48#));
reg_q218_in <= (reg_q218 AND symb_decoder(16#0c#)) OR
 					(reg_q218 AND symb_decoder(16#0d#)) OR
 					(reg_q218 AND symb_decoder(16#20#)) OR
 					(reg_q218 AND symb_decoder(16#09#)) OR
 					(reg_q218 AND symb_decoder(16#0a#)) OR
 					(reg_q216 AND symb_decoder(16#0a#)) OR
 					(reg_q216 AND symb_decoder(16#20#)) OR
 					(reg_q216 AND symb_decoder(16#09#)) OR
 					(reg_q216 AND symb_decoder(16#0d#)) OR
 					(reg_q216 AND symb_decoder(16#0c#));
reg_q220_in <= (reg_q218 AND symb_decoder(16#46#)) OR
 					(reg_q218 AND symb_decoder(16#66#));
reg_q1990_in <= (reg_q1988 AND symb_decoder(16#30#));
reg_q1992_in <= (reg_q1990 AND symb_decoder(16#30#)) OR
 					(reg_q1990 AND symb_decoder(16#61#)) OR
 					(reg_q1990 AND symb_decoder(16#65#)) OR
 					(reg_q1990 AND symb_decoder(16#64#)) OR
 					(reg_q1990 AND symb_decoder(16#34#)) OR
 					(reg_q1990 AND symb_decoder(16#44#)) OR
 					(reg_q1990 AND symb_decoder(16#45#)) OR
 					(reg_q1990 AND symb_decoder(16#43#)) OR
 					(reg_q1990 AND symb_decoder(16#46#)) OR
 					(reg_q1990 AND symb_decoder(16#36#)) OR
 					(reg_q1990 AND symb_decoder(16#66#)) OR
 					(reg_q1990 AND symb_decoder(16#63#)) OR
 					(reg_q1990 AND symb_decoder(16#35#)) OR
 					(reg_q1990 AND symb_decoder(16#37#)) OR
 					(reg_q1990 AND symb_decoder(16#39#)) OR
 					(reg_q1990 AND symb_decoder(16#42#)) OR
 					(reg_q1990 AND symb_decoder(16#41#)) OR
 					(reg_q1990 AND symb_decoder(16#32#)) OR
 					(reg_q1990 AND symb_decoder(16#33#)) OR
 					(reg_q1990 AND symb_decoder(16#31#)) OR
 					(reg_q1990 AND symb_decoder(16#38#)) OR
 					(reg_q1990 AND symb_decoder(16#62#));
reg_q2020_in <= (reg_q2018 AND symb_decoder(16#32#)) OR
 					(reg_q2018 AND symb_decoder(16#34#)) OR
 					(reg_q2018 AND symb_decoder(16#46#)) OR
 					(reg_q2018 AND symb_decoder(16#35#)) OR
 					(reg_q2018 AND symb_decoder(16#39#)) OR
 					(reg_q2018 AND symb_decoder(16#43#)) OR
 					(reg_q2018 AND symb_decoder(16#64#)) OR
 					(reg_q2018 AND symb_decoder(16#30#)) OR
 					(reg_q2018 AND symb_decoder(16#31#)) OR
 					(reg_q2018 AND symb_decoder(16#37#)) OR
 					(reg_q2018 AND symb_decoder(16#38#)) OR
 					(reg_q2018 AND symb_decoder(16#36#)) OR
 					(reg_q2018 AND symb_decoder(16#65#)) OR
 					(reg_q2018 AND symb_decoder(16#33#)) OR
 					(reg_q2018 AND symb_decoder(16#42#)) OR
 					(reg_q2018 AND symb_decoder(16#44#)) OR
 					(reg_q2018 AND symb_decoder(16#66#)) OR
 					(reg_q2018 AND symb_decoder(16#62#)) OR
 					(reg_q2018 AND symb_decoder(16#61#)) OR
 					(reg_q2018 AND symb_decoder(16#45#)) OR
 					(reg_q2018 AND symb_decoder(16#41#)) OR
 					(reg_q2018 AND symb_decoder(16#63#));
reg_q2022_in <= (reg_q2020 AND symb_decoder(16#62#)) OR
 					(reg_q2020 AND symb_decoder(16#65#)) OR
 					(reg_q2020 AND symb_decoder(16#37#)) OR
 					(reg_q2020 AND symb_decoder(16#34#)) OR
 					(reg_q2020 AND symb_decoder(16#44#)) OR
 					(reg_q2020 AND symb_decoder(16#41#)) OR
 					(reg_q2020 AND symb_decoder(16#66#)) OR
 					(reg_q2020 AND symb_decoder(16#39#)) OR
 					(reg_q2020 AND symb_decoder(16#31#)) OR
 					(reg_q2020 AND symb_decoder(16#45#)) OR
 					(reg_q2020 AND symb_decoder(16#63#)) OR
 					(reg_q2020 AND symb_decoder(16#38#)) OR
 					(reg_q2020 AND symb_decoder(16#33#)) OR
 					(reg_q2020 AND symb_decoder(16#43#)) OR
 					(reg_q2020 AND symb_decoder(16#35#)) OR
 					(reg_q2020 AND symb_decoder(16#61#)) OR
 					(reg_q2020 AND symb_decoder(16#46#)) OR
 					(reg_q2020 AND symb_decoder(16#36#)) OR
 					(reg_q2020 AND symb_decoder(16#32#)) OR
 					(reg_q2020 AND symb_decoder(16#64#)) OR
 					(reg_q2020 AND symb_decoder(16#42#)) OR
 					(reg_q2020 AND symb_decoder(16#30#));
reg_q214_in <= (reg_q214 AND symb_decoder(16#38#)) OR
 					(reg_q214 AND symb_decoder(16#33#)) OR
 					(reg_q214 AND symb_decoder(16#39#)) OR
 					(reg_q214 AND symb_decoder(16#34#)) OR
 					(reg_q214 AND symb_decoder(16#37#)) OR
 					(reg_q214 AND symb_decoder(16#30#)) OR
 					(reg_q214 AND symb_decoder(16#31#)) OR
 					(reg_q214 AND symb_decoder(16#32#)) OR
 					(reg_q214 AND symb_decoder(16#35#)) OR
 					(reg_q214 AND symb_decoder(16#36#)) OR
 					(reg_q212 AND symb_decoder(16#30#)) OR
 					(reg_q212 AND symb_decoder(16#34#)) OR
 					(reg_q212 AND symb_decoder(16#36#)) OR
 					(reg_q212 AND symb_decoder(16#38#)) OR
 					(reg_q212 AND symb_decoder(16#37#)) OR
 					(reg_q212 AND symb_decoder(16#35#)) OR
 					(reg_q212 AND symb_decoder(16#31#)) OR
 					(reg_q212 AND symb_decoder(16#39#)) OR
 					(reg_q212 AND symb_decoder(16#32#)) OR
 					(reg_q212 AND symb_decoder(16#33#));
reg_q2712_in <= (reg_q2710 AND symb_decoder(16#3a#));
reg_q2714_in <= (reg_q2712 AND symb_decoder(16#0a#)) OR
 					(reg_q2712 AND symb_decoder(16#0d#)) OR
 					(reg_q2712 AND symb_decoder(16#09#)) OR
 					(reg_q2712 AND symb_decoder(16#20#)) OR
 					(reg_q2712 AND symb_decoder(16#0c#));
reg_q2032_in <= (reg_q2030 AND symb_decoder(16#37#)) OR
 					(reg_q2030 AND symb_decoder(16#65#)) OR
 					(reg_q2030 AND symb_decoder(16#39#)) OR
 					(reg_q2030 AND symb_decoder(16#64#)) OR
 					(reg_q2030 AND symb_decoder(16#30#)) OR
 					(reg_q2030 AND symb_decoder(16#42#)) OR
 					(reg_q2030 AND symb_decoder(16#62#)) OR
 					(reg_q2030 AND symb_decoder(16#31#)) OR
 					(reg_q2030 AND symb_decoder(16#45#)) OR
 					(reg_q2030 AND symb_decoder(16#46#)) OR
 					(reg_q2030 AND symb_decoder(16#36#)) OR
 					(reg_q2030 AND symb_decoder(16#34#)) OR
 					(reg_q2030 AND symb_decoder(16#38#)) OR
 					(reg_q2030 AND symb_decoder(16#41#)) OR
 					(reg_q2030 AND symb_decoder(16#35#)) OR
 					(reg_q2030 AND symb_decoder(16#32#)) OR
 					(reg_q2030 AND symb_decoder(16#61#)) OR
 					(reg_q2030 AND symb_decoder(16#63#)) OR
 					(reg_q2030 AND symb_decoder(16#66#)) OR
 					(reg_q2030 AND symb_decoder(16#44#)) OR
 					(reg_q2030 AND symb_decoder(16#33#)) OR
 					(reg_q2030 AND symb_decoder(16#43#));
reg_q1945_in <= (reg_q1943 AND symb_decoder(16#33#));
reg_q1947_in <= (reg_q1945 AND symb_decoder(16#2a#));
reg_q124_in <= (reg_q122 AND symb_decoder(16#23#));
reg_q126_in <= (reg_q124 AND symb_decoder(16#51#)) OR
 					(reg_q124 AND symb_decoder(16#46#)) OR
 					(reg_q124 AND symb_decoder(16#56#)) OR
 					(reg_q124 AND symb_decoder(16#47#)) OR
 					(reg_q124 AND symb_decoder(16#6c#)) OR
 					(reg_q124 AND symb_decoder(16#68#)) OR
 					(reg_q124 AND symb_decoder(16#53#)) OR
 					(reg_q124 AND symb_decoder(16#79#)) OR
 					(reg_q124 AND symb_decoder(16#4d#)) OR
 					(reg_q124 AND symb_decoder(16#4f#)) OR
 					(reg_q124 AND symb_decoder(16#55#)) OR
 					(reg_q124 AND symb_decoder(16#42#)) OR
 					(reg_q124 AND symb_decoder(16#72#)) OR
 					(reg_q124 AND symb_decoder(16#4c#)) OR
 					(reg_q124 AND symb_decoder(16#52#)) OR
 					(reg_q124 AND symb_decoder(16#4e#)) OR
 					(reg_q124 AND symb_decoder(16#6d#)) OR
 					(reg_q124 AND symb_decoder(16#6e#)) OR
 					(reg_q124 AND symb_decoder(16#62#)) OR
 					(reg_q124 AND symb_decoder(16#6f#)) OR
 					(reg_q124 AND symb_decoder(16#57#)) OR
 					(reg_q124 AND symb_decoder(16#65#)) OR
 					(reg_q124 AND symb_decoder(16#54#)) OR
 					(reg_q124 AND symb_decoder(16#49#)) OR
 					(reg_q124 AND symb_decoder(16#45#)) OR
 					(reg_q124 AND symb_decoder(16#61#)) OR
 					(reg_q124 AND symb_decoder(16#78#)) OR
 					(reg_q124 AND symb_decoder(16#6a#)) OR
 					(reg_q124 AND symb_decoder(16#75#)) OR
 					(reg_q124 AND symb_decoder(16#41#)) OR
 					(reg_q124 AND symb_decoder(16#5a#)) OR
 					(reg_q124 AND symb_decoder(16#74#)) OR
 					(reg_q124 AND symb_decoder(16#43#)) OR
 					(reg_q124 AND symb_decoder(16#64#)) OR
 					(reg_q124 AND symb_decoder(16#67#)) OR
 					(reg_q124 AND symb_decoder(16#58#)) OR
 					(reg_q124 AND symb_decoder(16#59#)) OR
 					(reg_q124 AND symb_decoder(16#48#)) OR
 					(reg_q124 AND symb_decoder(16#6b#)) OR
 					(reg_q124 AND symb_decoder(16#76#)) OR
 					(reg_q124 AND symb_decoder(16#73#)) OR
 					(reg_q124 AND symb_decoder(16#7a#)) OR
 					(reg_q124 AND symb_decoder(16#4b#)) OR
 					(reg_q124 AND symb_decoder(16#50#)) OR
 					(reg_q124 AND symb_decoder(16#71#)) OR
 					(reg_q124 AND symb_decoder(16#63#)) OR
 					(reg_q124 AND symb_decoder(16#66#)) OR
 					(reg_q124 AND symb_decoder(16#77#)) OR
 					(reg_q124 AND symb_decoder(16#4a#)) OR
 					(reg_q124 AND symb_decoder(16#69#)) OR
 					(reg_q124 AND symb_decoder(16#70#)) OR
 					(reg_q124 AND symb_decoder(16#44#));
reg_q2272_in <= (reg_q2270 AND symb_decoder(16#45#)) OR
 					(reg_q2270 AND symb_decoder(16#65#));
reg_q2274_in <= (reg_q2272 AND symb_decoder(16#64#)) OR
 					(reg_q2272 AND symb_decoder(16#44#));
reg_q42_in <= (reg_q40 AND symb_decoder(16#70#)) OR
 					(reg_q40 AND symb_decoder(16#50#));
reg_q44_in <= (reg_q42 AND symb_decoder(16#61#)) OR
 					(reg_q42 AND symb_decoder(16#41#));
reg_q2028_in <= (reg_q2026 AND symb_decoder(16#44#)) OR
 					(reg_q2026 AND symb_decoder(16#30#)) OR
 					(reg_q2026 AND symb_decoder(16#61#)) OR
 					(reg_q2026 AND symb_decoder(16#35#)) OR
 					(reg_q2026 AND symb_decoder(16#66#)) OR
 					(reg_q2026 AND symb_decoder(16#36#)) OR
 					(reg_q2026 AND symb_decoder(16#42#)) OR
 					(reg_q2026 AND symb_decoder(16#31#)) OR
 					(reg_q2026 AND symb_decoder(16#41#)) OR
 					(reg_q2026 AND symb_decoder(16#63#)) OR
 					(reg_q2026 AND symb_decoder(16#37#)) OR
 					(reg_q2026 AND symb_decoder(16#64#)) OR
 					(reg_q2026 AND symb_decoder(16#62#)) OR
 					(reg_q2026 AND symb_decoder(16#46#)) OR
 					(reg_q2026 AND symb_decoder(16#34#)) OR
 					(reg_q2026 AND symb_decoder(16#43#)) OR
 					(reg_q2026 AND symb_decoder(16#45#)) OR
 					(reg_q2026 AND symb_decoder(16#39#)) OR
 					(reg_q2026 AND symb_decoder(16#38#)) OR
 					(reg_q2026 AND symb_decoder(16#65#)) OR
 					(reg_q2026 AND symb_decoder(16#33#)) OR
 					(reg_q2026 AND symb_decoder(16#32#));
reg_q2030_in <= (reg_q2028 AND symb_decoder(16#38#)) OR
 					(reg_q2028 AND symb_decoder(16#39#)) OR
 					(reg_q2028 AND symb_decoder(16#43#)) OR
 					(reg_q2028 AND symb_decoder(16#46#)) OR
 					(reg_q2028 AND symb_decoder(16#63#)) OR
 					(reg_q2028 AND symb_decoder(16#37#)) OR
 					(reg_q2028 AND symb_decoder(16#66#)) OR
 					(reg_q2028 AND symb_decoder(16#45#)) OR
 					(reg_q2028 AND symb_decoder(16#36#)) OR
 					(reg_q2028 AND symb_decoder(16#35#)) OR
 					(reg_q2028 AND symb_decoder(16#62#)) OR
 					(reg_q2028 AND symb_decoder(16#33#)) OR
 					(reg_q2028 AND symb_decoder(16#42#)) OR
 					(reg_q2028 AND symb_decoder(16#34#)) OR
 					(reg_q2028 AND symb_decoder(16#41#)) OR
 					(reg_q2028 AND symb_decoder(16#65#)) OR
 					(reg_q2028 AND symb_decoder(16#64#)) OR
 					(reg_q2028 AND symb_decoder(16#30#)) OR
 					(reg_q2028 AND symb_decoder(16#31#)) OR
 					(reg_q2028 AND symb_decoder(16#32#)) OR
 					(reg_q2028 AND symb_decoder(16#61#)) OR
 					(reg_q2028 AND symb_decoder(16#44#));
reg_q1315_in <= (reg_q1315 AND symb_decoder(16#09#)) OR
 					(reg_q1315 AND symb_decoder(16#0a#)) OR
 					(reg_q1315 AND symb_decoder(16#0c#)) OR
 					(reg_q1315 AND symb_decoder(16#20#)) OR
 					(reg_q1315 AND symb_decoder(16#0d#)) OR
 					(reg_q1313 AND symb_decoder(16#0d#)) OR
 					(reg_q1313 AND symb_decoder(16#0a#)) OR
 					(reg_q1313 AND symb_decoder(16#20#)) OR
 					(reg_q1313 AND symb_decoder(16#09#)) OR
 					(reg_q1313 AND symb_decoder(16#0c#));
reg_q2704_in <= (reg_q2702 AND symb_decoder(16#76#)) OR
 					(reg_q2702 AND symb_decoder(16#56#));
reg_q2706_in <= (reg_q2704 AND symb_decoder(16#65#)) OR
 					(reg_q2704 AND symb_decoder(16#45#));
reg_q1994_in <= (reg_q1992 AND symb_decoder(16#31#)) OR
 					(reg_q1992 AND symb_decoder(16#38#)) OR
 					(reg_q1992 AND symb_decoder(16#64#)) OR
 					(reg_q1992 AND symb_decoder(16#42#)) OR
 					(reg_q1992 AND symb_decoder(16#37#)) OR
 					(reg_q1992 AND symb_decoder(16#30#)) OR
 					(reg_q1992 AND symb_decoder(16#33#)) OR
 					(reg_q1992 AND symb_decoder(16#65#)) OR
 					(reg_q1992 AND symb_decoder(16#39#)) OR
 					(reg_q1992 AND symb_decoder(16#34#)) OR
 					(reg_q1992 AND symb_decoder(16#66#)) OR
 					(reg_q1992 AND symb_decoder(16#46#)) OR
 					(reg_q1992 AND symb_decoder(16#36#)) OR
 					(reg_q1992 AND symb_decoder(16#45#)) OR
 					(reg_q1992 AND symb_decoder(16#44#)) OR
 					(reg_q1992 AND symb_decoder(16#32#)) OR
 					(reg_q1992 AND symb_decoder(16#61#)) OR
 					(reg_q1992 AND symb_decoder(16#41#)) OR
 					(reg_q1992 AND symb_decoder(16#43#)) OR
 					(reg_q1992 AND symb_decoder(16#62#)) OR
 					(reg_q1992 AND symb_decoder(16#35#)) OR
 					(reg_q1992 AND symb_decoder(16#63#));
reg_q1804_in <= (reg_q1802 AND symb_decoder(16#76#)) OR
 					(reg_q1802 AND symb_decoder(16#56#));
reg_q1806_in <= (reg_q1804 AND symb_decoder(16#32#)) OR
 					(reg_q1804 AND symb_decoder(16#34#)) OR
 					(reg_q1804 AND symb_decoder(16#37#)) OR
 					(reg_q1804 AND symb_decoder(16#31#)) OR
 					(reg_q1804 AND symb_decoder(16#39#)) OR
 					(reg_q1804 AND symb_decoder(16#35#)) OR
 					(reg_q1804 AND symb_decoder(16#36#)) OR
 					(reg_q1804 AND symb_decoder(16#30#)) OR
 					(reg_q1804 AND symb_decoder(16#33#)) OR
 					(reg_q1804 AND symb_decoder(16#38#)) OR
 					(reg_q1806 AND symb_decoder(16#36#)) OR
 					(reg_q1806 AND symb_decoder(16#38#)) OR
 					(reg_q1806 AND symb_decoder(16#34#)) OR
 					(reg_q1806 AND symb_decoder(16#39#)) OR
 					(reg_q1806 AND symb_decoder(16#37#)) OR
 					(reg_q1806 AND symb_decoder(16#35#)) OR
 					(reg_q1806 AND symb_decoder(16#30#)) OR
 					(reg_q1806 AND symb_decoder(16#31#)) OR
 					(reg_q1806 AND symb_decoder(16#33#)) OR
 					(reg_q1806 AND symb_decoder(16#32#));
reg_q698_in <= (reg_q696 AND symb_decoder(16#54#)) OR
 					(reg_q696 AND symb_decoder(16#74#));
reg_q700_in <= (reg_q698 AND symb_decoder(16#61#)) OR
 					(reg_q698 AND symb_decoder(16#41#));
reg_q2617_in <= (reg_q2617 AND symb_decoder(16#20#)) OR
 					(reg_q2617 AND symb_decoder(16#0d#)) OR
 					(reg_q2617 AND symb_decoder(16#09#)) OR
 					(reg_q2617 AND symb_decoder(16#0a#)) OR
 					(reg_q2617 AND symb_decoder(16#0c#)) OR
 					(reg_q2615 AND symb_decoder(16#0d#)) OR
 					(reg_q2615 AND symb_decoder(16#20#)) OR
 					(reg_q2615 AND symb_decoder(16#0c#)) OR
 					(reg_q2615 AND symb_decoder(16#09#)) OR
 					(reg_q2615 AND symb_decoder(16#0a#));
reg_q768_in <= (reg_q767 AND symb_decoder(16#0d#));
reg_q2752_in <= (reg_q2750 AND symb_decoder(16#5c#));
reg_q2754_in <= (reg_q2752 AND symb_decoder(16#21#));
reg_q1701_in <= (reg_q1699 AND symb_decoder(16#58#)) OR
 					(reg_q1699 AND symb_decoder(16#78#));
reg_q1703_in <= (reg_q1701 AND symb_decoder(16#20#)) OR
 					(reg_q1701 AND symb_decoder(16#09#)) OR
 					(reg_q1701 AND symb_decoder(16#0a#)) OR
 					(reg_q1701 AND symb_decoder(16#0d#)) OR
 					(reg_q1701 AND symb_decoder(16#0c#)) OR
 					(reg_q1703 AND symb_decoder(16#20#)) OR
 					(reg_q1703 AND symb_decoder(16#09#)) OR
 					(reg_q1703 AND symb_decoder(16#0d#)) OR
 					(reg_q1703 AND symb_decoder(16#0c#)) OR
 					(reg_q1703 AND symb_decoder(16#0a#));
reg_q120_in <= (reg_q118 AND symb_decoder(16#65#)) OR
 					(reg_q118 AND symb_decoder(16#45#));
reg_q122_in <= (reg_q120 AND symb_decoder(16#51#)) OR
 					(reg_q120 AND symb_decoder(16#71#));
reg_q2726_in <= (reg_q2724 AND symb_decoder(16#47#)) OR
 					(reg_q2724 AND symb_decoder(16#67#));
reg_q2728_in <= (reg_q2726 AND symb_decoder(16#47#)) OR
 					(reg_q2726 AND symb_decoder(16#67#));
reg_q2040_in <= (reg_q2038 AND symb_decoder(16#41#)) OR
 					(reg_q2038 AND symb_decoder(16#32#)) OR
 					(reg_q2038 AND symb_decoder(16#44#)) OR
 					(reg_q2038 AND symb_decoder(16#42#)) OR
 					(reg_q2038 AND symb_decoder(16#66#)) OR
 					(reg_q2038 AND symb_decoder(16#65#)) OR
 					(reg_q2038 AND symb_decoder(16#34#)) OR
 					(reg_q2038 AND symb_decoder(16#33#)) OR
 					(reg_q2038 AND symb_decoder(16#36#)) OR
 					(reg_q2038 AND symb_decoder(16#35#)) OR
 					(reg_q2038 AND symb_decoder(16#30#)) OR
 					(reg_q2038 AND symb_decoder(16#37#)) OR
 					(reg_q2038 AND symb_decoder(16#45#)) OR
 					(reg_q2038 AND symb_decoder(16#61#)) OR
 					(reg_q2038 AND symb_decoder(16#39#)) OR
 					(reg_q2038 AND symb_decoder(16#62#)) OR
 					(reg_q2038 AND symb_decoder(16#64#)) OR
 					(reg_q2038 AND symb_decoder(16#63#)) OR
 					(reg_q2038 AND symb_decoder(16#43#)) OR
 					(reg_q2038 AND symb_decoder(16#31#)) OR
 					(reg_q2038 AND symb_decoder(16#38#)) OR
 					(reg_q2038 AND symb_decoder(16#46#));
reg_q2042_in <= (reg_q2040 AND symb_decoder(16#45#)) OR
 					(reg_q2040 AND symb_decoder(16#61#)) OR
 					(reg_q2040 AND symb_decoder(16#38#)) OR
 					(reg_q2040 AND symb_decoder(16#35#)) OR
 					(reg_q2040 AND symb_decoder(16#36#)) OR
 					(reg_q2040 AND symb_decoder(16#32#)) OR
 					(reg_q2040 AND symb_decoder(16#44#)) OR
 					(reg_q2040 AND symb_decoder(16#43#)) OR
 					(reg_q2040 AND symb_decoder(16#34#)) OR
 					(reg_q2040 AND symb_decoder(16#65#)) OR
 					(reg_q2040 AND symb_decoder(16#37#)) OR
 					(reg_q2040 AND symb_decoder(16#33#)) OR
 					(reg_q2040 AND symb_decoder(16#62#)) OR
 					(reg_q2040 AND symb_decoder(16#66#)) OR
 					(reg_q2040 AND symb_decoder(16#30#)) OR
 					(reg_q2040 AND symb_decoder(16#63#)) OR
 					(reg_q2040 AND symb_decoder(16#42#)) OR
 					(reg_q2040 AND symb_decoder(16#41#)) OR
 					(reg_q2040 AND symb_decoder(16#46#)) OR
 					(reg_q2040 AND symb_decoder(16#39#)) OR
 					(reg_q2040 AND symb_decoder(16#31#)) OR
 					(reg_q2040 AND symb_decoder(16#64#));
reg_q208_in <= (reg_q206 AND symb_decoder(16#2e#));
reg_q1126_in <= (reg_q1126 AND symb_decoder(16#20#)) OR
 					(reg_q1126 AND symb_decoder(16#0d#)) OR
 					(reg_q1126 AND symb_decoder(16#0a#)) OR
 					(reg_q1126 AND symb_decoder(16#09#)) OR
 					(reg_q1126 AND symb_decoder(16#0c#)) OR
 					(reg_q1124 AND symb_decoder(16#0a#)) OR
 					(reg_q1124 AND symb_decoder(16#09#)) OR
 					(reg_q1124 AND symb_decoder(16#0c#)) OR
 					(reg_q1124 AND symb_decoder(16#0d#)) OR
 					(reg_q1124 AND symb_decoder(16#20#));
reg_q1212_in <= (reg_q1210 AND symb_decoder(16#2e#));
reg_q1214_in <= (reg_q1212 AND symb_decoder(16#38#)) OR
 					(reg_q1212 AND symb_decoder(16#31#)) OR
 					(reg_q1212 AND symb_decoder(16#37#)) OR
 					(reg_q1212 AND symb_decoder(16#39#)) OR
 					(reg_q1212 AND symb_decoder(16#30#)) OR
 					(reg_q1212 AND symb_decoder(16#34#)) OR
 					(reg_q1212 AND symb_decoder(16#32#)) OR
 					(reg_q1212 AND symb_decoder(16#36#)) OR
 					(reg_q1212 AND symb_decoder(16#33#)) OR
 					(reg_q1212 AND symb_decoder(16#35#)) OR
 					(reg_q1214 AND symb_decoder(16#32#)) OR
 					(reg_q1214 AND symb_decoder(16#30#)) OR
 					(reg_q1214 AND symb_decoder(16#37#)) OR
 					(reg_q1214 AND symb_decoder(16#33#)) OR
 					(reg_q1214 AND symb_decoder(16#36#)) OR
 					(reg_q1214 AND symb_decoder(16#31#)) OR
 					(reg_q1214 AND symb_decoder(16#39#)) OR
 					(reg_q1214 AND symb_decoder(16#38#)) OR
 					(reg_q1214 AND symb_decoder(16#35#)) OR
 					(reg_q1214 AND symb_decoder(16#34#));
reg_q2316_in <= (reg_q2314 AND symb_decoder(16#73#)) OR
 					(reg_q2314 AND symb_decoder(16#53#));
reg_q2018_in <= (reg_q2016 AND symb_decoder(16#62#)) OR
 					(reg_q2016 AND symb_decoder(16#66#)) OR
 					(reg_q2016 AND symb_decoder(16#63#)) OR
 					(reg_q2016 AND symb_decoder(16#44#)) OR
 					(reg_q2016 AND symb_decoder(16#41#)) OR
 					(reg_q2016 AND symb_decoder(16#32#)) OR
 					(reg_q2016 AND symb_decoder(16#43#)) OR
 					(reg_q2016 AND symb_decoder(16#33#)) OR
 					(reg_q2016 AND symb_decoder(16#36#)) OR
 					(reg_q2016 AND symb_decoder(16#64#)) OR
 					(reg_q2016 AND symb_decoder(16#39#)) OR
 					(reg_q2016 AND symb_decoder(16#35#)) OR
 					(reg_q2016 AND symb_decoder(16#61#)) OR
 					(reg_q2016 AND symb_decoder(16#45#)) OR
 					(reg_q2016 AND symb_decoder(16#42#)) OR
 					(reg_q2016 AND symb_decoder(16#38#)) OR
 					(reg_q2016 AND symb_decoder(16#30#)) OR
 					(reg_q2016 AND symb_decoder(16#37#)) OR
 					(reg_q2016 AND symb_decoder(16#31#)) OR
 					(reg_q2016 AND symb_decoder(16#46#)) OR
 					(reg_q2016 AND symb_decoder(16#65#)) OR
 					(reg_q2016 AND symb_decoder(16#34#));
reg_q355_in <= (reg_q353 AND symb_decoder(16#45#)) OR
 					(reg_q353 AND symb_decoder(16#65#));
reg_q357_in <= (reg_q355 AND symb_decoder(16#72#)) OR
 					(reg_q355 AND symb_decoder(16#52#));
reg_q776_in <= (reg_q774 AND symb_decoder(16#75#)) OR
 					(reg_q774 AND symb_decoder(16#55#));
reg_q778_in <= (reg_q776 AND symb_decoder(16#62#)) OR
 					(reg_q776 AND symb_decoder(16#42#));
reg_q58_in <= (reg_q56 AND symb_decoder(16#0d#));
reg_q60_in <= (reg_q58 AND symb_decoder(16#0a#));
reg_q1183_in <= (reg_q1183 AND symb_decoder(16#37#)) OR
 					(reg_q1183 AND symb_decoder(16#32#)) OR
 					(reg_q1183 AND symb_decoder(16#39#)) OR
 					(reg_q1183 AND symb_decoder(16#35#)) OR
 					(reg_q1183 AND symb_decoder(16#33#)) OR
 					(reg_q1183 AND symb_decoder(16#38#)) OR
 					(reg_q1183 AND symb_decoder(16#34#)) OR
 					(reg_q1183 AND symb_decoder(16#30#)) OR
 					(reg_q1183 AND symb_decoder(16#36#)) OR
 					(reg_q1183 AND symb_decoder(16#31#)) OR
 					(reg_q1181 AND symb_decoder(16#39#)) OR
 					(reg_q1181 AND symb_decoder(16#36#)) OR
 					(reg_q1181 AND symb_decoder(16#31#)) OR
 					(reg_q1181 AND symb_decoder(16#32#)) OR
 					(reg_q1181 AND symb_decoder(16#34#)) OR
 					(reg_q1181 AND symb_decoder(16#37#)) OR
 					(reg_q1181 AND symb_decoder(16#30#)) OR
 					(reg_q1181 AND symb_decoder(16#33#)) OR
 					(reg_q1181 AND symb_decoder(16#38#)) OR
 					(reg_q1181 AND symb_decoder(16#35#));
reg_q718_in <= (reg_q718 AND symb_decoder(16#0d#)) OR
 					(reg_q718 AND symb_decoder(16#0a#)) OR
 					(reg_q718 AND symb_decoder(16#20#)) OR
 					(reg_q718 AND symb_decoder(16#0c#)) OR
 					(reg_q718 AND symb_decoder(16#09#)) OR
 					(reg_q716 AND symb_decoder(16#0c#)) OR
 					(reg_q716 AND symb_decoder(16#20#)) OR
 					(reg_q716 AND symb_decoder(16#0d#)) OR
 					(reg_q716 AND symb_decoder(16#0a#)) OR
 					(reg_q716 AND symb_decoder(16#09#));
reg_q972_in <= (reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q971 AND symb_decoder(16#74#)) OR
 					(reg_q971 AND symb_decoder(16#54#));
reg_q974_in <= (reg_q972 AND symb_decoder(16#46#)) OR
 					(reg_q972 AND symb_decoder(16#66#));
reg_q2012_in <= (reg_q2010 AND symb_decoder(16#45#)) OR
 					(reg_q2010 AND symb_decoder(16#64#)) OR
 					(reg_q2010 AND symb_decoder(16#41#)) OR
 					(reg_q2010 AND symb_decoder(16#46#)) OR
 					(reg_q2010 AND symb_decoder(16#35#)) OR
 					(reg_q2010 AND symb_decoder(16#43#)) OR
 					(reg_q2010 AND symb_decoder(16#31#)) OR
 					(reg_q2010 AND symb_decoder(16#63#)) OR
 					(reg_q2010 AND symb_decoder(16#62#)) OR
 					(reg_q2010 AND symb_decoder(16#30#)) OR
 					(reg_q2010 AND symb_decoder(16#37#)) OR
 					(reg_q2010 AND symb_decoder(16#33#)) OR
 					(reg_q2010 AND symb_decoder(16#32#)) OR
 					(reg_q2010 AND symb_decoder(16#38#)) OR
 					(reg_q2010 AND symb_decoder(16#44#)) OR
 					(reg_q2010 AND symb_decoder(16#66#)) OR
 					(reg_q2010 AND symb_decoder(16#36#)) OR
 					(reg_q2010 AND symb_decoder(16#42#)) OR
 					(reg_q2010 AND symb_decoder(16#61#)) OR
 					(reg_q2010 AND symb_decoder(16#65#)) OR
 					(reg_q2010 AND symb_decoder(16#34#)) OR
 					(reg_q2010 AND symb_decoder(16#39#));
reg_q2014_in <= (reg_q2012 AND symb_decoder(16#63#)) OR
 					(reg_q2012 AND symb_decoder(16#42#)) OR
 					(reg_q2012 AND symb_decoder(16#41#)) OR
 					(reg_q2012 AND symb_decoder(16#38#)) OR
 					(reg_q2012 AND symb_decoder(16#30#)) OR
 					(reg_q2012 AND symb_decoder(16#64#)) OR
 					(reg_q2012 AND symb_decoder(16#61#)) OR
 					(reg_q2012 AND symb_decoder(16#62#)) OR
 					(reg_q2012 AND symb_decoder(16#33#)) OR
 					(reg_q2012 AND symb_decoder(16#35#)) OR
 					(reg_q2012 AND symb_decoder(16#37#)) OR
 					(reg_q2012 AND symb_decoder(16#31#)) OR
 					(reg_q2012 AND symb_decoder(16#34#)) OR
 					(reg_q2012 AND symb_decoder(16#65#)) OR
 					(reg_q2012 AND symb_decoder(16#45#)) OR
 					(reg_q2012 AND symb_decoder(16#43#)) OR
 					(reg_q2012 AND symb_decoder(16#66#)) OR
 					(reg_q2012 AND symb_decoder(16#36#)) OR
 					(reg_q2012 AND symb_decoder(16#44#)) OR
 					(reg_q2012 AND symb_decoder(16#46#)) OR
 					(reg_q2012 AND symb_decoder(16#39#)) OR
 					(reg_q2012 AND symb_decoder(16#32#));
reg_q2383_in <= (reg_q2409 AND symb_decoder(16#73#)) OR
 					(reg_q2409 AND symb_decoder(16#53#)) OR
 					(reg_q2415 AND symb_decoder(16#73#)) OR
 					(reg_q2415 AND symb_decoder(16#53#)) OR
 					(reg_q2379 AND symb_decoder(16#53#)) OR
 					(reg_q2379 AND symb_decoder(16#73#));
reg_q2385_in <= (reg_q2383 AND symb_decoder(16#65#)) OR
 					(reg_q2383 AND symb_decoder(16#45#));
reg_q782_in <= (reg_q780 AND symb_decoder(16#45#)) OR
 					(reg_q780 AND symb_decoder(16#65#));
reg_q784_in <= (reg_q782 AND symb_decoder(16#43#)) OR
 					(reg_q782 AND symb_decoder(16#63#));
reg_q501_in <= (reg_q499 AND symb_decoder(16#49#)) OR
 					(reg_q499 AND symb_decoder(16#69#));
reg_q1707_in <= (reg_q1705 AND symb_decoder(16#52#)) OR
 					(reg_q1705 AND symb_decoder(16#72#));
reg_q1949_in <= (reg_q1947 AND symb_decoder(16#33#)) OR
 					(reg_q1947 AND symb_decoder(16#37#)) OR
 					(reg_q1947 AND symb_decoder(16#34#)) OR
 					(reg_q1947 AND symb_decoder(16#39#)) OR
 					(reg_q1947 AND symb_decoder(16#35#)) OR
 					(reg_q1947 AND symb_decoder(16#30#)) OR
 					(reg_q1947 AND symb_decoder(16#31#)) OR
 					(reg_q1947 AND symb_decoder(16#38#)) OR
 					(reg_q1947 AND symb_decoder(16#36#)) OR
 					(reg_q1947 AND symb_decoder(16#32#)) OR
 					(reg_q1949 AND symb_decoder(16#38#)) OR
 					(reg_q1949 AND symb_decoder(16#37#)) OR
 					(reg_q1949 AND symb_decoder(16#30#)) OR
 					(reg_q1949 AND symb_decoder(16#36#)) OR
 					(reg_q1949 AND symb_decoder(16#32#)) OR
 					(reg_q1949 AND symb_decoder(16#39#)) OR
 					(reg_q1949 AND symb_decoder(16#34#)) OR
 					(reg_q1949 AND symb_decoder(16#35#)) OR
 					(reg_q1949 AND symb_decoder(16#33#)) OR
 					(reg_q1949 AND symb_decoder(16#31#));
reg_q52_in <= (reg_q50 AND symb_decoder(16#6f#)) OR
 					(reg_q50 AND symb_decoder(16#4f#));
reg_q54_in <= (reg_q52 AND symb_decoder(16#72#)) OR
 					(reg_q52 AND symb_decoder(16#52#));
reg_q2621_in <= (reg_q2619 AND symb_decoder(16#2e#));
reg_q238_in <= (reg_q236 AND symb_decoder(16#47#)) OR
 					(reg_q236 AND symb_decoder(16#67#));
reg_q240_in <= (reg_q238 AND symb_decoder(16#75#)) OR
 					(reg_q238 AND symb_decoder(16#55#));
reg_q716_in <= (reg_q714 AND symb_decoder(16#53#)) OR
 					(reg_q714 AND symb_decoder(16#73#));
reg_q1187_in <= (reg_q1187 AND symb_decoder(16#38#)) OR
 					(reg_q1187 AND symb_decoder(16#36#)) OR
 					(reg_q1187 AND symb_decoder(16#31#)) OR
 					(reg_q1187 AND symb_decoder(16#30#)) OR
 					(reg_q1187 AND symb_decoder(16#37#)) OR
 					(reg_q1187 AND symb_decoder(16#33#)) OR
 					(reg_q1187 AND symb_decoder(16#32#)) OR
 					(reg_q1187 AND symb_decoder(16#35#)) OR
 					(reg_q1187 AND symb_decoder(16#34#)) OR
 					(reg_q1187 AND symb_decoder(16#39#)) OR
 					(reg_q1185 AND symb_decoder(16#32#)) OR
 					(reg_q1185 AND symb_decoder(16#31#)) OR
 					(reg_q1185 AND symb_decoder(16#35#)) OR
 					(reg_q1185 AND symb_decoder(16#39#)) OR
 					(reg_q1185 AND symb_decoder(16#38#)) OR
 					(reg_q1185 AND symb_decoder(16#33#)) OR
 					(reg_q1185 AND symb_decoder(16#34#)) OR
 					(reg_q1185 AND symb_decoder(16#36#)) OR
 					(reg_q1185 AND symb_decoder(16#37#)) OR
 					(reg_q1185 AND symb_decoder(16#30#));
reg_q1189_in <= (reg_q1187 AND symb_decoder(16#0d#)) OR
 					(reg_q1187 AND symb_decoder(16#0c#)) OR
 					(reg_q1187 AND symb_decoder(16#09#)) OR
 					(reg_q1187 AND symb_decoder(16#20#)) OR
 					(reg_q1187 AND symb_decoder(16#0a#)) OR
 					(reg_q1189 AND symb_decoder(16#20#)) OR
 					(reg_q1189 AND symb_decoder(16#0c#)) OR
 					(reg_q1189 AND symb_decoder(16#0d#)) OR
 					(reg_q1189 AND symb_decoder(16#0a#)) OR
 					(reg_q1189 AND symb_decoder(16#09#));
reg_q2597_in <= (reg_q2595 AND symb_decoder(16#43#)) OR
 					(reg_q2595 AND symb_decoder(16#63#));
reg_q2599_in <= (reg_q2597 AND symb_decoder(16#74#)) OR
 					(reg_q2597 AND symb_decoder(16#54#));
reg_q141_in <= (reg_q139 AND symb_decoder(16#45#)) OR
 					(reg_q139 AND symb_decoder(16#65#));
reg_q143_in <= (reg_q141 AND symb_decoder(16#52#)) OR
 					(reg_q141 AND symb_decoder(16#72#));
reg_q1768_in <= (reg_q1766 AND symb_decoder(16#66#)) OR
 					(reg_q1766 AND symb_decoder(16#46#));
reg_q1770_in <= (reg_q1768 AND symb_decoder(16#0c#)) OR
 					(reg_q1768 AND symb_decoder(16#09#)) OR
 					(reg_q1768 AND symb_decoder(16#0a#)) OR
 					(reg_q1768 AND symb_decoder(16#20#)) OR
 					(reg_q1768 AND symb_decoder(16#0d#)) OR
 					(reg_q1770 AND symb_decoder(16#0a#)) OR
 					(reg_q1770 AND symb_decoder(16#20#)) OR
 					(reg_q1770 AND symb_decoder(16#09#)) OR
 					(reg_q1770 AND symb_decoder(16#0c#)) OR
 					(reg_q1770 AND symb_decoder(16#0d#));
reg_q2288_in <= (reg_q2286 AND symb_decoder(16#3a#));
reg_q2000_in <= (reg_q1998 AND symb_decoder(16#41#)) OR
 					(reg_q1998 AND symb_decoder(16#62#)) OR
 					(reg_q1998 AND symb_decoder(16#63#)) OR
 					(reg_q1998 AND symb_decoder(16#61#)) OR
 					(reg_q1998 AND symb_decoder(16#66#)) OR
 					(reg_q1998 AND symb_decoder(16#33#)) OR
 					(reg_q1998 AND symb_decoder(16#65#)) OR
 					(reg_q1998 AND symb_decoder(16#42#)) OR
 					(reg_q1998 AND symb_decoder(16#38#)) OR
 					(reg_q1998 AND symb_decoder(16#32#)) OR
 					(reg_q1998 AND symb_decoder(16#64#)) OR
 					(reg_q1998 AND symb_decoder(16#34#)) OR
 					(reg_q1998 AND symb_decoder(16#46#)) OR
 					(reg_q1998 AND symb_decoder(16#30#)) OR
 					(reg_q1998 AND symb_decoder(16#39#)) OR
 					(reg_q1998 AND symb_decoder(16#43#)) OR
 					(reg_q1998 AND symb_decoder(16#36#)) OR
 					(reg_q1998 AND symb_decoder(16#44#)) OR
 					(reg_q1998 AND symb_decoder(16#45#)) OR
 					(reg_q1998 AND symb_decoder(16#35#)) OR
 					(reg_q1998 AND symb_decoder(16#31#)) OR
 					(reg_q1998 AND symb_decoder(16#37#));
reg_q1717_in <= (reg_q1715 AND symb_decoder(16#2e#));
reg_q2225_in <= (reg_q2223 AND symb_decoder(16#6c#)) OR
 					(reg_q2223 AND symb_decoder(16#67#)) OR
 					(reg_q2223 AND symb_decoder(16#4c#)) OR
 					(reg_q2223 AND symb_decoder(16#47#));
reg_q2227_in <= (reg_q2225 AND symb_decoder(16#72#)) OR
 					(reg_q2225 AND symb_decoder(16#52#));
reg_q50_in <= (reg_q48 AND symb_decoder(16#77#)) OR
 					(reg_q48 AND symb_decoder(16#57#));
reg_q557_in <= (reg_q555 AND symb_decoder(16#72#)) OR
 					(reg_q555 AND symb_decoder(16#52#));
reg_q559_in <= (reg_q557 AND symb_decoder(16#56#)) OR
 					(reg_q557 AND symb_decoder(16#76#));
reg_q478_in <= (reg_q478 AND symb_decoder(16#35#)) OR
 					(reg_q478 AND symb_decoder(16#33#)) OR
 					(reg_q478 AND symb_decoder(16#39#)) OR
 					(reg_q478 AND symb_decoder(16#32#)) OR
 					(reg_q478 AND symb_decoder(16#31#)) OR
 					(reg_q478 AND symb_decoder(16#34#)) OR
 					(reg_q478 AND symb_decoder(16#37#)) OR
 					(reg_q478 AND symb_decoder(16#38#)) OR
 					(reg_q478 AND symb_decoder(16#30#)) OR
 					(reg_q478 AND symb_decoder(16#36#)) OR
 					(reg_q476 AND symb_decoder(16#31#)) OR
 					(reg_q476 AND symb_decoder(16#35#)) OR
 					(reg_q476 AND symb_decoder(16#37#)) OR
 					(reg_q476 AND symb_decoder(16#34#)) OR
 					(reg_q476 AND symb_decoder(16#30#)) OR
 					(reg_q476 AND symb_decoder(16#39#)) OR
 					(reg_q476 AND symb_decoder(16#33#)) OR
 					(reg_q476 AND symb_decoder(16#32#)) OR
 					(reg_q476 AND symb_decoder(16#36#)) OR
 					(reg_q476 AND symb_decoder(16#38#));
reg_q2619_in <= (reg_q2617 AND symb_decoder(16#37#)) OR
 					(reg_q2617 AND symb_decoder(16#38#)) OR
 					(reg_q2617 AND symb_decoder(16#30#)) OR
 					(reg_q2617 AND symb_decoder(16#39#)) OR
 					(reg_q2617 AND symb_decoder(16#36#)) OR
 					(reg_q2617 AND symb_decoder(16#35#)) OR
 					(reg_q2617 AND symb_decoder(16#33#)) OR
 					(reg_q2617 AND symb_decoder(16#32#)) OR
 					(reg_q2617 AND symb_decoder(16#31#)) OR
 					(reg_q2617 AND symb_decoder(16#34#)) OR
 					(reg_q2619 AND symb_decoder(16#35#)) OR
 					(reg_q2619 AND symb_decoder(16#30#)) OR
 					(reg_q2619 AND symb_decoder(16#31#)) OR
 					(reg_q2619 AND symb_decoder(16#37#)) OR
 					(reg_q2619 AND symb_decoder(16#39#)) OR
 					(reg_q2619 AND symb_decoder(16#32#)) OR
 					(reg_q2619 AND symb_decoder(16#33#)) OR
 					(reg_q2619 AND symb_decoder(16#36#)) OR
 					(reg_q2619 AND symb_decoder(16#34#)) OR
 					(reg_q2619 AND symb_decoder(16#38#));
reg_q2004_in <= (reg_q2002 AND symb_decoder(16#41#)) OR
 					(reg_q2002 AND symb_decoder(16#32#)) OR
 					(reg_q2002 AND symb_decoder(16#61#)) OR
 					(reg_q2002 AND symb_decoder(16#63#)) OR
 					(reg_q2002 AND symb_decoder(16#66#)) OR
 					(reg_q2002 AND symb_decoder(16#42#)) OR
 					(reg_q2002 AND symb_decoder(16#30#)) OR
 					(reg_q2002 AND symb_decoder(16#39#)) OR
 					(reg_q2002 AND symb_decoder(16#64#)) OR
 					(reg_q2002 AND symb_decoder(16#62#)) OR
 					(reg_q2002 AND symb_decoder(16#35#)) OR
 					(reg_q2002 AND symb_decoder(16#44#)) OR
 					(reg_q2002 AND symb_decoder(16#45#)) OR
 					(reg_q2002 AND symb_decoder(16#37#)) OR
 					(reg_q2002 AND symb_decoder(16#34#)) OR
 					(reg_q2002 AND symb_decoder(16#33#)) OR
 					(reg_q2002 AND symb_decoder(16#43#)) OR
 					(reg_q2002 AND symb_decoder(16#65#)) OR
 					(reg_q2002 AND symb_decoder(16#31#)) OR
 					(reg_q2002 AND symb_decoder(16#38#)) OR
 					(reg_q2002 AND symb_decoder(16#36#)) OR
 					(reg_q2002 AND symb_decoder(16#46#));
reg_q212_in <= (reg_q210 AND symb_decoder(16#2e#));
reg_q2276_in <= (reg_q2274 AND symb_decoder(16#20#)) OR
 					(reg_q2274 AND symb_decoder(16#0a#)) OR
 					(reg_q2274 AND symb_decoder(16#09#)) OR
 					(reg_q2274 AND symb_decoder(16#0c#)) OR
 					(reg_q2274 AND symb_decoder(16#0d#)) OR
 					(reg_q2276 AND symb_decoder(16#0a#)) OR
 					(reg_q2276 AND symb_decoder(16#09#)) OR
 					(reg_q2276 AND symb_decoder(16#0c#)) OR
 					(reg_q2276 AND symb_decoder(16#20#)) OR
 					(reg_q2276 AND symb_decoder(16#0d#));
reg_q2278_in <= (reg_q2276 AND symb_decoder(16#6f#)) OR
 					(reg_q2276 AND symb_decoder(16#4f#));
reg_q1778_in <= (reg_q1776 AND symb_decoder(16#6f#)) OR
 					(reg_q1776 AND symb_decoder(16#4f#));
reg_q1780_in <= (reg_q1778 AND symb_decoder(16#74#)) OR
 					(reg_q1778 AND symb_decoder(16#54#));
reg_q2264_in <= (reg_q2262 AND symb_decoder(16#53#)) OR
 					(reg_q2262 AND symb_decoder(16#73#));
reg_q2266_in <= (reg_q2264 AND symb_decoder(16#74#)) OR
 					(reg_q2264 AND symb_decoder(16#54#));
reg_q1136_in <= (reg_q1136 AND symb_decoder(16#20#)) OR
 					(reg_q1136 AND symb_decoder(16#0d#)) OR
 					(reg_q1136 AND symb_decoder(16#09#)) OR
 					(reg_q1136 AND symb_decoder(16#0c#)) OR
 					(reg_q1136 AND symb_decoder(16#0a#)) OR
 					(reg_q1134 AND symb_decoder(16#0c#)) OR
 					(reg_q1134 AND symb_decoder(16#0a#)) OR
 					(reg_q1134 AND symb_decoder(16#0d#)) OR
 					(reg_q1134 AND symb_decoder(16#20#)) OR
 					(reg_q1134 AND symb_decoder(16#09#));
reg_q69_in <= (reg_q67 AND symb_decoder(16#2d#));
reg_q71_in <= (reg_q69 AND symb_decoder(16#0d#)) OR
 					(reg_q69 AND symb_decoder(16#0a#)) OR
 					(reg_q69 AND symb_decoder(16#2a#));
reg_q171_in <= (reg_q169 AND symb_decoder(16#2e#));
reg_q1721_in <= (reg_q1719 AND symb_decoder(16#0a#)) OR
 					(reg_q1719 AND symb_decoder(16#20#)) OR
 					(reg_q1719 AND symb_decoder(16#0c#)) OR
 					(reg_q1719 AND symb_decoder(16#09#)) OR
 					(reg_q1719 AND symb_decoder(16#0d#)) OR
 					(reg_q1721 AND symb_decoder(16#09#)) OR
 					(reg_q1721 AND symb_decoder(16#0a#)) OR
 					(reg_q1721 AND symb_decoder(16#20#)) OR
 					(reg_q1721 AND symb_decoder(16#0d#)) OR
 					(reg_q1721 AND symb_decoder(16#0c#));
reg_q2016_in <= (reg_q2014 AND symb_decoder(16#33#)) OR
 					(reg_q2014 AND symb_decoder(16#44#)) OR
 					(reg_q2014 AND symb_decoder(16#46#)) OR
 					(reg_q2014 AND symb_decoder(16#62#)) OR
 					(reg_q2014 AND symb_decoder(16#35#)) OR
 					(reg_q2014 AND symb_decoder(16#61#)) OR
 					(reg_q2014 AND symb_decoder(16#32#)) OR
 					(reg_q2014 AND symb_decoder(16#64#)) OR
 					(reg_q2014 AND symb_decoder(16#34#)) OR
 					(reg_q2014 AND symb_decoder(16#43#)) OR
 					(reg_q2014 AND symb_decoder(16#37#)) OR
 					(reg_q2014 AND symb_decoder(16#38#)) OR
 					(reg_q2014 AND symb_decoder(16#66#)) OR
 					(reg_q2014 AND symb_decoder(16#63#)) OR
 					(reg_q2014 AND symb_decoder(16#31#)) OR
 					(reg_q2014 AND symb_decoder(16#39#)) OR
 					(reg_q2014 AND symb_decoder(16#41#)) OR
 					(reg_q2014 AND symb_decoder(16#65#)) OR
 					(reg_q2014 AND symb_decoder(16#30#)) OR
 					(reg_q2014 AND symb_decoder(16#36#)) OR
 					(reg_q2014 AND symb_decoder(16#45#)) OR
 					(reg_q2014 AND symb_decoder(16#42#));
reg_q1100_in <= (reg_q1098 AND symb_decoder(16#74#)) OR
 					(reg_q1098 AND symb_decoder(16#54#));
reg_q1102_in <= (reg_q1100 AND symb_decoder(16#54#)) OR
 					(reg_q1100 AND symb_decoder(16#74#));
reg_q722_in <= (reg_q720 AND symb_decoder(16#52#)) OR
 					(reg_q720 AND symb_decoder(16#72#));
reg_q724_in <= (reg_q722 AND symb_decoder(16#4f#)) OR
 					(reg_q722 AND symb_decoder(16#6f#));
reg_q1073_in <= (reg_q1071 AND symb_decoder(16#4e#)) OR
 					(reg_q1071 AND symb_decoder(16#6e#));
reg_q1075_in <= (reg_q1073 AND symb_decoder(16#41#)) OR
 					(reg_q1073 AND symb_decoder(16#61#));
reg_q2044_in <= (reg_q2042 AND symb_decoder(16#61#)) OR
 					(reg_q2042 AND symb_decoder(16#37#)) OR
 					(reg_q2042 AND symb_decoder(16#44#)) OR
 					(reg_q2042 AND symb_decoder(16#63#)) OR
 					(reg_q2042 AND symb_decoder(16#62#)) OR
 					(reg_q2042 AND symb_decoder(16#42#)) OR
 					(reg_q2042 AND symb_decoder(16#31#)) OR
 					(reg_q2042 AND symb_decoder(16#45#)) OR
 					(reg_q2042 AND symb_decoder(16#35#)) OR
 					(reg_q2042 AND symb_decoder(16#34#)) OR
 					(reg_q2042 AND symb_decoder(16#46#)) OR
 					(reg_q2042 AND symb_decoder(16#38#)) OR
 					(reg_q2042 AND symb_decoder(16#33#)) OR
 					(reg_q2042 AND symb_decoder(16#39#)) OR
 					(reg_q2042 AND symb_decoder(16#32#)) OR
 					(reg_q2042 AND symb_decoder(16#30#)) OR
 					(reg_q2042 AND symb_decoder(16#36#)) OR
 					(reg_q2042 AND symb_decoder(16#43#)) OR
 					(reg_q2042 AND symb_decoder(16#66#)) OR
 					(reg_q2042 AND symb_decoder(16#65#)) OR
 					(reg_q2042 AND symb_decoder(16#64#)) OR
 					(reg_q2042 AND symb_decoder(16#41#));
reg_q2046_in <= (reg_q2044 AND symb_decoder(16#63#)) OR
 					(reg_q2044 AND symb_decoder(16#46#)) OR
 					(reg_q2044 AND symb_decoder(16#64#)) OR
 					(reg_q2044 AND symb_decoder(16#45#)) OR
 					(reg_q2044 AND symb_decoder(16#41#)) OR
 					(reg_q2044 AND symb_decoder(16#38#)) OR
 					(reg_q2044 AND symb_decoder(16#66#)) OR
 					(reg_q2044 AND symb_decoder(16#43#)) OR
 					(reg_q2044 AND symb_decoder(16#32#)) OR
 					(reg_q2044 AND symb_decoder(16#30#)) OR
 					(reg_q2044 AND symb_decoder(16#42#)) OR
 					(reg_q2044 AND symb_decoder(16#34#)) OR
 					(reg_q2044 AND symb_decoder(16#36#)) OR
 					(reg_q2044 AND symb_decoder(16#65#)) OR
 					(reg_q2044 AND symb_decoder(16#35#)) OR
 					(reg_q2044 AND symb_decoder(16#37#)) OR
 					(reg_q2044 AND symb_decoder(16#44#)) OR
 					(reg_q2044 AND symb_decoder(16#62#)) OR
 					(reg_q2044 AND symb_decoder(16#33#)) OR
 					(reg_q2044 AND symb_decoder(16#61#)) OR
 					(reg_q2044 AND symb_decoder(16#39#)) OR
 					(reg_q2044 AND symb_decoder(16#31#));
reg_q258_in <= (reg_q256 AND symb_decoder(16#52#)) OR
 					(reg_q256 AND symb_decoder(16#72#));
reg_q260_in <= (reg_q258 AND symb_decoder(16#54#)) OR
 					(reg_q258 AND symb_decoder(16#74#));
reg_q236_in <= (reg_q236 AND symb_decoder(16#0a#)) OR
 					(reg_q236 AND symb_decoder(16#20#)) OR
 					(reg_q236 AND symb_decoder(16#09#)) OR
 					(reg_q236 AND symb_decoder(16#0d#)) OR
 					(reg_q236 AND symb_decoder(16#0c#)) OR
 					(reg_q234 AND symb_decoder(16#0a#)) OR
 					(reg_q234 AND symb_decoder(16#20#)) OR
 					(reg_q234 AND symb_decoder(16#0d#)) OR
 					(reg_q234 AND symb_decoder(16#09#)) OR
 					(reg_q234 AND symb_decoder(16#0c#));
reg_q1800_in <= (reg_q1798 AND symb_decoder(16#22#));
reg_q1802_in <= (reg_q1800 AND symb_decoder(16#0c#)) OR
 					(reg_q1800 AND symb_decoder(16#0a#)) OR
 					(reg_q1800 AND symb_decoder(16#0d#)) OR
 					(reg_q1800 AND symb_decoder(16#20#)) OR
 					(reg_q1800 AND symb_decoder(16#09#)) OR
 					(reg_q1802 AND symb_decoder(16#20#)) OR
 					(reg_q1802 AND symb_decoder(16#0d#)) OR
 					(reg_q1802 AND symb_decoder(16#0c#)) OR
 					(reg_q1802 AND symb_decoder(16#0a#)) OR
 					(reg_q1802 AND symb_decoder(16#09#));
reg_q145_in <= (reg_q143 AND symb_decoder(16#56#)) OR
 					(reg_q143 AND symb_decoder(16#76#));
reg_q1723_in <= (reg_q1721 AND symb_decoder(16#73#)) OR
 					(reg_q1721 AND symb_decoder(16#53#));
reg_q511_in <= (reg_q511 AND symb_decoder(16#30#)) OR
 					(reg_q511 AND symb_decoder(16#39#)) OR
 					(reg_q511 AND symb_decoder(16#34#)) OR
 					(reg_q511 AND symb_decoder(16#33#)) OR
 					(reg_q511 AND symb_decoder(16#36#)) OR
 					(reg_q511 AND symb_decoder(16#32#)) OR
 					(reg_q511 AND symb_decoder(16#35#)) OR
 					(reg_q511 AND symb_decoder(16#37#)) OR
 					(reg_q511 AND symb_decoder(16#38#)) OR
 					(reg_q511 AND symb_decoder(16#31#)) OR
 					(reg_q509 AND symb_decoder(16#35#)) OR
 					(reg_q509 AND symb_decoder(16#32#)) OR
 					(reg_q509 AND symb_decoder(16#30#)) OR
 					(reg_q509 AND symb_decoder(16#36#)) OR
 					(reg_q509 AND symb_decoder(16#37#)) OR
 					(reg_q509 AND symb_decoder(16#33#)) OR
 					(reg_q509 AND symb_decoder(16#34#)) OR
 					(reg_q509 AND symb_decoder(16#31#)) OR
 					(reg_q509 AND symb_decoder(16#38#)) OR
 					(reg_q509 AND symb_decoder(16#39#));
reg_q1010_in <= (reg_q1010 AND symb_decoder(16#0a#)) OR
 					(reg_q1010 AND symb_decoder(16#0c#)) OR
 					(reg_q1010 AND symb_decoder(16#0d#)) OR
 					(reg_q1010 AND symb_decoder(16#09#)) OR
 					(reg_q1010 AND symb_decoder(16#20#)) OR
 					(reg_q1008 AND symb_decoder(16#20#)) OR
 					(reg_q1008 AND symb_decoder(16#0c#)) OR
 					(reg_q1008 AND symb_decoder(16#0d#)) OR
 					(reg_q1008 AND symb_decoder(16#0a#)) OR
 					(reg_q1008 AND symb_decoder(16#09#));
reg_q555_in <= (reg_q553 AND symb_decoder(16#45#)) OR
 					(reg_q553 AND symb_decoder(16#65#));
reg_q167_in <= (reg_q165 AND symb_decoder(16#3a#));
reg_q169_in <= (reg_q167 AND symb_decoder(16#31#)) OR
 					(reg_q167 AND symb_decoder(16#39#)) OR
 					(reg_q167 AND symb_decoder(16#35#)) OR
 					(reg_q167 AND symb_decoder(16#34#)) OR
 					(reg_q167 AND symb_decoder(16#38#)) OR
 					(reg_q167 AND symb_decoder(16#33#)) OR
 					(reg_q167 AND symb_decoder(16#30#)) OR
 					(reg_q167 AND symb_decoder(16#36#)) OR
 					(reg_q167 AND symb_decoder(16#32#)) OR
 					(reg_q167 AND symb_decoder(16#37#)) OR
 					(reg_q169 AND symb_decoder(16#38#)) OR
 					(reg_q169 AND symb_decoder(16#35#)) OR
 					(reg_q169 AND symb_decoder(16#31#)) OR
 					(reg_q169 AND symb_decoder(16#36#)) OR
 					(reg_q169 AND symb_decoder(16#32#)) OR
 					(reg_q169 AND symb_decoder(16#34#)) OR
 					(reg_q169 AND symb_decoder(16#39#)) OR
 					(reg_q169 AND symb_decoder(16#30#)) OR
 					(reg_q169 AND symb_decoder(16#37#)) OR
 					(reg_q169 AND symb_decoder(16#33#));
reg_q2304_in <= (reg_q2302 AND symb_decoder(16#52#)) OR
 					(reg_q2302 AND symb_decoder(16#72#));
reg_q2306_in <= (reg_q2304 AND symb_decoder(16#65#)) OR
 					(reg_q2304 AND symb_decoder(16#45#));
reg_q2223_in <= (reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2222 AND symb_decoder(16#2f#));
reg_q1171_in <= (reg_q1169 AND symb_decoder(16#52#)) OR
 					(reg_q1169 AND symb_decoder(16#72#));
reg_q1173_in <= (reg_q1171 AND symb_decoder(16#73#)) OR
 					(reg_q1171 AND symb_decoder(16#53#));
reg_q1520_in <= (reg_q1520 AND symb_decoder(16#34#)) OR
 					(reg_q1520 AND symb_decoder(16#38#)) OR
 					(reg_q1520 AND symb_decoder(16#32#)) OR
 					(reg_q1520 AND symb_decoder(16#33#)) OR
 					(reg_q1520 AND symb_decoder(16#31#)) OR
 					(reg_q1520 AND symb_decoder(16#36#)) OR
 					(reg_q1520 AND symb_decoder(16#37#)) OR
 					(reg_q1520 AND symb_decoder(16#39#)) OR
 					(reg_q1520 AND symb_decoder(16#30#)) OR
 					(reg_q1520 AND symb_decoder(16#35#)) OR
 					(reg_q1518 AND symb_decoder(16#31#)) OR
 					(reg_q1518 AND symb_decoder(16#36#)) OR
 					(reg_q1518 AND symb_decoder(16#37#)) OR
 					(reg_q1518 AND symb_decoder(16#34#)) OR
 					(reg_q1518 AND symb_decoder(16#33#)) OR
 					(reg_q1518 AND symb_decoder(16#35#)) OR
 					(reg_q1518 AND symb_decoder(16#39#)) OR
 					(reg_q1518 AND symb_decoder(16#30#)) OR
 					(reg_q1518 AND symb_decoder(16#38#)) OR
 					(reg_q1518 AND symb_decoder(16#32#));
reg_q147_in <= (reg_q145 AND symb_decoder(16#45#)) OR
 					(reg_q145 AND symb_decoder(16#65#));
reg_q79_in <= (reg_q77 AND symb_decoder(16#53#)) OR
 					(reg_q77 AND symb_decoder(16#73#));
reg_q81_in <= (reg_q79 AND symb_decoder(16#57#)) OR
 					(reg_q79 AND symb_decoder(16#77#));
reg_q242_in <= (reg_q240 AND symb_decoder(16#41#)) OR
 					(reg_q240 AND symb_decoder(16#61#));
reg_q244_in <= (reg_q242 AND symb_decoder(16#52#)) OR
 					(reg_q242 AND symb_decoder(16#72#));
reg_q1911_in <= (reg_q1909 AND symb_decoder(16#31#));
reg_q1913_in <= (reg_q1911 AND symb_decoder(16#2a#));
reg_q190_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q189 AND symb_decoder(16#72#)) OR
 					(reg_q189 AND symb_decoder(16#52#));
reg_q2024_in <= (reg_q2022 AND symb_decoder(16#35#)) OR
 					(reg_q2022 AND symb_decoder(16#65#)) OR
 					(reg_q2022 AND symb_decoder(16#33#)) OR
 					(reg_q2022 AND symb_decoder(16#41#)) OR
 					(reg_q2022 AND symb_decoder(16#37#)) OR
 					(reg_q2022 AND symb_decoder(16#31#)) OR
 					(reg_q2022 AND symb_decoder(16#36#)) OR
 					(reg_q2022 AND symb_decoder(16#46#)) OR
 					(reg_q2022 AND symb_decoder(16#42#)) OR
 					(reg_q2022 AND symb_decoder(16#45#)) OR
 					(reg_q2022 AND symb_decoder(16#61#)) OR
 					(reg_q2022 AND symb_decoder(16#30#)) OR
 					(reg_q2022 AND symb_decoder(16#44#)) OR
 					(reg_q2022 AND symb_decoder(16#66#)) OR
 					(reg_q2022 AND symb_decoder(16#62#)) OR
 					(reg_q2022 AND symb_decoder(16#38#)) OR
 					(reg_q2022 AND symb_decoder(16#39#)) OR
 					(reg_q2022 AND symb_decoder(16#32#)) OR
 					(reg_q2022 AND symb_decoder(16#43#)) OR
 					(reg_q2022 AND symb_decoder(16#34#)) OR
 					(reg_q2022 AND symb_decoder(16#63#)) OR
 					(reg_q2022 AND symb_decoder(16#64#));
reg_q2026_in <= (reg_q2024 AND symb_decoder(16#44#)) OR
 					(reg_q2024 AND symb_decoder(16#65#)) OR
 					(reg_q2024 AND symb_decoder(16#32#)) OR
 					(reg_q2024 AND symb_decoder(16#45#)) OR
 					(reg_q2024 AND symb_decoder(16#66#)) OR
 					(reg_q2024 AND symb_decoder(16#63#)) OR
 					(reg_q2024 AND symb_decoder(16#41#)) OR
 					(reg_q2024 AND symb_decoder(16#42#)) OR
 					(reg_q2024 AND symb_decoder(16#36#)) OR
 					(reg_q2024 AND symb_decoder(16#61#)) OR
 					(reg_q2024 AND symb_decoder(16#34#)) OR
 					(reg_q2024 AND symb_decoder(16#35#)) OR
 					(reg_q2024 AND symb_decoder(16#38#)) OR
 					(reg_q2024 AND symb_decoder(16#43#)) OR
 					(reg_q2024 AND symb_decoder(16#64#)) OR
 					(reg_q2024 AND symb_decoder(16#46#)) OR
 					(reg_q2024 AND symb_decoder(16#30#)) OR
 					(reg_q2024 AND symb_decoder(16#37#)) OR
 					(reg_q2024 AND symb_decoder(16#33#)) OR
 					(reg_q2024 AND symb_decoder(16#39#)) OR
 					(reg_q2024 AND symb_decoder(16#31#)) OR
 					(reg_q2024 AND symb_decoder(16#62#));
reg_q1159_in <= (reg_q1157 AND symb_decoder(16#6f#)) OR
 					(reg_q1157 AND symb_decoder(16#4f#));
reg_q1161_in <= (reg_q1159 AND symb_decoder(16#73#)) OR
 					(reg_q1159 AND symb_decoder(16#53#));
reg_q1918_in <= (reg_q2757 AND symb_decoder(16#2a#));
reg_q1766_in <= (reg_q1764 AND symb_decoder(16#4c#)) OR
 					(reg_q1764 AND symb_decoder(16#6c#));
reg_q1715_in <= (reg_q1715 AND symb_decoder(16#30#)) OR
 					(reg_q1715 AND symb_decoder(16#39#)) OR
 					(reg_q1715 AND symb_decoder(16#31#)) OR
 					(reg_q1715 AND symb_decoder(16#34#)) OR
 					(reg_q1715 AND symb_decoder(16#36#)) OR
 					(reg_q1715 AND symb_decoder(16#32#)) OR
 					(reg_q1715 AND symb_decoder(16#33#)) OR
 					(reg_q1715 AND symb_decoder(16#37#)) OR
 					(reg_q1715 AND symb_decoder(16#35#)) OR
 					(reg_q1715 AND symb_decoder(16#38#)) OR
 					(reg_q1713 AND symb_decoder(16#38#)) OR
 					(reg_q1713 AND symb_decoder(16#33#)) OR
 					(reg_q1713 AND symb_decoder(16#39#)) OR
 					(reg_q1713 AND symb_decoder(16#36#)) OR
 					(reg_q1713 AND symb_decoder(16#34#)) OR
 					(reg_q1713 AND symb_decoder(16#30#)) OR
 					(reg_q1713 AND symb_decoder(16#31#)) OR
 					(reg_q1713 AND symb_decoder(16#35#)) OR
 					(reg_q1713 AND symb_decoder(16#37#)) OR
 					(reg_q1713 AND symb_decoder(16#32#));
reg_q530_in <= (reg_q526 AND symb_decoder(16#0d#)) OR
 					(reg_q540 AND symb_decoder(16#0d#));
reg_q32_in <= (reg_q30 AND symb_decoder(16#52#)) OR
 					(reg_q30 AND symb_decoder(16#72#));
reg_q34_in <= (reg_q32 AND symb_decoder(16#6f#)) OR
 					(reg_q32 AND symb_decoder(16#4f#));
reg_q990_in <= (reg_q988 AND symb_decoder(16#72#)) OR
 					(reg_q988 AND symb_decoder(16#52#));
reg_q992_in <= (reg_q990 AND symb_decoder(16#52#)) OR
 					(reg_q990 AND symb_decoder(16#72#));
reg_q18_in <= (reg_q16 AND symb_decoder(16#52#)) OR
 					(reg_q16 AND symb_decoder(16#72#));
reg_q20_in <= (reg_q18 AND symb_decoder(16#4f#)) OR
 					(reg_q18 AND symb_decoder(16#6f#));
reg_q9_in <= (reg_q7 AND symb_decoder(16#77#)) OR
 					(reg_q7 AND symb_decoder(16#57#));
reg_q11_in <= (reg_q9 AND symb_decoder(16#64#)) OR
 					(reg_q9 AND symb_decoder(16#44#));
reg_q1735_in <= (reg_q1735 AND symb_decoder(16#0a#)) OR
 					(reg_q1735 AND symb_decoder(16#0d#)) OR
 					(reg_q1735 AND symb_decoder(16#20#)) OR
 					(reg_q1735 AND symb_decoder(16#09#)) OR
 					(reg_q1735 AND symb_decoder(16#0c#)) OR
 					(reg_q1733 AND symb_decoder(16#20#)) OR
 					(reg_q1733 AND symb_decoder(16#0a#)) OR
 					(reg_q1733 AND symb_decoder(16#09#)) OR
 					(reg_q1733 AND symb_decoder(16#0c#)) OR
 					(reg_q1733 AND symb_decoder(16#0d#));
reg_q1737_in <= (reg_q1735 AND symb_decoder(16#4f#)) OR
 					(reg_q1735 AND symb_decoder(16#6f#));
reg_q1331_in <= (reg_q1329 AND symb_decoder(16#53#)) OR
 					(reg_q1329 AND symb_decoder(16#73#));
reg_q1333_in <= (reg_q1331 AND symb_decoder(16#0d#)) OR
 					(reg_q1331 AND symb_decoder(16#0a#)) OR
 					(reg_q1331 AND symb_decoder(16#09#)) OR
 					(reg_q1331 AND symb_decoder(16#20#)) OR
 					(reg_q1331 AND symb_decoder(16#0c#)) OR
 					(reg_q1333 AND symb_decoder(16#0d#)) OR
 					(reg_q1333 AND symb_decoder(16#0c#)) OR
 					(reg_q1333 AND symb_decoder(16#0a#)) OR
 					(reg_q1333 AND symb_decoder(16#09#)) OR
 					(reg_q1333 AND symb_decoder(16#20#));
reg_q1713_in <= (reg_q1711 AND symb_decoder(16#56#)) OR
 					(reg_q1711 AND symb_decoder(16#76#));
reg_q373_in <= (reg_q395 AND symb_decoder(16#4b#)) OR
 					(reg_q395 AND symb_decoder(16#6b#)) OR
 					(reg_q369 AND symb_decoder(16#6b#)) OR
 					(reg_q369 AND symb_decoder(16#4b#));
reg_q375_in <= (reg_q373 AND symb_decoder(16#49#)) OR
 					(reg_q373 AND symb_decoder(16#69#));
reg_q2395_in <= (reg_q2393 AND symb_decoder(16#65#)) OR
 					(reg_q2393 AND symb_decoder(16#45#));
reg_q2397_in <= (reg_q2395 AND symb_decoder(16#73#)) OR
 					(reg_q2395 AND symb_decoder(16#53#));
reg_q2601_in <= (reg_q2599 AND symb_decoder(16#45#)) OR
 					(reg_q2599 AND symb_decoder(16#65#));
reg_q77_in <= (reg_q75 AND symb_decoder(16#73#)) OR
 					(reg_q75 AND symb_decoder(16#53#));
reg_q2694_in <= (reg_q2692 AND symb_decoder(16#53#)) OR
 					(reg_q2692 AND symb_decoder(16#73#));
reg_q2696_in <= (reg_q2694 AND symb_decoder(16#c0#));
reg_q2310_in <= (reg_q2308 AND symb_decoder(16#74#)) OR
 					(reg_q2308 AND symb_decoder(16#54#));
reg_q1012_in <= (reg_q1010 AND symb_decoder(16#66#)) OR
 					(reg_q1010 AND symb_decoder(16#46#));
reg_q1014_in <= (reg_q1012 AND symb_decoder(16#52#)) OR
 					(reg_q1012 AND symb_decoder(16#72#));
reg_q1193_in <= (reg_q1191 AND symb_decoder(16#65#)) OR
 					(reg_q1191 AND symb_decoder(16#45#));
reg_q1195_in <= (reg_q1193 AND symb_decoder(16#52#)) OR
 					(reg_q1193 AND symb_decoder(16#72#));
reg_q2407_in <= (reg_q2405 AND symb_decoder(16#76#)) OR
 					(reg_q2405 AND symb_decoder(16#56#));
reg_q2409_in <= (reg_q2407 AND symb_decoder(16#65#)) OR
 					(reg_q2407 AND symb_decoder(16#45#));
reg_q2718_in <= (reg_q2716 AND symb_decoder(16#65#)) OR
 					(reg_q2716 AND symb_decoder(16#45#));
reg_q2720_in <= (reg_q2718 AND symb_decoder(16#59#)) OR
 					(reg_q2718 AND symb_decoder(16#79#));
reg_q216_in <= (reg_q214 AND symb_decoder(16#3b#));
reg_q1327_in <= (reg_q1325 AND symb_decoder(16#68#)) OR
 					(reg_q1325 AND symb_decoder(16#48#));
reg_q551_in <= (reg_q549 AND symb_decoder(16#23#));
reg_q2048_in <= (reg_q2046 AND symb_decoder(16#35#)) OR
 					(reg_q2046 AND symb_decoder(16#66#)) OR
 					(reg_q2046 AND symb_decoder(16#43#)) OR
 					(reg_q2046 AND symb_decoder(16#45#)) OR
 					(reg_q2046 AND symb_decoder(16#63#)) OR
 					(reg_q2046 AND symb_decoder(16#44#)) OR
 					(reg_q2046 AND symb_decoder(16#36#)) OR
 					(reg_q2046 AND symb_decoder(16#42#)) OR
 					(reg_q2046 AND symb_decoder(16#37#)) OR
 					(reg_q2046 AND symb_decoder(16#46#)) OR
 					(reg_q2046 AND symb_decoder(16#41#)) OR
 					(reg_q2046 AND symb_decoder(16#31#)) OR
 					(reg_q2046 AND symb_decoder(16#64#)) OR
 					(reg_q2046 AND symb_decoder(16#34#)) OR
 					(reg_q2046 AND symb_decoder(16#38#)) OR
 					(reg_q2046 AND symb_decoder(16#39#)) OR
 					(reg_q2046 AND symb_decoder(16#65#)) OR
 					(reg_q2046 AND symb_decoder(16#30#)) OR
 					(reg_q2046 AND symb_decoder(16#62#)) OR
 					(reg_q2046 AND symb_decoder(16#33#)) OR
 					(reg_q2046 AND symb_decoder(16#61#)) OR
 					(reg_q2046 AND symb_decoder(16#32#));
reg_q105_in <= (reg_q103 AND symb_decoder(16#44#)) OR
 					(reg_q103 AND symb_decoder(16#64#));
reg_q1484_in <= (reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q1483 AND symb_decoder(16#57#)) OR
 					(reg_q1483 AND symb_decoder(16#77#));
reg_q250_in <= (reg_q248 AND symb_decoder(16#44#)) OR
 					(reg_q248 AND symb_decoder(16#64#));
reg_q252_in <= (reg_q250 AND symb_decoder(16#09#)) OR
 					(reg_q250 AND symb_decoder(16#0a#)) OR
 					(reg_q250 AND symb_decoder(16#20#)) OR
 					(reg_q250 AND symb_decoder(16#0c#)) OR
 					(reg_q250 AND symb_decoder(16#0d#)) OR
 					(reg_q252 AND symb_decoder(16#0a#)) OR
 					(reg_q252 AND symb_decoder(16#0d#)) OR
 					(reg_q252 AND symb_decoder(16#0c#)) OR
 					(reg_q252 AND symb_decoder(16#20#)) OR
 					(reg_q252 AND symb_decoder(16#09#));
reg_q2415_in <= (reg_q2413 AND symb_decoder(16#6c#)) OR
 					(reg_q2413 AND symb_decoder(16#4c#));
reg_q2010_in <= (reg_q2008 AND symb_decoder(16#66#)) OR
 					(reg_q2008 AND symb_decoder(16#64#)) OR
 					(reg_q2008 AND symb_decoder(16#39#)) OR
 					(reg_q2008 AND symb_decoder(16#37#)) OR
 					(reg_q2008 AND symb_decoder(16#62#)) OR
 					(reg_q2008 AND symb_decoder(16#43#)) OR
 					(reg_q2008 AND symb_decoder(16#45#)) OR
 					(reg_q2008 AND symb_decoder(16#34#)) OR
 					(reg_q2008 AND symb_decoder(16#33#)) OR
 					(reg_q2008 AND symb_decoder(16#61#)) OR
 					(reg_q2008 AND symb_decoder(16#41#)) OR
 					(reg_q2008 AND symb_decoder(16#63#)) OR
 					(reg_q2008 AND symb_decoder(16#32#)) OR
 					(reg_q2008 AND symb_decoder(16#30#)) OR
 					(reg_q2008 AND symb_decoder(16#38#)) OR
 					(reg_q2008 AND symb_decoder(16#31#)) OR
 					(reg_q2008 AND symb_decoder(16#65#)) OR
 					(reg_q2008 AND symb_decoder(16#42#)) OR
 					(reg_q2008 AND symb_decoder(16#35#)) OR
 					(reg_q2008 AND symb_decoder(16#36#)) OR
 					(reg_q2008 AND symb_decoder(16#44#)) OR
 					(reg_q2008 AND symb_decoder(16#46#));
reg_q2585_in <= (reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2584 AND symb_decoder(16#7c#));
reg_q2682_in <= (reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2681 AND symb_decoder(16#c0#));
reg_q996_in <= (reg_q994 AND symb_decoder(16#4e#)) OR
 					(reg_q994 AND symb_decoder(16#6e#));
reg_q998_in <= (reg_q996 AND symb_decoder(16#67#)) OR
 					(reg_q996 AND symb_decoder(16#47#));
reg_q1808_in <= (reg_q1806 AND symb_decoder(16#2e#));
reg_q1810_in <= (reg_q1808 AND symb_decoder(16#34#)) OR
 					(reg_q1808 AND symb_decoder(16#36#)) OR
 					(reg_q1808 AND symb_decoder(16#33#)) OR
 					(reg_q1808 AND symb_decoder(16#30#)) OR
 					(reg_q1808 AND symb_decoder(16#35#)) OR
 					(reg_q1808 AND symb_decoder(16#32#)) OR
 					(reg_q1808 AND symb_decoder(16#31#)) OR
 					(reg_q1808 AND symb_decoder(16#38#)) OR
 					(reg_q1808 AND symb_decoder(16#37#)) OR
 					(reg_q1808 AND symb_decoder(16#39#)) OR
 					(reg_q1810 AND symb_decoder(16#37#)) OR
 					(reg_q1810 AND symb_decoder(16#36#)) OR
 					(reg_q1810 AND symb_decoder(16#38#)) OR
 					(reg_q1810 AND symb_decoder(16#35#)) OR
 					(reg_q1810 AND symb_decoder(16#34#)) OR
 					(reg_q1810 AND symb_decoder(16#32#)) OR
 					(reg_q1810 AND symb_decoder(16#39#)) OR
 					(reg_q1810 AND symb_decoder(16#31#)) OR
 					(reg_q1810 AND symb_decoder(16#33#)) OR
 					(reg_q1810 AND symb_decoder(16#30#));
reg_q1725_in <= (reg_q1723 AND symb_decoder(16#45#)) OR
 					(reg_q1723 AND symb_decoder(16#65#));
reg_q1727_in <= (reg_q1725 AND symb_decoder(16#72#)) OR
 					(reg_q1725 AND symb_decoder(16#52#));
reg_q1743_in <= (reg_q1741 AND symb_decoder(16#49#)) OR
 					(reg_q1741 AND symb_decoder(16#69#));
reg_q1745_in <= (reg_q1743 AND symb_decoder(16#4e#)) OR
 					(reg_q1743 AND symb_decoder(16#6e#));
reg_q204_in <= (reg_q204 AND symb_decoder(16#0a#)) OR
 					(reg_q204 AND symb_decoder(16#0d#)) OR
 					(reg_q204 AND symb_decoder(16#20#)) OR
 					(reg_q204 AND symb_decoder(16#0c#)) OR
 					(reg_q204 AND symb_decoder(16#09#)) OR
 					(reg_q202 AND symb_decoder(16#0c#)) OR
 					(reg_q202 AND symb_decoder(16#09#)) OR
 					(reg_q202 AND symb_decoder(16#0a#)) OR
 					(reg_q202 AND symb_decoder(16#20#)) OR
 					(reg_q202 AND symb_decoder(16#0d#));
reg_q206_in <= (reg_q204 AND symb_decoder(16#76#)) OR
 					(reg_q204 AND symb_decoder(16#56#));
reg_q2393_in <= (reg_q2391 AND symb_decoder(16#63#)) OR
 					(reg_q2391 AND symb_decoder(16#43#));
reg_q1762_in <= (reg_q1760 AND symb_decoder(16#4f#)) OR
 					(reg_q1760 AND symb_decoder(16#6f#));
reg_q1764_in <= (reg_q1762 AND symb_decoder(16#6c#)) OR
 					(reg_q1762 AND symb_decoder(16#4c#));
reg_q868_in <= (reg_q866 AND symb_decoder(16#6a#)) OR
 					(reg_q866 AND symb_decoder(16#4a#));
reg_q2684_in <= (reg_q2682 AND symb_decoder(16#73#)) OR
 					(reg_q2682 AND symb_decoder(16#53#));
reg_q2686_in <= (reg_q2684 AND symb_decoder(16#74#)) OR
 					(reg_q2684 AND symb_decoder(16#54#));
reg_q746_in <= (reg_q746 AND symb_decoder(16#0c#)) OR
 					(reg_q746 AND symb_decoder(16#0a#)) OR
 					(reg_q746 AND symb_decoder(16#20#)) OR
 					(reg_q746 AND symb_decoder(16#09#)) OR
 					(reg_q746 AND symb_decoder(16#0d#)) OR
 					(reg_q744 AND symb_decoder(16#0c#)) OR
 					(reg_q744 AND symb_decoder(16#0a#)) OR
 					(reg_q744 AND symb_decoder(16#09#)) OR
 					(reg_q744 AND symb_decoder(16#0d#)) OR
 					(reg_q744 AND symb_decoder(16#20#));
reg_q87_in <= (reg_q85 AND symb_decoder(16#64#)) OR
 					(reg_q85 AND symb_decoder(16#44#));
reg_q89_in <= (reg_q87 AND symb_decoder(16#0d#)) OR
 					(reg_q87 AND symb_decoder(16#0c#)) OR
 					(reg_q87 AND symb_decoder(16#0a#)) OR
 					(reg_q87 AND symb_decoder(16#20#)) OR
 					(reg_q87 AND symb_decoder(16#09#)) OR
 					(reg_q89 AND symb_decoder(16#0a#)) OR
 					(reg_q89 AND symb_decoder(16#0c#)) OR
 					(reg_q89 AND symb_decoder(16#20#)) OR
 					(reg_q89 AND symb_decoder(16#0d#)) OR
 					(reg_q89 AND symb_decoder(16#09#));
reg_q5_in <= (reg_q3 AND symb_decoder(16#73#)) OR
 					(reg_q3 AND symb_decoder(16#53#));
reg_q1165_in <= (reg_q1165 AND symb_decoder(16#0c#)) OR
 					(reg_q1165 AND symb_decoder(16#0d#)) OR
 					(reg_q1165 AND symb_decoder(16#20#)) OR
 					(reg_q1165 AND symb_decoder(16#0a#)) OR
 					(reg_q1165 AND symb_decoder(16#09#)) OR
 					(reg_q1163 AND symb_decoder(16#20#)) OR
 					(reg_q1163 AND symb_decoder(16#09#)) OR
 					(reg_q1163 AND symb_decoder(16#0a#)) OR
 					(reg_q1163 AND symb_decoder(16#0c#)) OR
 					(reg_q1163 AND symb_decoder(16#0d#));
reg_q1167_in <= (reg_q1165 AND symb_decoder(16#56#)) OR
 					(reg_q1165 AND symb_decoder(16#76#));
reg_q1208_in <= (reg_q1206 AND symb_decoder(16#3b#));
reg_q1210_in <= (reg_q1208 AND symb_decoder(16#32#)) OR
 					(reg_q1208 AND symb_decoder(16#39#)) OR
 					(reg_q1208 AND symb_decoder(16#38#)) OR
 					(reg_q1208 AND symb_decoder(16#31#)) OR
 					(reg_q1208 AND symb_decoder(16#30#)) OR
 					(reg_q1208 AND symb_decoder(16#33#)) OR
 					(reg_q1208 AND symb_decoder(16#34#)) OR
 					(reg_q1208 AND symb_decoder(16#36#)) OR
 					(reg_q1208 AND symb_decoder(16#37#)) OR
 					(reg_q1208 AND symb_decoder(16#35#)) OR
 					(reg_q1210 AND symb_decoder(16#31#)) OR
 					(reg_q1210 AND symb_decoder(16#37#)) OR
 					(reg_q1210 AND symb_decoder(16#34#)) OR
 					(reg_q1210 AND symb_decoder(16#39#)) OR
 					(reg_q1210 AND symb_decoder(16#32#)) OR
 					(reg_q1210 AND symb_decoder(16#30#)) OR
 					(reg_q1210 AND symb_decoder(16#38#)) OR
 					(reg_q1210 AND symb_decoder(16#35#)) OR
 					(reg_q1210 AND symb_decoder(16#33#)) OR
 					(reg_q1210 AND symb_decoder(16#36#));
reg_q254_in <= (reg_q252 AND symb_decoder(16#70#)) OR
 					(reg_q252 AND symb_decoder(16#50#));
reg_q1313_in <= (reg_q1311 AND symb_decoder(16#45#)) OR
 					(reg_q1311 AND symb_decoder(16#65#));
reg_q1132_in <= (reg_q1130 AND symb_decoder(16#4c#)) OR
 					(reg_q1130 AND symb_decoder(16#6c#));
reg_q2308_in <= (reg_q2306 AND symb_decoder(16#6e#)) OR
 					(reg_q2306 AND symb_decoder(16#4e#));
reg_q702_in <= (reg_q700 AND symb_decoder(16#6c#)) OR
 					(reg_q700 AND symb_decoder(16#4c#));
reg_q1081_in <= (reg_q1081 AND symb_decoder(16#0d#)) OR
 					(reg_q1081 AND symb_decoder(16#09#)) OR
 					(reg_q1081 AND symb_decoder(16#0c#)) OR
 					(reg_q1081 AND symb_decoder(16#20#)) OR
 					(reg_q1081 AND symb_decoder(16#0a#)) OR
 					(reg_q1079 AND symb_decoder(16#0a#)) OR
 					(reg_q1079 AND symb_decoder(16#0c#)) OR
 					(reg_q1079 AND symb_decoder(16#09#)) OR
 					(reg_q1079 AND symb_decoder(16#20#)) OR
 					(reg_q1079 AND symb_decoder(16#0d#));
reg_q988_in <= (reg_q986 AND symb_decoder(16#45#)) OR
 					(reg_q986 AND symb_decoder(16#65#));
reg_q1689_in <= (reg_q1687 AND symb_decoder(16#21#));
reg_q1691_in <= (reg_q1689 AND symb_decoder(16#21#));
reg_q2615_in <= (reg_q2613 AND symb_decoder(16#3a#));
reg_q1514_in <= (reg_q1514 AND symb_decoder(16#0c#)) OR
 					(reg_q1514 AND symb_decoder(16#0d#)) OR
 					(reg_q1514 AND symb_decoder(16#09#)) OR
 					(reg_q1514 AND symb_decoder(16#20#)) OR
 					(reg_q1514 AND symb_decoder(16#0a#)) OR
 					(reg_q1512 AND symb_decoder(16#0d#)) OR
 					(reg_q1512 AND symb_decoder(16#0a#)) OR
 					(reg_q1512 AND symb_decoder(16#0c#)) OR
 					(reg_q1512 AND symb_decoder(16#09#)) OR
 					(reg_q1512 AND symb_decoder(16#20#));
reg_q1516_in <= (reg_q1514 AND symb_decoder(16#30#)) OR
 					(reg_q1514 AND symb_decoder(16#31#)) OR
 					(reg_q1514 AND symb_decoder(16#34#)) OR
 					(reg_q1514 AND symb_decoder(16#39#)) OR
 					(reg_q1514 AND symb_decoder(16#38#)) OR
 					(reg_q1514 AND symb_decoder(16#37#)) OR
 					(reg_q1514 AND symb_decoder(16#36#)) OR
 					(reg_q1514 AND symb_decoder(16#35#)) OR
 					(reg_q1514 AND symb_decoder(16#33#)) OR
 					(reg_q1514 AND symb_decoder(16#32#)) OR
 					(reg_q1516 AND symb_decoder(16#33#)) OR
 					(reg_q1516 AND symb_decoder(16#38#)) OR
 					(reg_q1516 AND symb_decoder(16#37#)) OR
 					(reg_q1516 AND symb_decoder(16#31#)) OR
 					(reg_q1516 AND symb_decoder(16#34#)) OR
 					(reg_q1516 AND symb_decoder(16#32#)) OR
 					(reg_q1516 AND symb_decoder(16#39#)) OR
 					(reg_q1516 AND symb_decoder(16#35#)) OR
 					(reg_q1516 AND symb_decoder(16#36#)) OR
 					(reg_q1516 AND symb_decoder(16#30#));
reg_q740_in <= (reg_q738 AND symb_decoder(16#76#)) OR
 					(reg_q738 AND symb_decoder(16#56#));
reg_q563_in <= (reg_q561 AND symb_decoder(16#52#)) OR
 					(reg_q561 AND symb_decoder(16#72#));
reg_q994_in <= (reg_q992 AND symb_decoder(16#69#)) OR
 					(reg_q992 AND symb_decoder(16#49#));
reg_q2002_in <= (reg_q2000 AND symb_decoder(16#32#)) OR
 					(reg_q2000 AND symb_decoder(16#41#)) OR
 					(reg_q2000 AND symb_decoder(16#66#)) OR
 					(reg_q2000 AND symb_decoder(16#31#)) OR
 					(reg_q2000 AND symb_decoder(16#39#)) OR
 					(reg_q2000 AND symb_decoder(16#33#)) OR
 					(reg_q2000 AND symb_decoder(16#61#)) OR
 					(reg_q2000 AND symb_decoder(16#42#)) OR
 					(reg_q2000 AND symb_decoder(16#46#)) OR
 					(reg_q2000 AND symb_decoder(16#34#)) OR
 					(reg_q2000 AND symb_decoder(16#38#)) OR
 					(reg_q2000 AND symb_decoder(16#63#)) OR
 					(reg_q2000 AND symb_decoder(16#64#)) OR
 					(reg_q2000 AND symb_decoder(16#30#)) OR
 					(reg_q2000 AND symb_decoder(16#36#)) OR
 					(reg_q2000 AND symb_decoder(16#62#)) OR
 					(reg_q2000 AND symb_decoder(16#35#)) OR
 					(reg_q2000 AND symb_decoder(16#44#)) OR
 					(reg_q2000 AND symb_decoder(16#43#)) OR
 					(reg_q2000 AND symb_decoder(16#45#)) OR
 					(reg_q2000 AND symb_decoder(16#65#)) OR
 					(reg_q2000 AND symb_decoder(16#37#));
reg_q708_in <= (reg_q706 AND symb_decoder(16#55#)) OR
 					(reg_q706 AND symb_decoder(16#75#));
reg_q710_in <= (reg_q708 AND symb_decoder(16#53#)) OR
 					(reg_q708 AND symb_decoder(16#73#));
reg_q1185_in <= (reg_q1183 AND symb_decoder(16#2e#));
reg_q2357_in <= (reg_q2355 AND symb_decoder(16#55#)) OR
 					(reg_q2355 AND symb_decoder(16#75#));
reg_q2359_in <= (reg_q2357 AND symb_decoder(16#53#)) OR
 					(reg_q2357 AND symb_decoder(16#73#));
reg_q226_in <= (reg_q224 AND symb_decoder(16#65#)) OR
 					(reg_q224 AND symb_decoder(16#45#));
reg_q228_in <= (reg_q226 AND symb_decoder(16#57#)) OR
 					(reg_q226 AND symb_decoder(16#77#));
reg_q1339_in <= (reg_q1337 AND symb_decoder(16#65#)) OR
 					(reg_q1337 AND symb_decoder(16#45#));
reg_q1341_in <= (reg_q1339 AND symb_decoder(16#61#)) OR
 					(reg_q1339 AND symb_decoder(16#41#));
reg_q1124_in <= (reg_q1122 AND symb_decoder(16#67#)) OR
 					(reg_q1122 AND symb_decoder(16#47#));
reg_q1317_in <= (reg_q1315 AND symb_decoder(16#67#)) OR
 					(reg_q1315 AND symb_decoder(16#47#));
reg_q38_in <= (reg_q36 AND symb_decoder(16#47#)) OR
 					(reg_q36 AND symb_decoder(16#67#));
reg_q673_in <= (reg_q671 AND symb_decoder(16#09#)) OR
 					(reg_q671 AND symb_decoder(16#0a#)) OR
 					(reg_q671 AND symb_decoder(16#0d#)) OR
 					(reg_q671 AND symb_decoder(16#0c#)) OR
 					(reg_q671 AND symb_decoder(16#20#));
reg_q1349_in <= (reg_q1347 AND symb_decoder(16#41#)) OR
 					(reg_q1347 AND symb_decoder(16#61#));
reg_q1351_in <= (reg_q1349 AND symb_decoder(16#65#)) OR
 					(reg_q1349 AND symb_decoder(16#45#));
reg_q1494_in <= (reg_q1492 AND symb_decoder(16#61#)) OR
 					(reg_q1492 AND symb_decoder(16#41#));
reg_q1496_in <= (reg_q1494 AND symb_decoder(16#73#)) OR
 					(reg_q1494 AND symb_decoder(16#53#));
reg_q532_in <= (reg_q530 AND symb_decoder(16#0a#));
reg_q534_in <= (reg_q532 AND symb_decoder(16#31#)) OR
 					(reg_q532 AND symb_decoder(16#32#)) OR
 					(reg_q532 AND symb_decoder(16#35#)) OR
 					(reg_q532 AND symb_decoder(16#37#)) OR
 					(reg_q532 AND symb_decoder(16#34#)) OR
 					(reg_q532 AND symb_decoder(16#36#)) OR
 					(reg_q532 AND symb_decoder(16#33#)) OR
 					(reg_q532 AND symb_decoder(16#30#)) OR
 					(reg_q532 AND symb_decoder(16#39#)) OR
 					(reg_q532 AND symb_decoder(16#38#)) OR
 					(reg_q534 AND symb_decoder(16#35#)) OR
 					(reg_q534 AND symb_decoder(16#33#)) OR
 					(reg_q534 AND symb_decoder(16#30#)) OR
 					(reg_q534 AND symb_decoder(16#32#)) OR
 					(reg_q534 AND symb_decoder(16#37#)) OR
 					(reg_q534 AND symb_decoder(16#31#)) OR
 					(reg_q534 AND symb_decoder(16#34#)) OR
 					(reg_q534 AND symb_decoder(16#38#)) OR
 					(reg_q534 AND symb_decoder(16#39#)) OR
 					(reg_q534 AND symb_decoder(16#36#));
reg_q967_in <= (reg_q965 AND symb_decoder(16#53#));
reg_q955_in <= (reg_q967 AND symb_decoder(16#44#)) OR
 					(reg_q952 AND symb_decoder(16#44#));
reg_q270_in <= (reg_q268 AND symb_decoder(16#55#)) OR
 					(reg_q268 AND symb_decoder(16#75#));
reg_q272_in <= (reg_q270 AND symb_decoder(16#72#)) OR
 					(reg_q270 AND symb_decoder(16#52#));
reg_q734_in <= (reg_q732 AND symb_decoder(16#73#)) OR
 					(reg_q732 AND symb_decoder(16#53#));
reg_q736_in <= (reg_q734 AND symb_decoder(16#65#)) OR
 					(reg_q734 AND symb_decoder(16#45#));
reg_q1004_in <= (reg_q1002 AND symb_decoder(16#69#)) OR
 					(reg_q1002 AND symb_decoder(16#49#));
reg_q1006_in <= (reg_q1004 AND symb_decoder(16#6c#)) OR
 					(reg_q1004 AND symb_decoder(16#4c#));
reg_q1077_in <= (reg_q1075 AND symb_decoder(16#4b#)) OR
 					(reg_q1075 AND symb_decoder(16#6b#));
reg_q1079_in <= (reg_q1077 AND symb_decoder(16#45#)) OR
 					(reg_q1077 AND symb_decoder(16#65#));
reg_q2268_in <= (reg_q2266 AND symb_decoder(16#65#)) OR
 					(reg_q2266 AND symb_decoder(16#45#));
reg_q2270_in <= (reg_q2268 AND symb_decoder(16#72#)) OR
 					(reg_q2268 AND symb_decoder(16#52#));
reg_q2298_in <= (reg_q2296 AND symb_decoder(16#63#)) OR
 					(reg_q2296 AND symb_decoder(16#43#));
reg_q2300_in <= (reg_q2298 AND symb_decoder(16#55#)) OR
 					(reg_q2298 AND symb_decoder(16#75#));
reg_q1905_in <= (reg_q1903 AND symb_decoder(16#4f#));
reg_q1163_in <= (reg_q1161 AND symb_decoder(16#54#)) OR
 					(reg_q1161 AND symb_decoder(16#74#));
reg_q1812_in <= (reg_q1810 AND symb_decoder(16#0d#));
reg_q1814_in <= (reg_q1812 AND symb_decoder(16#0a#));
reg_q1000_in <= (reg_q998 AND symb_decoder(16#20#)) OR
 					(reg_q998 AND symb_decoder(16#0d#)) OR
 					(reg_q998 AND symb_decoder(16#0c#)) OR
 					(reg_q998 AND symb_decoder(16#0a#)) OR
 					(reg_q998 AND symb_decoder(16#09#)) OR
 					(reg_q1000 AND symb_decoder(16#0d#)) OR
 					(reg_q1000 AND symb_decoder(16#20#)) OR
 					(reg_q1000 AND symb_decoder(16#09#)) OR
 					(reg_q1000 AND symb_decoder(16#0a#)) OR
 					(reg_q1000 AND symb_decoder(16#0c#));
reg_q1069_in <= (reg_q1069 AND symb_decoder(16#20#)) OR
 					(reg_q1069 AND symb_decoder(16#0d#)) OR
 					(reg_q1069 AND symb_decoder(16#0c#)) OR
 					(reg_q1069 AND symb_decoder(16#09#)) OR
 					(reg_q1069 AND symb_decoder(16#0a#)) OR
 					(reg_q1067 AND symb_decoder(16#0d#)) OR
 					(reg_q1067 AND symb_decoder(16#0a#)) OR
 					(reg_q1067 AND symb_decoder(16#09#)) OR
 					(reg_q1067 AND symb_decoder(16#0c#)) OR
 					(reg_q1067 AND symb_decoder(16#20#));
reg_q274_in <= (reg_q272 AND symb_decoder(16#0a#)) OR
 					(reg_q272 AND symb_decoder(16#20#)) OR
 					(reg_q272 AND symb_decoder(16#0d#)) OR
 					(reg_q272 AND symb_decoder(16#0c#)) OR
 					(reg_q272 AND symb_decoder(16#09#)) OR
 					(reg_q274 AND symb_decoder(16#0c#)) OR
 					(reg_q274 AND symb_decoder(16#0d#)) OR
 					(reg_q274 AND symb_decoder(16#20#)) OR
 					(reg_q274 AND symb_decoder(16#0a#)) OR
 					(reg_q274 AND symb_decoder(16#09#));
reg_q1794_in <= (reg_q1792 AND symb_decoder(16#47#)) OR
 					(reg_q1792 AND symb_decoder(16#67#));
reg_q1796_in <= (reg_q1794 AND symb_decoder(16#45#)) OR
 					(reg_q1794 AND symb_decoder(16#65#));
reg_q280_in <= (reg_q280 AND symb_decoder(16#20#)) OR
 					(reg_q280 AND symb_decoder(16#0d#)) OR
 					(reg_q280 AND symb_decoder(16#0c#)) OR
 					(reg_q280 AND symb_decoder(16#09#)) OR
 					(reg_q280 AND symb_decoder(16#0a#)) OR
 					(reg_q278 AND symb_decoder(16#0c#)) OR
 					(reg_q278 AND symb_decoder(16#0a#)) OR
 					(reg_q278 AND symb_decoder(16#0d#)) OR
 					(reg_q278 AND symb_decoder(16#20#)) OR
 					(reg_q278 AND symb_decoder(16#09#));
reg_q2347_in <= (reg_q2345 AND symb_decoder(16#73#)) OR
 					(reg_q2345 AND symb_decoder(16#53#));
reg_q2349_in <= (reg_q2347 AND symb_decoder(16#73#)) OR
 					(reg_q2347 AND symb_decoder(16#53#));
reg_q387_in <= (reg_q385 AND symb_decoder(16#6e#)) OR
 					(reg_q385 AND symb_decoder(16#4e#));
reg_q389_in <= (reg_q387 AND symb_decoder(16#45#)) OR
 					(reg_q387 AND symb_decoder(16#65#));
reg_q1343_in <= (reg_q1341 AND symb_decoder(16#54#)) OR
 					(reg_q1341 AND symb_decoder(16#74#));
reg_q1729_in <= (reg_q1727 AND symb_decoder(16#76#)) OR
 					(reg_q1727 AND symb_decoder(16#56#));
reg_q2522_in <= (reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2521 AND symb_decoder(16#3c#));
reg_q2722_in <= (reg_q2720 AND symb_decoder(16#6c#)) OR
 					(reg_q2720 AND symb_decoder(16#4c#));
reg_q2724_in <= (reg_q2722 AND symb_decoder(16#6f#)) OR
 					(reg_q2722 AND symb_decoder(16#4f#));
reg_q1776_in <= (reg_q1774 AND symb_decoder(16#6d#)) OR
 					(reg_q1774 AND symb_decoder(16#4d#));
reg_q2286_in <= (reg_q2284 AND symb_decoder(16#52#)) OR
 					(reg_q2284 AND symb_decoder(16#72#));
reg_q264_in <= (reg_q264 AND symb_decoder(16#09#)) OR
 					(reg_q264 AND symb_decoder(16#20#)) OR
 					(reg_q264 AND symb_decoder(16#0d#)) OR
 					(reg_q264 AND symb_decoder(16#0c#)) OR
 					(reg_q264 AND symb_decoder(16#0a#)) OR
 					(reg_q262 AND symb_decoder(16#0a#)) OR
 					(reg_q262 AND symb_decoder(16#0c#)) OR
 					(reg_q262 AND symb_decoder(16#09#)) OR
 					(reg_q262 AND symb_decoder(16#20#)) OR
 					(reg_q262 AND symb_decoder(16#0d#));
reg_q2373_in <= (reg_q2371 AND symb_decoder(16#54#)) OR
 					(reg_q2371 AND symb_decoder(16#74#));
reg_q2375_in <= (reg_q2373 AND symb_decoder(16#69#)) OR
 					(reg_q2373 AND symb_decoder(16#49#));
reg_q2702_in <= (reg_q2700 AND symb_decoder(16#52#)) OR
 					(reg_q2700 AND symb_decoder(16#72#));
reg_q276_in <= (reg_q274 AND symb_decoder(16#69#)) OR
 					(reg_q274 AND symb_decoder(16#49#));
reg_q278_in <= (reg_q276 AND symb_decoder(16#50#)) OR
 					(reg_q276 AND symb_decoder(16#70#));
reg_q383_in <= (reg_q381 AND symb_decoder(16#43#)) OR
 					(reg_q381 AND symb_decoder(16#63#));
reg_q385_in <= (reg_q383 AND symb_decoder(16#41#)) OR
 					(reg_q383 AND symb_decoder(16#61#));
reg_q679_in <= (reg_q679 AND symb_decoder(16#32#)) OR
 					(reg_q679 AND symb_decoder(16#35#)) OR
 					(reg_q679 AND symb_decoder(16#36#)) OR
 					(reg_q679 AND symb_decoder(16#31#)) OR
 					(reg_q679 AND symb_decoder(16#30#)) OR
 					(reg_q679 AND symb_decoder(16#33#)) OR
 					(reg_q679 AND symb_decoder(16#34#)) OR
 					(reg_q679 AND symb_decoder(16#37#)) OR
 					(reg_q679 AND symb_decoder(16#38#)) OR
 					(reg_q679 AND symb_decoder(16#39#)) OR
 					(reg_q677 AND symb_decoder(16#33#)) OR
 					(reg_q677 AND symb_decoder(16#38#)) OR
 					(reg_q677 AND symb_decoder(16#37#)) OR
 					(reg_q677 AND symb_decoder(16#30#)) OR
 					(reg_q677 AND symb_decoder(16#36#)) OR
 					(reg_q677 AND symb_decoder(16#32#)) OR
 					(reg_q677 AND symb_decoder(16#34#)) OR
 					(reg_q677 AND symb_decoder(16#35#)) OR
 					(reg_q677 AND symb_decoder(16#39#)) OR
 					(reg_q677 AND symb_decoder(16#31#));
reg_q2284_in <= (reg_q2282 AND symb_decoder(16#65#)) OR
 					(reg_q2282 AND symb_decoder(16#45#));
reg_q1008_in <= (reg_q1006 AND symb_decoder(16#65#)) OR
 					(reg_q1006 AND symb_decoder(16#45#));
reg_q83_in <= (reg_q81 AND symb_decoder(16#6f#)) OR
 					(reg_q81 AND symb_decoder(16#4f#));
reg_q85_in <= (reg_q83 AND symb_decoder(16#52#)) OR
 					(reg_q83 AND symb_decoder(16#72#));
reg_q1181_in <= (reg_q1181 AND symb_decoder(16#0d#)) OR
 					(reg_q1181 AND symb_decoder(16#0a#)) OR
 					(reg_q1181 AND symb_decoder(16#0c#)) OR
 					(reg_q1181 AND symb_decoder(16#09#)) OR
 					(reg_q1181 AND symb_decoder(16#20#)) OR
 					(reg_q1179 AND symb_decoder(16#0d#)) OR
 					(reg_q1179 AND symb_decoder(16#09#)) OR
 					(reg_q1179 AND symb_decoder(16#20#)) OR
 					(reg_q1179 AND symb_decoder(16#0a#)) OR
 					(reg_q1179 AND symb_decoder(16#0c#));
reg_q1345_in <= (reg_q1343 AND symb_decoder(16#0d#)) OR
 					(reg_q1343 AND symb_decoder(16#20#)) OR
 					(reg_q1343 AND symb_decoder(16#0a#)) OR
 					(reg_q1343 AND symb_decoder(16#0c#)) OR
 					(reg_q1343 AND symb_decoder(16#09#)) OR
 					(reg_q1345 AND symb_decoder(16#20#)) OR
 					(reg_q1345 AND symb_decoder(16#0a#)) OR
 					(reg_q1345 AND symb_decoder(16#0c#)) OR
 					(reg_q1345 AND symb_decoder(16#0d#)) OR
 					(reg_q1345 AND symb_decoder(16#09#));
reg_q730_in <= (reg_q728 AND symb_decoder(16#4e#)) OR
 					(reg_q728 AND symb_decoder(16#6e#));
reg_q2341_in <= (reg_q2339 AND symb_decoder(16#49#)) OR
 					(reg_q2339 AND symb_decoder(16#69#));
reg_q2343_in <= (reg_q2341 AND symb_decoder(16#43#)) OR
 					(reg_q2341 AND symb_decoder(16#63#));
reg_q669_in <= (reg_q667 AND symb_decoder(16#41#)) OR
 					(reg_q667 AND symb_decoder(16#61#));
reg_q1518_in <= (reg_q1516 AND symb_decoder(16#2e#));
reg_q1112_in <= (reg_q1110 AND symb_decoder(16#66#)) OR
 					(reg_q1110 AND symb_decoder(16#46#));
reg_q1114_in <= (reg_q1112 AND symb_decoder(16#65#)) OR
 					(reg_q1112 AND symb_decoder(16#45#));
reg_q230_in <= (reg_q228 AND symb_decoder(16#61#)) OR
 					(reg_q228 AND symb_decoder(16#41#));
reg_q1118_in <= (reg_q1116 AND symb_decoder(16#72#)) OR
 					(reg_q1116 AND symb_decoder(16#52#));
reg_q1120_in <= (reg_q1118 AND symb_decoder(16#49#)) OR
 					(reg_q1118 AND symb_decoder(16#69#));
reg_q14_in <= (reg_q11 AND symb_decoder(16#65#)) OR
 					(reg_q11 AND symb_decoder(16#45#));
reg_q16_in <= (reg_q14 AND symb_decoder(16#72#)) OR
 					(reg_q14 AND symb_decoder(16#52#));
reg_q1071_in <= (reg_q1069 AND symb_decoder(16#53#)) OR
 					(reg_q1069 AND symb_decoder(16#73#));
reg_q2256_in <= (reg_q2254 AND symb_decoder(16#72#)) OR
 					(reg_q2254 AND symb_decoder(16#52#));
reg_q2258_in <= (reg_q2256 AND symb_decoder(16#65#)) OR
 					(reg_q2256 AND symb_decoder(16#45#));
reg_q1335_in <= (reg_q1333 AND symb_decoder(16#67#)) OR
 					(reg_q1333 AND symb_decoder(16#47#));
reg_q681_in <= (reg_q679 AND symb_decoder(16#2e#));
reg_q683_in <= (reg_q681 AND symb_decoder(16#31#)) OR
 					(reg_q681 AND symb_decoder(16#39#)) OR
 					(reg_q681 AND symb_decoder(16#34#)) OR
 					(reg_q681 AND symb_decoder(16#38#)) OR
 					(reg_q681 AND symb_decoder(16#32#)) OR
 					(reg_q681 AND symb_decoder(16#35#)) OR
 					(reg_q681 AND symb_decoder(16#33#)) OR
 					(reg_q681 AND symb_decoder(16#30#)) OR
 					(reg_q681 AND symb_decoder(16#36#)) OR
 					(reg_q681 AND symb_decoder(16#37#)) OR
 					(reg_q683 AND symb_decoder(16#35#)) OR
 					(reg_q683 AND symb_decoder(16#32#)) OR
 					(reg_q683 AND symb_decoder(16#39#)) OR
 					(reg_q683 AND symb_decoder(16#37#)) OR
 					(reg_q683 AND symb_decoder(16#30#)) OR
 					(reg_q683 AND symb_decoder(16#38#)) OR
 					(reg_q683 AND symb_decoder(16#33#)) OR
 					(reg_q683 AND symb_decoder(16#31#)) OR
 					(reg_q683 AND symb_decoder(16#36#)) OR
 					(reg_q683 AND symb_decoder(16#34#));
reg_q1984_in <= (reg_q1982 AND symb_decoder(16#45#)) OR
 					(reg_q1982 AND symb_decoder(16#65#));
reg_q1986_in <= (reg_q1984 AND symb_decoder(16#38#));
reg_q26_in <= (reg_q24 AND symb_decoder(16#2d#));
reg_q28_in <= (reg_q26 AND symb_decoder(16#0a#)) OR
 					(reg_q26 AND symb_decoder(16#2a#)) OR
 					(reg_q26 AND symb_decoder(16#0d#));
reg_q22_in <= (reg_q20 AND symb_decoder(16#72#)) OR
 					(reg_q20 AND symb_decoder(16#52#));
reg_q1699_in <= (reg_q1697 AND symb_decoder(16#69#)) OR
 					(reg_q1697 AND symb_decoder(16#49#));
reg_q1175_in <= (reg_q1173 AND symb_decoder(16#49#)) OR
 					(reg_q1173 AND symb_decoder(16#69#));
reg_q1177_in <= (reg_q1175 AND symb_decoder(16#6f#)) OR
 					(reg_q1175 AND symb_decoder(16#4f#));
reg_q381_in <= (reg_q377 AND symb_decoder(16#73#)) OR
 					(reg_q377 AND symb_decoder(16#53#)) OR
 					(reg_q393 AND symb_decoder(16#53#)) OR
 					(reg_q393 AND symb_decoder(16#73#));
reg_q2365_in <= (reg_q2361 AND symb_decoder(16#49#)) OR
 					(reg_q2361 AND symb_decoder(16#69#));
reg_q2367_in <= (reg_q2365 AND symb_decoder(16#4e#)) OR
 					(reg_q2365 AND symb_decoder(16#6e#));
reg_q192_in <= (reg_q190 AND symb_decoder(16#74#)) OR
 					(reg_q190 AND symb_decoder(16#54#));
reg_q194_in <= (reg_q192 AND symb_decoder(16#42#)) OR
 					(reg_q192 AND symb_decoder(16#62#));
reg_q1488_in <= (reg_q1486 AND symb_decoder(16#4e#)) OR
 					(reg_q1486 AND symb_decoder(16#6e#));
reg_q1490_in <= (reg_q1488 AND symb_decoder(16#43#)) OR
 					(reg_q1488 AND symb_decoder(16#63#));
reg_q1758_in <= (reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q1757 AND symb_decoder(16#22#));
reg_q1760_in <= (reg_q1758 AND symb_decoder(16#57#)) OR
 					(reg_q1758 AND symb_decoder(16#77#));
reg_q2331_in <= (reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2330 AND symb_decoder(16#3b#));
reg_q2333_in <= (reg_q2331 AND symb_decoder(16#73#)) OR
 					(reg_q2331 AND symb_decoder(16#53#));
reg_q163_in <= (reg_q161 AND symb_decoder(16#4f#)) OR
 					(reg_q161 AND symb_decoder(16#6f#));
reg_q165_in <= (reg_q163 AND symb_decoder(16#4e#)) OR
 					(reg_q163 AND symb_decoder(16#6e#));
reg_q2252_in <= (reg_q2250 AND symb_decoder(16#4f#)) OR
 					(reg_q2250 AND symb_decoder(16#6f#));
reg_q2254_in <= (reg_q2252 AND symb_decoder(16#2c#));
reg_q1988_in <= (reg_q1986 AND symb_decoder(16#30#));
reg_q553_in <= (reg_q551 AND symb_decoder(16#73#)) OR
 					(reg_q551 AND symb_decoder(16#53#));
reg_q671_in <= (reg_q669 AND symb_decoder(16#44#)) OR
 					(reg_q669 AND symb_decoder(16#64#));
reg_q2716_in <= (reg_q2714 AND symb_decoder(16#6b#)) OR
 					(reg_q2714 AND symb_decoder(16#4b#));
reg_q2690_in <= (reg_q2688 AND symb_decoder(16#74#)) OR
 					(reg_q2688 AND symb_decoder(16#54#));
reg_q2692_in <= (reg_q2690 AND symb_decoder(16#75#)) OR
 					(reg_q2690 AND symb_decoder(16#55#));
reg_q1741_in <= (reg_q1739 AND symb_decoder(16#6c#)) OR
 					(reg_q1739 AND symb_decoder(16#4c#));
reg_q1337_in <= (reg_q1335 AND symb_decoder(16#52#)) OR
 					(reg_q1335 AND symb_decoder(16#72#));
reg_q75_in <= (reg_q73 AND symb_decoder(16#61#)) OR
 					(reg_q73 AND symb_decoder(16#41#));
reg_q24_in <= (reg_q22 AND symb_decoder(16#2a#)) OR
 					(reg_q22 AND symb_decoder(16#0d#)) OR
 					(reg_q22 AND symb_decoder(16#0a#));
reg_q1191_in <= (reg_q1189 AND symb_decoder(16#53#)) OR
 					(reg_q1189 AND symb_decoder(16#73#));
reg_q2603_in <= (reg_q2601 AND symb_decoder(16#64#)) OR
 					(reg_q2601 AND symb_decoder(16#44#));
reg_q2605_in <= (reg_q2603 AND symb_decoder(16#20#));
reg_q1932_in <= (reg_q1932 AND symb_decoder(16#39#)) OR
 					(reg_q1932 AND symb_decoder(16#37#)) OR
 					(reg_q1932 AND symb_decoder(16#35#)) OR
 					(reg_q1932 AND symb_decoder(16#32#)) OR
 					(reg_q1932 AND symb_decoder(16#30#)) OR
 					(reg_q1932 AND symb_decoder(16#36#)) OR
 					(reg_q1932 AND symb_decoder(16#33#)) OR
 					(reg_q1932 AND symb_decoder(16#34#)) OR
 					(reg_q1932 AND symb_decoder(16#38#)) OR
 					(reg_q1932 AND symb_decoder(16#31#)) OR
 					(reg_q1930 AND symb_decoder(16#38#)) OR
 					(reg_q1930 AND symb_decoder(16#37#)) OR
 					(reg_q1930 AND symb_decoder(16#33#)) OR
 					(reg_q1930 AND symb_decoder(16#35#)) OR
 					(reg_q1930 AND symb_decoder(16#39#)) OR
 					(reg_q1930 AND symb_decoder(16#36#)) OR
 					(reg_q1930 AND symb_decoder(16#32#)) OR
 					(reg_q1930 AND symb_decoder(16#30#)) OR
 					(reg_q1930 AND symb_decoder(16#31#)) OR
 					(reg_q1930 AND symb_decoder(16#34#));
reg_q950_in <= (reg_q948 AND symb_decoder(16#49#));
reg_q2710_in <= (reg_q2708 AND symb_decoder(16#20#)) OR
 					(reg_q2708 AND symb_decoder(16#0a#)) OR
 					(reg_q2708 AND symb_decoder(16#0d#)) OR
 					(reg_q2708 AND symb_decoder(16#09#)) OR
 					(reg_q2708 AND symb_decoder(16#0c#));
reg_q36_in <= (reg_q34 AND symb_decoder(16#4e#)) OR
 					(reg_q34 AND symb_decoder(16#6e#));
reg_q1155_in <= (reg_q1153 AND symb_decoder(16#47#)) OR
 					(reg_q1153 AND symb_decoder(16#67#));
reg_q1157_in <= (reg_q1155 AND symb_decoder(16#48#)) OR
 					(reg_q1155 AND symb_decoder(16#68#));
reg_q153_in <= (reg_q151 AND symb_decoder(16#56#)) OR
 					(reg_q151 AND symb_decoder(16#76#));
reg_q1169_in <= (reg_q1167 AND symb_decoder(16#65#)) OR
 					(reg_q1167 AND symb_decoder(16#45#));
reg_q266_in <= (reg_q264 AND symb_decoder(16#79#)) OR
 					(reg_q264 AND symb_decoder(16#59#));
reg_q507_in <= (reg_q505 AND symb_decoder(16#6f#)) OR
 					(reg_q505 AND symb_decoder(16#4f#));
reg_q509_in <= (reg_q507 AND symb_decoder(16#3b#));
reg_q2611_in <= (reg_q2609 AND symb_decoder(16#54#)) OR
 					(reg_q2609 AND symb_decoder(16#74#));
reg_q2613_in <= (reg_q2611 AND symb_decoder(16#68#)) OR
 					(reg_q2611 AND symb_decoder(16#48#));
reg_q2700_in <= (reg_q2698 AND symb_decoder(16#45#)) OR
 					(reg_q2698 AND symb_decoder(16#65#));
reg_q196_in <= (reg_q194 AND symb_decoder(16#0a#)) OR
 					(reg_q194 AND symb_decoder(16#0c#)) OR
 					(reg_q194 AND symb_decoder(16#20#)) OR
 					(reg_q194 AND symb_decoder(16#09#)) OR
 					(reg_q194 AND symb_decoder(16#0d#)) OR
 					(reg_q196 AND symb_decoder(16#09#)) OR
 					(reg_q196 AND symb_decoder(16#0c#)) OR
 					(reg_q196 AND symb_decoder(16#0d#)) OR
 					(reg_q196 AND symb_decoder(16#20#)) OR
 					(reg_q196 AND symb_decoder(16#0a#));
reg_q2708_in <= (reg_q2706 AND symb_decoder(16#52#)) OR
 					(reg_q2706 AND symb_decoder(16#72#));
reg_q561_in <= (reg_q559 AND symb_decoder(16#65#)) OR
 					(reg_q559 AND symb_decoder(16#45#));
reg_q161_in <= (reg_q159 AND symb_decoder(16#69#)) OR
 					(reg_q159 AND symb_decoder(16#49#));
reg_q224_in <= (reg_q222 AND symb_decoder(16#72#)) OR
 					(reg_q222 AND symb_decoder(16#52#));
reg_q232_in <= (reg_q230 AND symb_decoder(16#4c#)) OR
 					(reg_q230 AND symb_decoder(16#6c#));
reg_q234_in <= (reg_q232 AND symb_decoder(16#4c#)) OR
 					(reg_q232 AND symb_decoder(16#6c#));
reg_q2593_in <= (reg_q2591 AND symb_decoder(16#6e#)) OR
 					(reg_q2591 AND symb_decoder(16#4e#));
reg_q2595_in <= (reg_q2593 AND symb_decoder(16#65#)) OR
 					(reg_q2593 AND symb_decoder(16#45#));
reg_q594_in <= (reg_q592 AND symb_decoder(16#70#)) OR
 					(reg_q592 AND symb_decoder(16#50#));
reg_q2698_in <= (reg_q2696 AND symb_decoder(16#73#)) OR
 					(reg_q2696 AND symb_decoder(16#53#));
reg_q67_in <= (reg_q65 AND symb_decoder(16#0d#)) OR
 					(reg_q65 AND symb_decoder(16#2a#)) OR
 					(reg_q65 AND symb_decoder(16#0a#));
reg_q2302_in <= (reg_q2300 AND symb_decoder(16#52#)) OR
 					(reg_q2300 AND symb_decoder(16#72#));
reg_q2351_in <= (reg_q2349 AND symb_decoder(16#74#)) OR
 					(reg_q2349 AND symb_decoder(16#54#));
reg_q2353_in <= (reg_q2351 AND symb_decoder(16#61#)) OR
 					(reg_q2351 AND symb_decoder(16#41#));
reg_q1930_in <= (reg_q1928 AND symb_decoder(16#2a#));
reg_q1695_in <= (reg_q1693 AND symb_decoder(16#50#)) OR
 					(reg_q1693 AND symb_decoder(16#70#));
reg_q1697_in <= (reg_q1695 AND symb_decoder(16#74#)) OR
 					(reg_q1695 AND symb_decoder(16#54#));
reg_q268_in <= (reg_q266 AND symb_decoder(16#6f#)) OR
 					(reg_q266 AND symb_decoder(16#4f#));
reg_q1085_in <= (reg_q1083 AND symb_decoder(16#52#)) OR
 					(reg_q1083 AND symb_decoder(16#72#));
reg_q685_in <= (reg_q683 AND symb_decoder(16#0d#)) OR
 					(reg_q683 AND symb_decoder(16#0c#)) OR
 					(reg_q683 AND symb_decoder(16#09#)) OR
 					(reg_q683 AND symb_decoder(16#20#)) OR
 					(reg_q683 AND symb_decoder(16#0a#));
reg_q1739_in <= (reg_q1737 AND symb_decoder(16#6e#)) OR
 					(reg_q1737 AND symb_decoder(16#4e#));
reg_q2361_in <= (reg_q2359 AND symb_decoder(16#3b#));
reg_q262_in <= (reg_q260 AND symb_decoder(16#2e#));
reg_q46_in <= (reg_q44 AND symb_decoder(16#53#)) OR
 					(reg_q44 AND symb_decoder(16#73#));
reg_q1747_in <= (reg_q1745 AND symb_decoder(16#65#)) OR
 					(reg_q1745 AND symb_decoder(16#45#));
reg_q2371_in <= (reg_q2369 AND symb_decoder(16#43#)) OR
 					(reg_q2369 AND symb_decoder(16#63#));
reg_q2324_in <= (reg_q2324 AND symb_decoder(16#0a#)) OR
 					(reg_q2324 AND symb_decoder(16#09#)) OR
 					(reg_q2324 AND symb_decoder(16#0c#)) OR
 					(reg_q2324 AND symb_decoder(16#20#)) OR
 					(reg_q2324 AND symb_decoder(16#0d#)) OR
 					(reg_q2322 AND symb_decoder(16#20#)) OR
 					(reg_q2322 AND symb_decoder(16#09#)) OR
 					(reg_q2322 AND symb_decoder(16#0c#)) OR
 					(reg_q2322 AND symb_decoder(16#0a#)) OR
 					(reg_q2322 AND symb_decoder(16#0d#));
reg_q1980_in <= (reg_q1978 AND symb_decoder(16#34#));
reg_q2379_in <= (reg_q2377 AND symb_decoder(16#65#)) OR
 					(reg_q2377 AND symb_decoder(16#45#));
reg_q139_in <= (reg_q137 AND symb_decoder(16#73#)) OR
 					(reg_q137 AND symb_decoder(16#53#));
reg_q2377_in <= (reg_q2375 AND symb_decoder(16#76#)) OR
 					(reg_q2375 AND symb_decoder(16#56#));
reg_q93_in <= (reg_q91 AND symb_decoder(16#6b#)) OR
 					(reg_q91 AND symb_decoder(16#4b#));
reg_q95_in <= (reg_q93 AND symb_decoder(16#0d#));
reg_q1798_in <= (reg_q1796 AND symb_decoder(16#72#)) OR
 					(reg_q1796 AND symb_decoder(16#52#));
reg_q2730_in <= (reg_q2728 AND symb_decoder(16#49#)) OR
 					(reg_q2728 AND symb_decoder(16#69#));
reg_q2732_in <= (reg_q2730 AND symb_decoder(16#6e#)) OR
 					(reg_q2730 AND symb_decoder(16#4e#));
reg_q1329_in <= (reg_q1327 AND symb_decoder(16#49#)) OR
 					(reg_q1327 AND symb_decoder(16#69#));
reg_q155_in <= (reg_q153 AND symb_decoder(16#65#)) OR
 					(reg_q153 AND symb_decoder(16#45#));
reg_q157_in <= (reg_q155 AND symb_decoder(16#52#)) OR
 					(reg_q155 AND symb_decoder(16#72#));
reg_q1784_in <= (reg_q1784 AND symb_decoder(16#09#)) OR
 					(reg_q1784 AND symb_decoder(16#20#)) OR
 					(reg_q1784 AND symb_decoder(16#0a#)) OR
 					(reg_q1784 AND symb_decoder(16#0d#)) OR
 					(reg_q1784 AND symb_decoder(16#0c#)) OR
 					(reg_q1782 AND symb_decoder(16#20#)) OR
 					(reg_q1782 AND symb_decoder(16#0d#)) OR
 					(reg_q1782 AND symb_decoder(16#09#)) OR
 					(reg_q1782 AND symb_decoder(16#0a#)) OR
 					(reg_q1782 AND symb_decoder(16#0c#));
reg_q202_in <= (reg_q200 AND symb_decoder(16#36#));
reg_q1002_in <= (reg_q1000 AND symb_decoder(16#46#)) OR
 					(reg_q1000 AND symb_decoder(16#66#));
reg_q2335_in <= (reg_q2333 AND symb_decoder(16#45#)) OR
 					(reg_q2333 AND symb_decoder(16#65#));
reg_q1792_in <= (reg_q1790 AND symb_decoder(16#61#)) OR
 					(reg_q1790 AND symb_decoder(16#41#));
reg_q1134_in <= (reg_q1132 AND symb_decoder(16#45#)) OR
 					(reg_q1132 AND symb_decoder(16#65#));
reg_q677_in <= (reg_q675 AND symb_decoder(16#2e#));
reg_q2734_in <= (reg_q2732 AND symb_decoder(16#67#)) OR
 					(reg_q2732 AND symb_decoder(16#47#));
reg_q2322_in <= (reg_q2320 AND symb_decoder(16#3a#));
reg_q1140_in <= (reg_q1138 AND symb_decoder(16#6f#)) OR
 					(reg_q1138 AND symb_decoder(16#4f#));
reg_q2403_in <= (reg_q2401 AND symb_decoder(16#54#)) OR
 					(reg_q2401 AND symb_decoder(16#74#));
reg_q2405_in <= (reg_q2403 AND symb_decoder(16#69#)) OR
 					(reg_q2403 AND symb_decoder(16#49#));
reg_q2320_in <= (reg_q2318 AND symb_decoder(16#72#)) OR
 					(reg_q2318 AND symb_decoder(16#52#));
reg_q1153_in <= (reg_q1151 AND symb_decoder(16#3a#));
reg_q505_in <= (reg_q503 AND symb_decoder(16#46#)) OR
 					(reg_q503 AND symb_decoder(16#66#));
reg_q1687_in <= (reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q1686 AND symb_decoder(16#21#));
reg_q65_in <= (reg_q63 AND symb_decoder(16#6b#)) OR
 					(reg_q63 AND symb_decoder(16#4b#));
reg_q56_in <= (reg_q54 AND symb_decoder(16#44#)) OR
 					(reg_q54 AND symb_decoder(16#64#));
reg_q687_in <= (reg_q685 AND symb_decoder(16#0d#)) OR
 					(reg_q685 AND symb_decoder(16#09#)) OR
 					(reg_q685 AND symb_decoder(16#20#)) OR
 					(reg_q685 AND symb_decoder(16#0a#)) OR
 					(reg_q685 AND symb_decoder(16#0c#));
reg_q365_in <= (reg_q363 AND symb_decoder(16#6f#)) OR
 					(reg_q363 AND symb_decoder(16#4f#));
reg_q367_in <= (reg_q365 AND symb_decoder(16#4f#)) OR
 					(reg_q365 AND symb_decoder(16#6f#));
reg_q2260_in <= (reg_q2258 AND symb_decoder(16#67#)) OR
 					(reg_q2258 AND symb_decoder(16#47#));
reg_q2262_in <= (reg_q2260 AND symb_decoder(16#69#)) OR
 					(reg_q2260 AND symb_decoder(16#49#));
reg_q363_in <= (reg_q359 AND symb_decoder(16#52#)) OR
 					(reg_q359 AND symb_decoder(16#72#)) OR
 					(reg_q397 AND symb_decoder(16#72#)) OR
 					(reg_q397 AND symb_decoder(16#52#));
reg_q1104_in <= (reg_q1102 AND symb_decoder(16#52#)) OR
 					(reg_q1102 AND symb_decoder(16#72#));
reg_q1106_in <= (reg_q1104 AND symb_decoder(16#61#)) OR
 					(reg_q1104 AND symb_decoder(16#41#));
reg_q728_in <= (reg_q726 AND symb_decoder(16#61#)) OR
 					(reg_q726 AND symb_decoder(16#41#));
reg_q957_in <= (reg_q955 AND symb_decoder(16#49#));
reg_q1506_in <= (reg_q1504 AND symb_decoder(16#52#)) OR
 					(reg_q1504 AND symb_decoder(16#72#));
reg_q137_in <= (reg_q135 AND symb_decoder(16#5f#));
reg_q2337_in <= (reg_q2335 AND symb_decoder(16#52#)) OR
 					(reg_q2335 AND symb_decoder(16#72#));
reg_q2339_in <= (reg_q2337 AND symb_decoder(16#76#)) OR
 					(reg_q2337 AND symb_decoder(16#56#));
reg_q986_in <= (reg_q984 AND symb_decoder(16#46#)) OR
 					(reg_q984 AND symb_decoder(16#66#));
reg_q738_in <= (reg_q736 AND symb_decoder(16#52#)) OR
 					(reg_q736 AND symb_decoder(16#72#));
reg_q1116_in <= (reg_q1114 AND symb_decoder(16#72#)) OR
 					(reg_q1114 AND symb_decoder(16#52#));
reg_q91_in <= (reg_q89 AND symb_decoder(16#4f#)) OR
 					(reg_q89 AND symb_decoder(16#6f#));
reg_q1179_in <= (reg_q1177 AND symb_decoder(16#4e#)) OR
 					(reg_q1177 AND symb_decoder(16#6e#));
reg_q1693_in <= (reg_q1691 AND symb_decoder(16#6f#)) OR
 					(reg_q1691 AND symb_decoder(16#4f#));
reg_q2391_in <= (reg_q2389 AND symb_decoder(16#49#)) OR
 					(reg_q2389 AND symb_decoder(16#69#));
reg_q2607_in <= (reg_q2605 AND symb_decoder(16#57#)) OR
 					(reg_q2605 AND symb_decoder(16#77#));
reg_q2609_in <= (reg_q2607 AND symb_decoder(16#69#)) OR
 					(reg_q2607 AND symb_decoder(16#49#));
reg_q1087_in <= (reg_q1085 AND symb_decoder(16#4f#)) OR
 					(reg_q1085 AND symb_decoder(16#6f#));
reg_q1786_in <= (reg_q1784 AND symb_decoder(16#6d#)) OR
 					(reg_q1784 AND symb_decoder(16#4d#));
reg_q1788_in <= (reg_q1786 AND symb_decoder(16#61#)) OR
 					(reg_q1786 AND symb_decoder(16#41#));
reg_q1016_in <= (reg_q1014 AND symb_decoder(16#6f#)) OR
 					(reg_q1014 AND symb_decoder(16#4f#));
reg_q706_in <= (reg_q704 AND symb_decoder(16#47#)) OR
 					(reg_q704 AND symb_decoder(16#67#));
reg_q2355_in <= (reg_q2353 AND symb_decoder(16#74#)) OR
 					(reg_q2353 AND symb_decoder(16#54#));
reg_q2688_in <= (reg_q2686 AND symb_decoder(16#41#)) OR
 					(reg_q2686 AND symb_decoder(16#61#));
reg_q222_in <= (reg_q220 AND symb_decoder(16#49#)) OR
 					(reg_q220 AND symb_decoder(16#69#));
reg_q248_in <= (reg_q246 AND symb_decoder(16#65#)) OR
 					(reg_q246 AND symb_decoder(16#45#));
reg_q1353_in <= (reg_q1351 AND symb_decoder(16#6d#)) OR
 					(reg_q1351 AND symb_decoder(16#4d#));
reg_q63_in <= (reg_q11 AND symb_decoder(16#4f#)) OR
 					(reg_q11 AND symb_decoder(16#6f#));
reg_q984_in <= (reg_q982 AND symb_decoder(16#73#)) OR
 					(reg_q982 AND symb_decoder(16#53#));
reg_q2748_in <= (reg_q2746 AND symb_decoder(16#65#)) OR
 					(reg_q2746 AND symb_decoder(16#45#));
reg_q1018_in <= (reg_q1016 AND symb_decoder(16#4d#)) OR
 					(reg_q1016 AND symb_decoder(16#6d#));
reg_q2411_in <= (reg_q2361 AND symb_decoder(16#61#)) OR
 					(reg_q2361 AND symb_decoder(16#41#));
reg_q2589_in <= (reg_q2587 AND symb_decoder(16#4f#)) OR
 					(reg_q2587 AND symb_decoder(16#6f#));
reg_q2591_in <= (reg_q2589 AND symb_decoder(16#4e#)) OR
 					(reg_q2589 AND symb_decoder(16#6e#));
reg_q1982_in <= (reg_q1980 AND symb_decoder(16#30#));
reg_q2401_in <= (reg_q2399 AND symb_decoder(16#43#)) OR
 					(reg_q2399 AND symb_decoder(16#63#));
reg_q1319_in <= (reg_q1317 AND symb_decoder(16#6f#)) OR
 					(reg_q1317 AND symb_decoder(16#4f#));
reg_q726_in <= (reg_q724 AND symb_decoder(16#4a#)) OR
 					(reg_q724 AND symb_decoder(16#6a#));
reg_q1108_in <= (reg_q1106 AND symb_decoder(16#4e#)) OR
 					(reg_q1106 AND symb_decoder(16#6e#));
reg_q1110_in <= (reg_q1108 AND symb_decoder(16#53#)) OR
 					(reg_q1108 AND symb_decoder(16#73#));
reg_q1355_in <= (reg_q1353 AND symb_decoder(16#4f#)) OR
 					(reg_q1353 AND symb_decoder(16#6f#));
reg_q704_in <= (reg_q702 AND symb_decoder(16#56#)) OR
 					(reg_q702 AND symb_decoder(16#76#));
reg_q1122_in <= (reg_q1120 AND symb_decoder(16#4e#)) OR
 					(reg_q1120 AND symb_decoder(16#6e#));
reg_q1749_in <= (reg_q1747 AND symb_decoder(16#21#));
reg_q159_in <= (reg_q157 AND symb_decoder(16#73#)) OR
 					(reg_q157 AND symb_decoder(16#53#));
reg_q2587_in <= (reg_q2585 AND symb_decoder(16#63#)) OR
 					(reg_q2585 AND symb_decoder(16#43#));
reg_q2345_in <= (reg_q2343 AND symb_decoder(16#45#)) OR
 					(reg_q2343 AND symb_decoder(16#65#));
reg_q2750_in <= (reg_q2748 AND symb_decoder(16#64#)) OR
 					(reg_q2748 AND symb_decoder(16#44#));
reg_q1937_in <= (reg_q1935 AND symb_decoder(16#50#));
reg_q1705_in <= (reg_q1703 AND symb_decoder(16#50#)) OR
 					(reg_q1703 AND symb_decoder(16#70#));
reg_q748_in <= (reg_q746 AND symb_decoder(16#32#));
reg_q2369_in <= (reg_q2367 AND symb_decoder(16#61#)) OR
 					(reg_q2367 AND symb_decoder(16#41#));
reg_q596_in <= (reg_q594 AND symb_decoder(16#61#)) OR
 					(reg_q594 AND symb_decoder(16#41#));
reg_q598_in <= (reg_q596 AND symb_decoder(16#73#)) OR
 					(reg_q596 AND symb_decoder(16#53#));
reg_q1321_in <= (reg_q1319 AND symb_decoder(16#74#)) OR
 					(reg_q1319 AND symb_decoder(16#54#));
reg_q2318_in <= (reg_q2316 AND symb_decoder(16#65#)) OR
 					(reg_q2316 AND symb_decoder(16#45#));
reg_q976_in <= (reg_q974 AND symb_decoder(16#54#)) OR
 					(reg_q974 AND symb_decoder(16#74#));
reg_q1782_in <= (reg_q1780 AND symb_decoder(16#65#)) OR
 					(reg_q1780 AND symb_decoder(16#45#));
reg_q7_in <= (reg_q5 AND symb_decoder(16#73#)) OR
 					(reg_q5 AND symb_decoder(16#53#));
reg_q2248_in <= (reg_q2246 AND symb_decoder(16#6e#)) OR
 					(reg_q2246 AND symb_decoder(16#4e#));
reg_q103_in <= (reg_q101 AND symb_decoder(16#57#)) OR
 					(reg_q101 AND symb_decoder(16#77#));
reg_q513_in <= (reg_q511 AND symb_decoder(16#3b#));
reg_q980_in <= (reg_q978 AND symb_decoder(16#61#)) OR
 					(reg_q978 AND symb_decoder(16#41#));
reg_q982_in <= (reg_q980 AND symb_decoder(16#4e#)) OR
 					(reg_q980 AND symb_decoder(16#6e#));
reg_q246_in <= (reg_q244 AND symb_decoder(16#44#)) OR
 					(reg_q244 AND symb_decoder(16#64#));
reg_q965_in <= (reg_q963 AND symb_decoder(16#59#));
reg_q1508_in <= (reg_q1506 AND symb_decoder(16#56#)) OR
 					(reg_q1506 AND symb_decoder(16#76#));
reg_q1067_in <= (reg_q1065 AND symb_decoder(16#65#)) OR
 					(reg_q1065 AND symb_decoder(16#45#));
reg_q48_in <= (reg_q46 AND symb_decoder(16#53#)) OR
 					(reg_q46 AND symb_decoder(16#73#));
reg_q1347_in <= (reg_q1345 AND symb_decoder(16#44#)) OR
 					(reg_q1345 AND symb_decoder(16#64#));
reg_q1091_in <= (reg_q1089 AND symb_decoder(16#41#)) OR
 					(reg_q1089 AND symb_decoder(16#61#));
reg_q1093_in <= (reg_q1091 AND symb_decoder(16#6e#)) OR
 					(reg_q1091 AND symb_decoder(16#4e#));
reg_q1751_in <= (reg_q1749 AND symb_decoder(16#21#));
reg_q1790_in <= (reg_q1788 AND symb_decoder(16#4e#)) OR
 					(reg_q1788 AND symb_decoder(16#6e#));
reg_q750_in <= (reg_q748 AND symb_decoder(16#30#));
reg_q1492_in <= (reg_q1490 AND symb_decoder(16#72#)) OR
 					(reg_q1490 AND symb_decoder(16#52#));
reg_q1928_in <= (reg_q1926 AND symb_decoder(16#32#));
reg_q1089_in <= (reg_q1087 AND symb_decoder(16#4a#)) OR
 					(reg_q1087 AND symb_decoder(16#6a#));
reg_q1197_in <= (reg_q1195 AND symb_decoder(16#76#)) OR
 					(reg_q1195 AND symb_decoder(16#56#));
reg_q600_in <= (reg_q598 AND symb_decoder(16#32#)) OR
 					(reg_q598 AND symb_decoder(16#33#));
reg_q602_in <= (reg_q600 AND symb_decoder(16#3a#));
reg_q536_in <= (reg_q534 AND symb_decoder(16#0d#));
reg_q538_in <= (reg_q536 AND symb_decoder(16#0a#));
reg_q2250_in <= (reg_q2248 AND symb_decoder(16#46#)) OR
 					(reg_q2248 AND symb_decoder(16#66#));
reg_q73_in <= (reg_q71 AND symb_decoder(16#70#)) OR
 					(reg_q71 AND symb_decoder(16#50#));
reg_q978_in <= (reg_q976 AND symb_decoder(16#72#)) OR
 					(reg_q976 AND symb_decoder(16#52#));
reg_q256_in <= (reg_q254 AND symb_decoder(16#6f#)) OR
 					(reg_q254 AND symb_decoder(16#4f#));
reg_q128_in <= (reg_q126 AND symb_decoder(16#3a#));
reg_q130_in <= (reg_q128 AND symb_decoder(16#5c#));
reg_q959_in <= (reg_q957 AND symb_decoder(16#52#));
reg_q960_in <= (reg_q959 AND symb_decoder(16#0d#));
reg_q2413_in <= (reg_q2411 AND symb_decoder(16#4c#)) OR
 					(reg_q2411 AND symb_decoder(16#6c#));
reg_q752_in <= (reg_q750 AND symb_decoder(16#30#));
reg_q1216_in <= (reg_q1214 AND symb_decoder(16#3b#));
reg_q198_in <= (reg_q196 AND symb_decoder(16#36#));
reg_q1142_in <= (reg_q1140 AND symb_decoder(16#3a#));
reg_q2755_in <= (reg_q2754 AND symb_decoder(16#0d#));
reg_q689_in <= (reg_q687 AND symb_decoder(16#3e#));
reg_q97_in <= (reg_q95 AND symb_decoder(16#0a#));
reg_q754_in <= (reg_q752 AND symb_decoder(16#30#));
reg_q1753_in <= (reg_q1751 AND symb_decoder(16#21#));
reg_q691_in <= (reg_q689 AND symb_decoder(16#3c#));
reg_q200_in <= (reg_q198 AND symb_decoder(16#36#));
reg_q1020_in <= (reg_q1018 AND symb_decoder(16#3a#));
reg_fullgraph1_init <= "0000000000";

reg_fullgraph1_sel <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & reg_q1020_in & reg_q200_in & reg_q691_in & reg_q1753_in & reg_q754_in & reg_q97_in & reg_q689_in & reg_q2755_in & reg_q1142_in & reg_q198_in & reg_q1216_in & reg_q752_in & reg_q2413_in & reg_q960_in & reg_q959_in & reg_q130_in & reg_q128_in & reg_q256_in & reg_q978_in & reg_q73_in & reg_q2250_in & reg_q538_in & reg_q536_in & reg_q602_in & reg_q600_in & reg_q1197_in & reg_q1089_in & reg_q1928_in & reg_q1492_in & reg_q750_in & reg_q1790_in & reg_q1751_in & reg_q1093_in & reg_q1091_in & reg_q1347_in & reg_q48_in & reg_q1067_in & reg_q1508_in & reg_q965_in & reg_q246_in & reg_q982_in & reg_q980_in & reg_q513_in & reg_q103_in & reg_q2248_in & reg_q7_in & reg_q1782_in & reg_q976_in & reg_q2318_in & reg_q1321_in & reg_q598_in & reg_q596_in & reg_q2369_in & reg_q748_in & reg_q1705_in & reg_q1937_in & reg_q2750_in & reg_q2345_in & reg_q2587_in & reg_q159_in & reg_q1749_in & reg_q1122_in & reg_q704_in & reg_q1355_in & reg_q1110_in & reg_q1108_in & reg_q726_in & reg_q1319_in & reg_q2401_in & reg_q1982_in & reg_q2591_in & reg_q2589_in & reg_q2411_in & reg_q1018_in & reg_q2748_in & reg_q984_in & reg_q63_in & reg_q1353_in & reg_q248_in & reg_q222_in & reg_q2688_in & reg_q2355_in & reg_q706_in & reg_q1016_in & reg_q1788_in & reg_q1786_in & reg_q1087_in & reg_q2609_in & reg_q2607_in & reg_q2391_in & reg_q1693_in & reg_q1179_in & reg_q91_in & reg_q1116_in & reg_q738_in & reg_q986_in & reg_q2339_in & reg_q2337_in & reg_q137_in & reg_q1506_in & reg_q957_in & reg_q728_in & reg_q1106_in & reg_q1104_in & reg_q363_in & reg_q2262_in & reg_q2260_in & reg_q367_in & reg_q365_in & reg_q687_in & reg_q56_in & reg_q65_in & reg_q1687_in & reg_q505_in & reg_q1153_in & reg_q2320_in & reg_q2405_in & reg_q2403_in & reg_q1140_in & reg_q2322_in & reg_q2734_in & reg_q677_in & reg_q1134_in & reg_q1792_in & reg_q2335_in & reg_q1002_in & reg_q202_in & reg_q1784_in & reg_q157_in & reg_q155_in & reg_q1329_in & reg_q2732_in & reg_q2730_in & reg_q1798_in & reg_q95_in & reg_q93_in & reg_q2377_in & reg_q139_in & reg_q2379_in & reg_q1980_in & reg_q2324_in & reg_q2371_in & reg_q1747_in & reg_q46_in & reg_q262_in & reg_q2361_in & reg_q1739_in & reg_q685_in & reg_q1085_in & reg_q268_in & reg_q1697_in & reg_q1695_in & reg_q1930_in & reg_q2353_in & reg_q2351_in & reg_q2302_in & reg_q67_in & reg_q2698_in & reg_q594_in & reg_q2595_in & reg_q2593_in & reg_q234_in & reg_q232_in & reg_q224_in & reg_q161_in & reg_q561_in & reg_q2708_in & reg_q196_in & reg_q2700_in & reg_q2613_in & reg_q2611_in & reg_q509_in & reg_q507_in & reg_q266_in & reg_q1169_in & reg_q153_in & reg_q1157_in & reg_q1155_in & reg_q36_in & reg_q2710_in & reg_q950_in & reg_q1932_in & reg_q2605_in & reg_q2603_in & reg_q1191_in & reg_q24_in & reg_q75_in & reg_q1337_in & reg_q1741_in & reg_q2692_in & reg_q2690_in & reg_q2716_in & reg_q671_in & reg_q553_in & reg_q1988_in & reg_q2254_in & reg_q2252_in & reg_q165_in & reg_q163_in & reg_q2333_in & reg_q2331_in & reg_q1760_in & reg_q1758_in & reg_q1490_in & reg_q1488_in & reg_q194_in & reg_q192_in & reg_q2367_in & reg_q2365_in & reg_q381_in & reg_q1177_in & reg_q1175_in & reg_q1699_in & reg_q22_in & reg_q28_in & reg_q26_in & reg_q1986_in & reg_q1984_in & reg_q683_in & reg_q681_in & reg_q1335_in & reg_q2258_in & reg_q2256_in & reg_q1071_in & reg_q16_in & reg_q14_in & reg_q1120_in & reg_q1118_in & reg_q230_in & reg_q1114_in & reg_q1112_in & reg_q1518_in & reg_q669_in & reg_q2343_in & reg_q2341_in & reg_q730_in & reg_q1345_in & reg_q1181_in & reg_q85_in & reg_q83_in & reg_q1008_in & reg_q2284_in & reg_q679_in & reg_q385_in & reg_q383_in & reg_q278_in & reg_q276_in & reg_q2702_in & reg_q2375_in & reg_q2373_in & reg_q264_in & reg_q2286_in & reg_q1776_in & reg_q2724_in & reg_q2722_in & reg_q2522_in & reg_q1729_in & reg_q1343_in & reg_q389_in & reg_q387_in & reg_q2349_in & reg_q2347_in & reg_q280_in & reg_q1796_in & reg_q1794_in & reg_q274_in & reg_q1069_in & reg_q1000_in & reg_q1814_in & reg_q1812_in & reg_q1163_in & reg_q1905_in & reg_q2300_in & reg_q2298_in & reg_q2270_in & reg_q2268_in & reg_q1079_in & reg_q1077_in & reg_q1006_in & reg_q1004_in & reg_q736_in & reg_q734_in & reg_q272_in & reg_q270_in & reg_q955_in & reg_q967_in & reg_q534_in & reg_q532_in & reg_q1496_in & reg_q1494_in & reg_q1351_in & reg_q1349_in & reg_q673_in & reg_q38_in & reg_q1317_in & reg_q1124_in & reg_q1341_in & reg_q1339_in & reg_q228_in & reg_q226_in & reg_q2359_in & reg_q2357_in & reg_q1185_in & reg_q710_in & reg_q708_in & reg_q2002_in & reg_q994_in & reg_q563_in & reg_q740_in & reg_q1516_in & reg_q1514_in & reg_q2615_in & reg_q1691_in & reg_q1689_in & reg_q988_in & reg_q1081_in & reg_q702_in & reg_q2308_in & reg_q1132_in & reg_q1313_in & reg_q254_in & reg_q1210_in & reg_q1208_in & reg_q1167_in & reg_q1165_in & reg_q5_in & reg_q89_in & reg_q87_in & reg_q746_in & reg_q2686_in & reg_q2684_in & reg_q868_in & reg_q1764_in & reg_q1762_in & reg_q2393_in & reg_q206_in & reg_q204_in & reg_q1745_in & reg_q1743_in & reg_q1727_in & reg_q1725_in & reg_q1810_in & reg_q1808_in & reg_q998_in & reg_q996_in & reg_q2682_in & reg_q2585_in & reg_q2010_in & reg_q2415_in & reg_q252_in & reg_q250_in & reg_q1484_in & reg_q105_in & reg_q2048_in & reg_q551_in & reg_q1327_in & reg_q216_in & reg_q2720_in & reg_q2718_in & reg_q2409_in & reg_q2407_in & reg_q1195_in & reg_q1193_in & reg_q1014_in & reg_q1012_in & reg_q2310_in & reg_q2696_in & reg_q2694_in & reg_q77_in & reg_q2601_in & reg_q2397_in & reg_q2395_in & reg_q375_in & reg_q373_in & reg_q1713_in & reg_q1333_in & reg_q1331_in & reg_q1737_in & reg_q1735_in & reg_q11_in & reg_q9_in & reg_q20_in & reg_q18_in & reg_q992_in & reg_q990_in & reg_q34_in & reg_q32_in & reg_q530_in & reg_q1715_in & reg_q1766_in & reg_q1918_in & reg_q1161_in & reg_q1159_in & reg_q2026_in & reg_q2024_in & reg_q190_in & reg_q1913_in & reg_q1911_in & reg_q244_in & reg_q242_in & reg_q81_in & reg_q79_in & reg_q147_in & reg_q1520_in & reg_q1173_in & reg_q1171_in & reg_q2223_in & reg_q2306_in & reg_q2304_in & reg_q169_in & reg_q167_in & reg_q555_in & reg_q1010_in & reg_q511_in & reg_q1723_in & reg_q145_in & reg_q1802_in & reg_q1800_in & reg_q236_in & reg_q260_in & reg_q258_in & reg_q2046_in & reg_q2044_in & reg_q1075_in & reg_q1073_in & reg_q724_in & reg_q722_in & reg_q1102_in & reg_q1100_in & reg_q2016_in & reg_q1721_in & reg_q171_in & reg_q71_in & reg_q69_in & reg_q1136_in & reg_q2266_in & reg_q2264_in & reg_q1780_in & reg_q1778_in & reg_q2278_in & reg_q2276_in & reg_q212_in & reg_q2004_in & reg_q2619_in & reg_q478_in & reg_q559_in & reg_q557_in & reg_q50_in & reg_q2227_in & reg_q2225_in & reg_q1717_in & reg_q2000_in & reg_q2288_in & reg_q1770_in & reg_q1768_in & reg_q143_in & reg_q141_in & reg_q2599_in & reg_q2597_in & reg_q1189_in & reg_q1187_in & reg_q716_in & reg_q240_in & reg_q238_in & reg_q2621_in & reg_q54_in & reg_q52_in & reg_q1949_in & reg_q1707_in & reg_q501_in & reg_q784_in & reg_q782_in & reg_q2385_in & reg_q2383_in & reg_q2014_in & reg_q2012_in & reg_q974_in & reg_q972_in & reg_q718_in & reg_q1183_in & reg_q60_in & reg_q58_in & reg_q778_in & reg_q776_in & reg_q357_in & reg_q355_in & reg_q2018_in & reg_q2316_in & reg_q1214_in & reg_q1212_in & reg_q1126_in & reg_q208_in & reg_q2042_in & reg_q2040_in & reg_q2728_in & reg_q2726_in & reg_q122_in & reg_q120_in & reg_q1703_in & reg_q1701_in & reg_q2754_in & reg_q2752_in & reg_q768_in & reg_q2617_in & reg_q700_in & reg_q698_in & reg_q1806_in & reg_q1804_in & reg_q1994_in & reg_q2706_in & reg_q2704_in & reg_q1315_in & reg_q2030_in & reg_q2028_in & reg_q44_in & reg_q42_in & reg_q2274_in & reg_q2272_in & reg_q126_in & reg_q124_in & reg_q1947_in & reg_q1945_in & reg_q2032_in & reg_q2714_in & reg_q2712_in & reg_q214_in & reg_q2022_in & reg_q2020_in & reg_q1992_in & reg_q1990_in & reg_q220_in & reg_q218_in & reg_q1498_in & reg_q1915_in & reg_q2746_in & reg_q2744_in & reg_q1500_in & reg_q2389_in & reg_q2387_in & reg_q284_in & reg_q282_in & reg_q2282_in & reg_q2280_in & reg_q1711_in & reg_q1709_in & reg_q1926_in & reg_q1924_in & reg_q714_in & reg_q712_in & reg_q369_in & reg_q210_in & reg_q2054_in & reg_q2050_in & reg_q1130_in & reg_q1128_in & reg_q817_in & reg_q2008_in & reg_q2006_in & reg_q1998_in & reg_q1996_in & reg_q1504_in & reg_q1502_in & reg_q2038_in & reg_q2314_in & reg_q2312_in & reg_q2290_in & reg_q107_in & reg_q1357_in & reg_q732_in & reg_q40_in & reg_q480_in & reg_q151_in & reg_q149_in & reg_q675_in & reg_q2623_in & reg_q2036_in & reg_q2034_in & reg_q359_in & reg_q2524_in & reg_q942_in & reg_q876_in & reg_q2738_in & reg_q2736_in & reg_q1719_in & reg_q522_in & reg_q185_in & reg_q377_in & reg_q2526_in & reg_q494_in & reg_q1323_in & reg_q587_in & reg_q565_in;

	--coder fullgraph1
with reg_fullgraph1_sel select
reg_fullgraph1_in <=
	"0000000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001",
	"0000000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010",
	"0000000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100",
	"0000000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000",
	"0000000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000",
	"0000000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000",
	"0000000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000",
	"0000001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000",
	"0000001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
	"0000001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000",
	"0000001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000",
	"0000001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000",
	"0000001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000",
	"0000001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000",
	"0000001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000",
	"0000010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000",
	"0000010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000",
	"0000010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000",
	"0000010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000",
	"0000010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000",
	"0000010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000",
	"0000010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000",
	"0000010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000",
	"0000011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000",
	"0000011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000",
	"0000011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000",
	"0000011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000",
	"0000011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000",
	"0000011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000",
	"0000011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000",
	"0000011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000",
	"0000100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000",
	"0000100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000",
	"0000100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000",
	"0000100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000",
	"0000100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000",
	"0000100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000",
	"0000100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000",
	"0000100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000",
	"0000101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000",
	"0000101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000",
	"0000101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000",
	"0000101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000",
	"0000101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000",
	"0000101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"0000101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000",
	"0000101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000",
	"0000110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000",
	"0000110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000",
	"0000110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000",
	"0000110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000",
	"0000110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000",
	"0000110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000",
	"0000110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000",
	"0000110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000",
	"0000111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000",
	"0000111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000",
	"0000111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000",
	"0000111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000",
	"0000111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000",
	"0000111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000",
	"0000111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000",
	"0000111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000",
	"0001000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000",
	"0001000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000",
	"0001000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000",
	"0001000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000",
	"0001000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000",
	"0001000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000",
	"0001000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000",
	"0001000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0000000000" when others;
 --end coder

	p_reg_fullgraph1: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph1 <= reg_fullgraph1_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph1 <= reg_fullgraph1_init;
        else
          reg_fullgraph1 <= reg_fullgraph1_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph1

		reg_q565 <= '1' when reg_fullgraph1 = "0000000001" else '0'; 
		reg_q587 <= '1' when reg_fullgraph1 = "0000000010" else '0'; 
		reg_q1323 <= '1' when reg_fullgraph1 = "0000000011" else '0'; 
		reg_q494 <= '1' when reg_fullgraph1 = "0000000100" else '0'; 
		reg_q2526 <= '1' when reg_fullgraph1 = "0000000101" else '0'; 
		reg_q377 <= '1' when reg_fullgraph1 = "0000000110" else '0'; 
		reg_q185 <= '1' when reg_fullgraph1 = "0000000111" else '0'; 
		reg_q522 <= '1' when reg_fullgraph1 = "0000001000" else '0'; 
		reg_q1719 <= '1' when reg_fullgraph1 = "0000001001" else '0'; 
		reg_q2736 <= '1' when reg_fullgraph1 = "0000001010" else '0'; 
		reg_q2738 <= '1' when reg_fullgraph1 = "0000001011" else '0'; 
		reg_q876 <= '1' when reg_fullgraph1 = "0000001100" else '0'; 
		reg_q942 <= '1' when reg_fullgraph1 = "0000001101" else '0'; 
		reg_q2524 <= '1' when reg_fullgraph1 = "0000001110" else '0'; 
		reg_q359 <= '1' when reg_fullgraph1 = "0000001111" else '0'; 
		reg_q2034 <= '1' when reg_fullgraph1 = "0000010000" else '0'; 
		reg_q2036 <= '1' when reg_fullgraph1 = "0000010001" else '0'; 
		reg_q2623 <= '1' when reg_fullgraph1 = "0000010010" else '0'; 
		reg_q675 <= '1' when reg_fullgraph1 = "0000010011" else '0'; 
		reg_q149 <= '1' when reg_fullgraph1 = "0000010100" else '0'; 
		reg_q151 <= '1' when reg_fullgraph1 = "0000010101" else '0'; 
		reg_q480 <= '1' when reg_fullgraph1 = "0000010110" else '0'; 
		reg_q40 <= '1' when reg_fullgraph1 = "0000010111" else '0'; 
		reg_q732 <= '1' when reg_fullgraph1 = "0000011000" else '0'; 
		reg_q1357 <= '1' when reg_fullgraph1 = "0000011001" else '0'; 
		reg_q107 <= '1' when reg_fullgraph1 = "0000011010" else '0'; 
		reg_q2290 <= '1' when reg_fullgraph1 = "0000011011" else '0'; 
		reg_q2312 <= '1' when reg_fullgraph1 = "0000011100" else '0'; 
		reg_q2314 <= '1' when reg_fullgraph1 = "0000011101" else '0'; 
		reg_q2038 <= '1' when reg_fullgraph1 = "0000011110" else '0'; 
		reg_q1502 <= '1' when reg_fullgraph1 = "0000011111" else '0'; 
		reg_q1504 <= '1' when reg_fullgraph1 = "0000100000" else '0'; 
		reg_q1996 <= '1' when reg_fullgraph1 = "0000100001" else '0'; 
		reg_q1998 <= '1' when reg_fullgraph1 = "0000100010" else '0'; 
		reg_q2006 <= '1' when reg_fullgraph1 = "0000100011" else '0'; 
		reg_q2008 <= '1' when reg_fullgraph1 = "0000100100" else '0'; 
		reg_q817 <= '1' when reg_fullgraph1 = "0000100101" else '0'; 
		reg_q1128 <= '1' when reg_fullgraph1 = "0000100110" else '0'; 
		reg_q1130 <= '1' when reg_fullgraph1 = "0000100111" else '0'; 
		reg_q2050 <= '1' when reg_fullgraph1 = "0000101000" else '0'; 
		reg_q2054 <= '1' when reg_fullgraph1 = "0000101001" else '0'; 
		reg_q210 <= '1' when reg_fullgraph1 = "0000101010" else '0'; 
		reg_q369 <= '1' when reg_fullgraph1 = "0000101011" else '0'; 
		reg_q712 <= '1' when reg_fullgraph1 = "0000101100" else '0'; 
		reg_q714 <= '1' when reg_fullgraph1 = "0000101101" else '0'; 
		reg_q1924 <= '1' when reg_fullgraph1 = "0000101110" else '0'; 
		reg_q1926 <= '1' when reg_fullgraph1 = "0000101111" else '0'; 
		reg_q1709 <= '1' when reg_fullgraph1 = "0000110000" else '0'; 
		reg_q1711 <= '1' when reg_fullgraph1 = "0000110001" else '0'; 
		reg_q2280 <= '1' when reg_fullgraph1 = "0000110010" else '0'; 
		reg_q2282 <= '1' when reg_fullgraph1 = "0000110011" else '0'; 
		reg_q282 <= '1' when reg_fullgraph1 = "0000110100" else '0'; 
		reg_q284 <= '1' when reg_fullgraph1 = "0000110101" else '0'; 
		reg_q2387 <= '1' when reg_fullgraph1 = "0000110110" else '0'; 
		reg_q2389 <= '1' when reg_fullgraph1 = "0000110111" else '0'; 
		reg_q1500 <= '1' when reg_fullgraph1 = "0000111000" else '0'; 
		reg_q2744 <= '1' when reg_fullgraph1 = "0000111001" else '0'; 
		reg_q2746 <= '1' when reg_fullgraph1 = "0000111010" else '0'; 
		reg_q1915 <= '1' when reg_fullgraph1 = "0000111011" else '0'; 
		reg_q1498 <= '1' when reg_fullgraph1 = "0000111100" else '0'; 
		reg_q218 <= '1' when reg_fullgraph1 = "0000111101" else '0'; 
		reg_q220 <= '1' when reg_fullgraph1 = "0000111110" else '0'; 
		reg_q1990 <= '1' when reg_fullgraph1 = "0000111111" else '0'; 
		reg_q1992 <= '1' when reg_fullgraph1 = "0001000000" else '0'; 
		reg_q2020 <= '1' when reg_fullgraph1 = "0001000001" else '0'; 
		reg_q2022 <= '1' when reg_fullgraph1 = "0001000010" else '0'; 
		reg_q214 <= '1' when reg_fullgraph1 = "0001000011" else '0'; 
		reg_q2712 <= '1' when reg_fullgraph1 = "0001000100" else '0'; 
		reg_q2714 <= '1' when reg_fullgraph1 = "0001000101" else '0'; 
		reg_q2032 <= '1' when reg_fullgraph1 = "0001000110" else '0'; 
		reg_q1945 <= '1' when reg_fullgraph1 = "0001000111" else '0'; 
		reg_q1947 <= '1' when reg_fullgraph1 = "0001001000" else '0'; 
		reg_q124 <= '1' when reg_fullgraph1 = "0001001001" else '0'; 
		reg_q126 <= '1' when reg_fullgraph1 = "0001001010" else '0'; 
		reg_q2272 <= '1' when reg_fullgraph1 = "0001001011" else '0'; 
		reg_q2274 <= '1' when reg_fullgraph1 = "0001001100" else '0'; 
		reg_q42 <= '1' when reg_fullgraph1 = "0001001101" else '0'; 
		reg_q44 <= '1' when reg_fullgraph1 = "0001001110" else '0'; 
		reg_q2028 <= '1' when reg_fullgraph1 = "0001001111" else '0'; 
		reg_q2030 <= '1' when reg_fullgraph1 = "0001010000" else '0'; 
		reg_q1315 <= '1' when reg_fullgraph1 = "0001010001" else '0'; 
		reg_q2704 <= '1' when reg_fullgraph1 = "0001010010" else '0'; 
		reg_q2706 <= '1' when reg_fullgraph1 = "0001010011" else '0'; 
		reg_q1994 <= '1' when reg_fullgraph1 = "0001010100" else '0'; 
		reg_q1804 <= '1' when reg_fullgraph1 = "0001010101" else '0'; 
		reg_q1806 <= '1' when reg_fullgraph1 = "0001010110" else '0'; 
		reg_q698 <= '1' when reg_fullgraph1 = "0001010111" else '0'; 
		reg_q700 <= '1' when reg_fullgraph1 = "0001011000" else '0'; 
		reg_q2617 <= '1' when reg_fullgraph1 = "0001011001" else '0'; 
		reg_q768 <= '1' when reg_fullgraph1 = "0001011010" else '0'; 
		reg_q2752 <= '1' when reg_fullgraph1 = "0001011011" else '0'; 
		reg_q2754 <= '1' when reg_fullgraph1 = "0001011100" else '0'; 
		reg_q1701 <= '1' when reg_fullgraph1 = "0001011101" else '0'; 
		reg_q1703 <= '1' when reg_fullgraph1 = "0001011110" else '0'; 
		reg_q120 <= '1' when reg_fullgraph1 = "0001011111" else '0'; 
		reg_q122 <= '1' when reg_fullgraph1 = "0001100000" else '0'; 
		reg_q2726 <= '1' when reg_fullgraph1 = "0001100001" else '0'; 
		reg_q2728 <= '1' when reg_fullgraph1 = "0001100010" else '0'; 
		reg_q2040 <= '1' when reg_fullgraph1 = "0001100011" else '0'; 
		reg_q2042 <= '1' when reg_fullgraph1 = "0001100100" else '0'; 
		reg_q208 <= '1' when reg_fullgraph1 = "0001100101" else '0'; 
		reg_q1126 <= '1' when reg_fullgraph1 = "0001100110" else '0'; 
		reg_q1212 <= '1' when reg_fullgraph1 = "0001100111" else '0'; 
		reg_q1214 <= '1' when reg_fullgraph1 = "0001101000" else '0'; 
		reg_q2316 <= '1' when reg_fullgraph1 = "0001101001" else '0'; 
		reg_q2018 <= '1' when reg_fullgraph1 = "0001101010" else '0'; 
		reg_q355 <= '1' when reg_fullgraph1 = "0001101011" else '0'; 
		reg_q357 <= '1' when reg_fullgraph1 = "0001101100" else '0'; 
		reg_q776 <= '1' when reg_fullgraph1 = "0001101101" else '0'; 
		reg_q778 <= '1' when reg_fullgraph1 = "0001101110" else '0'; 
		reg_q58 <= '1' when reg_fullgraph1 = "0001101111" else '0'; 
		reg_q60 <= '1' when reg_fullgraph1 = "0001110000" else '0'; 
		reg_q1183 <= '1' when reg_fullgraph1 = "0001110001" else '0'; 
		reg_q718 <= '1' when reg_fullgraph1 = "0001110010" else '0'; 
		reg_q972 <= '1' when reg_fullgraph1 = "0001110011" else '0'; 
		reg_q974 <= '1' when reg_fullgraph1 = "0001110100" else '0'; 
		reg_q2012 <= '1' when reg_fullgraph1 = "0001110101" else '0'; 
		reg_q2014 <= '1' when reg_fullgraph1 = "0001110110" else '0'; 
		reg_q2383 <= '1' when reg_fullgraph1 = "0001110111" else '0'; 
		reg_q2385 <= '1' when reg_fullgraph1 = "0001111000" else '0'; 
		reg_q782 <= '1' when reg_fullgraph1 = "0001111001" else '0'; 
		reg_q784 <= '1' when reg_fullgraph1 = "0001111010" else '0'; 
		reg_q501 <= '1' when reg_fullgraph1 = "0001111011" else '0'; 
		reg_q1707 <= '1' when reg_fullgraph1 = "0001111100" else '0'; 
		reg_q1949 <= '1' when reg_fullgraph1 = "0001111101" else '0'; 
		reg_q52 <= '1' when reg_fullgraph1 = "0001111110" else '0'; 
		reg_q54 <= '1' when reg_fullgraph1 = "0001111111" else '0'; 
		reg_q2621 <= '1' when reg_fullgraph1 = "0010000000" else '0'; 
		reg_q238 <= '1' when reg_fullgraph1 = "0010000001" else '0'; 
		reg_q240 <= '1' when reg_fullgraph1 = "0010000010" else '0'; 
		reg_q716 <= '1' when reg_fullgraph1 = "0010000011" else '0'; 
		reg_q1187 <= '1' when reg_fullgraph1 = "0010000100" else '0'; 
		reg_q1189 <= '1' when reg_fullgraph1 = "0010000101" else '0'; 
		reg_q2597 <= '1' when reg_fullgraph1 = "0010000110" else '0'; 
		reg_q2599 <= '1' when reg_fullgraph1 = "0010000111" else '0'; 
		reg_q141 <= '1' when reg_fullgraph1 = "0010001000" else '0'; 
		reg_q143 <= '1' when reg_fullgraph1 = "0010001001" else '0'; 
		reg_q1768 <= '1' when reg_fullgraph1 = "0010001010" else '0'; 
		reg_q1770 <= '1' when reg_fullgraph1 = "0010001011" else '0'; 
		reg_q2288 <= '1' when reg_fullgraph1 = "0010001100" else '0'; 
		reg_q2000 <= '1' when reg_fullgraph1 = "0010001101" else '0'; 
		reg_q1717 <= '1' when reg_fullgraph1 = "0010001110" else '0'; 
		reg_q2225 <= '1' when reg_fullgraph1 = "0010001111" else '0'; 
		reg_q2227 <= '1' when reg_fullgraph1 = "0010010000" else '0'; 
		reg_q50 <= '1' when reg_fullgraph1 = "0010010001" else '0'; 
		reg_q557 <= '1' when reg_fullgraph1 = "0010010010" else '0'; 
		reg_q559 <= '1' when reg_fullgraph1 = "0010010011" else '0'; 
		reg_q478 <= '1' when reg_fullgraph1 = "0010010100" else '0'; 
		reg_q2619 <= '1' when reg_fullgraph1 = "0010010101" else '0'; 
		reg_q2004 <= '1' when reg_fullgraph1 = "0010010110" else '0'; 
		reg_q212 <= '1' when reg_fullgraph1 = "0010010111" else '0'; 
		reg_q2276 <= '1' when reg_fullgraph1 = "0010011000" else '0'; 
		reg_q2278 <= '1' when reg_fullgraph1 = "0010011001" else '0'; 
		reg_q1778 <= '1' when reg_fullgraph1 = "0010011010" else '0'; 
		reg_q1780 <= '1' when reg_fullgraph1 = "0010011011" else '0'; 
		reg_q2264 <= '1' when reg_fullgraph1 = "0010011100" else '0'; 
		reg_q2266 <= '1' when reg_fullgraph1 = "0010011101" else '0'; 
		reg_q1136 <= '1' when reg_fullgraph1 = "0010011110" else '0'; 
		reg_q69 <= '1' when reg_fullgraph1 = "0010011111" else '0'; 
		reg_q71 <= '1' when reg_fullgraph1 = "0010100000" else '0'; 
		reg_q171 <= '1' when reg_fullgraph1 = "0010100001" else '0'; 
		reg_q1721 <= '1' when reg_fullgraph1 = "0010100010" else '0'; 
		reg_q2016 <= '1' when reg_fullgraph1 = "0010100011" else '0'; 
		reg_q1100 <= '1' when reg_fullgraph1 = "0010100100" else '0'; 
		reg_q1102 <= '1' when reg_fullgraph1 = "0010100101" else '0'; 
		reg_q722 <= '1' when reg_fullgraph1 = "0010100110" else '0'; 
		reg_q724 <= '1' when reg_fullgraph1 = "0010100111" else '0'; 
		reg_q1073 <= '1' when reg_fullgraph1 = "0010101000" else '0'; 
		reg_q1075 <= '1' when reg_fullgraph1 = "0010101001" else '0'; 
		reg_q2044 <= '1' when reg_fullgraph1 = "0010101010" else '0'; 
		reg_q2046 <= '1' when reg_fullgraph1 = "0010101011" else '0'; 
		reg_q258 <= '1' when reg_fullgraph1 = "0010101100" else '0'; 
		reg_q260 <= '1' when reg_fullgraph1 = "0010101101" else '0'; 
		reg_q236 <= '1' when reg_fullgraph1 = "0010101110" else '0'; 
		reg_q1800 <= '1' when reg_fullgraph1 = "0010101111" else '0'; 
		reg_q1802 <= '1' when reg_fullgraph1 = "0010110000" else '0'; 
		reg_q145 <= '1' when reg_fullgraph1 = "0010110001" else '0'; 
		reg_q1723 <= '1' when reg_fullgraph1 = "0010110010" else '0'; 
		reg_q511 <= '1' when reg_fullgraph1 = "0010110011" else '0'; 
		reg_q1010 <= '1' when reg_fullgraph1 = "0010110100" else '0'; 
		reg_q555 <= '1' when reg_fullgraph1 = "0010110101" else '0'; 
		reg_q167 <= '1' when reg_fullgraph1 = "0010110110" else '0'; 
		reg_q169 <= '1' when reg_fullgraph1 = "0010110111" else '0'; 
		reg_q2304 <= '1' when reg_fullgraph1 = "0010111000" else '0'; 
		reg_q2306 <= '1' when reg_fullgraph1 = "0010111001" else '0'; 
		reg_q2223 <= '1' when reg_fullgraph1 = "0010111010" else '0'; 
		reg_q1171 <= '1' when reg_fullgraph1 = "0010111011" else '0'; 
		reg_q1173 <= '1' when reg_fullgraph1 = "0010111100" else '0'; 
		reg_q1520 <= '1' when reg_fullgraph1 = "0010111101" else '0'; 
		reg_q147 <= '1' when reg_fullgraph1 = "0010111110" else '0'; 
		reg_q79 <= '1' when reg_fullgraph1 = "0010111111" else '0'; 
		reg_q81 <= '1' when reg_fullgraph1 = "0011000000" else '0'; 
		reg_q242 <= '1' when reg_fullgraph1 = "0011000001" else '0'; 
		reg_q244 <= '1' when reg_fullgraph1 = "0011000010" else '0'; 
		reg_q1911 <= '1' when reg_fullgraph1 = "0011000011" else '0'; 
		reg_q1913 <= '1' when reg_fullgraph1 = "0011000100" else '0'; 
		reg_q190 <= '1' when reg_fullgraph1 = "0011000101" else '0'; 
		reg_q2024 <= '1' when reg_fullgraph1 = "0011000110" else '0'; 
		reg_q2026 <= '1' when reg_fullgraph1 = "0011000111" else '0'; 
		reg_q1159 <= '1' when reg_fullgraph1 = "0011001000" else '0'; 
		reg_q1161 <= '1' when reg_fullgraph1 = "0011001001" else '0'; 
		reg_q1918 <= '1' when reg_fullgraph1 = "0011001010" else '0'; 
		reg_q1766 <= '1' when reg_fullgraph1 = "0011001011" else '0'; 
		reg_q1715 <= '1' when reg_fullgraph1 = "0011001100" else '0'; 
		reg_q530 <= '1' when reg_fullgraph1 = "0011001101" else '0'; 
		reg_q32 <= '1' when reg_fullgraph1 = "0011001110" else '0'; 
		reg_q34 <= '1' when reg_fullgraph1 = "0011001111" else '0'; 
		reg_q990 <= '1' when reg_fullgraph1 = "0011010000" else '0'; 
		reg_q992 <= '1' when reg_fullgraph1 = "0011010001" else '0'; 
		reg_q18 <= '1' when reg_fullgraph1 = "0011010010" else '0'; 
		reg_q20 <= '1' when reg_fullgraph1 = "0011010011" else '0'; 
		reg_q9 <= '1' when reg_fullgraph1 = "0011010100" else '0'; 
		reg_q11 <= '1' when reg_fullgraph1 = "0011010101" else '0'; 
		reg_q1735 <= '1' when reg_fullgraph1 = "0011010110" else '0'; 
		reg_q1737 <= '1' when reg_fullgraph1 = "0011010111" else '0'; 
		reg_q1331 <= '1' when reg_fullgraph1 = "0011011000" else '0'; 
		reg_q1333 <= '1' when reg_fullgraph1 = "0011011001" else '0'; 
		reg_q1713 <= '1' when reg_fullgraph1 = "0011011010" else '0'; 
		reg_q373 <= '1' when reg_fullgraph1 = "0011011011" else '0'; 
		reg_q375 <= '1' when reg_fullgraph1 = "0011011100" else '0'; 
		reg_q2395 <= '1' when reg_fullgraph1 = "0011011101" else '0'; 
		reg_q2397 <= '1' when reg_fullgraph1 = "0011011110" else '0'; 
		reg_q2601 <= '1' when reg_fullgraph1 = "0011011111" else '0'; 
		reg_q77 <= '1' when reg_fullgraph1 = "0011100000" else '0'; 
		reg_q2694 <= '1' when reg_fullgraph1 = "0011100001" else '0'; 
		reg_q2696 <= '1' when reg_fullgraph1 = "0011100010" else '0'; 
		reg_q2310 <= '1' when reg_fullgraph1 = "0011100011" else '0'; 
		reg_q1012 <= '1' when reg_fullgraph1 = "0011100100" else '0'; 
		reg_q1014 <= '1' when reg_fullgraph1 = "0011100101" else '0'; 
		reg_q1193 <= '1' when reg_fullgraph1 = "0011100110" else '0'; 
		reg_q1195 <= '1' when reg_fullgraph1 = "0011100111" else '0'; 
		reg_q2407 <= '1' when reg_fullgraph1 = "0011101000" else '0'; 
		reg_q2409 <= '1' when reg_fullgraph1 = "0011101001" else '0'; 
		reg_q2718 <= '1' when reg_fullgraph1 = "0011101010" else '0'; 
		reg_q2720 <= '1' when reg_fullgraph1 = "0011101011" else '0'; 
		reg_q216 <= '1' when reg_fullgraph1 = "0011101100" else '0'; 
		reg_q1327 <= '1' when reg_fullgraph1 = "0011101101" else '0'; 
		reg_q551 <= '1' when reg_fullgraph1 = "0011101110" else '0'; 
		reg_q2048 <= '1' when reg_fullgraph1 = "0011101111" else '0'; 
		reg_q105 <= '1' when reg_fullgraph1 = "0011110000" else '0'; 
		reg_q1484 <= '1' when reg_fullgraph1 = "0011110001" else '0'; 
		reg_q250 <= '1' when reg_fullgraph1 = "0011110010" else '0'; 
		reg_q252 <= '1' when reg_fullgraph1 = "0011110011" else '0'; 
		reg_q2415 <= '1' when reg_fullgraph1 = "0011110100" else '0'; 
		reg_q2010 <= '1' when reg_fullgraph1 = "0011110101" else '0'; 
		reg_q2585 <= '1' when reg_fullgraph1 = "0011110110" else '0'; 
		reg_q2682 <= '1' when reg_fullgraph1 = "0011110111" else '0'; 
		reg_q996 <= '1' when reg_fullgraph1 = "0011111000" else '0'; 
		reg_q998 <= '1' when reg_fullgraph1 = "0011111001" else '0'; 
		reg_q1808 <= '1' when reg_fullgraph1 = "0011111010" else '0'; 
		reg_q1810 <= '1' when reg_fullgraph1 = "0011111011" else '0'; 
		reg_q1725 <= '1' when reg_fullgraph1 = "0011111100" else '0'; 
		reg_q1727 <= '1' when reg_fullgraph1 = "0011111101" else '0'; 
		reg_q1743 <= '1' when reg_fullgraph1 = "0011111110" else '0'; 
		reg_q1745 <= '1' when reg_fullgraph1 = "0011111111" else '0'; 
		reg_q204 <= '1' when reg_fullgraph1 = "0100000000" else '0'; 
		reg_q206 <= '1' when reg_fullgraph1 = "0100000001" else '0'; 
		reg_q2393 <= '1' when reg_fullgraph1 = "0100000010" else '0'; 
		reg_q1762 <= '1' when reg_fullgraph1 = "0100000011" else '0'; 
		reg_q1764 <= '1' when reg_fullgraph1 = "0100000100" else '0'; 
		reg_q868 <= '1' when reg_fullgraph1 = "0100000101" else '0'; 
		reg_q2684 <= '1' when reg_fullgraph1 = "0100000110" else '0'; 
		reg_q2686 <= '1' when reg_fullgraph1 = "0100000111" else '0'; 
		reg_q746 <= '1' when reg_fullgraph1 = "0100001000" else '0'; 
		reg_q87 <= '1' when reg_fullgraph1 = "0100001001" else '0'; 
		reg_q89 <= '1' when reg_fullgraph1 = "0100001010" else '0'; 
		reg_q5 <= '1' when reg_fullgraph1 = "0100001011" else '0'; 
		reg_q1165 <= '1' when reg_fullgraph1 = "0100001100" else '0'; 
		reg_q1167 <= '1' when reg_fullgraph1 = "0100001101" else '0'; 
		reg_q1208 <= '1' when reg_fullgraph1 = "0100001110" else '0'; 
		reg_q1210 <= '1' when reg_fullgraph1 = "0100001111" else '0'; 
		reg_q254 <= '1' when reg_fullgraph1 = "0100010000" else '0'; 
		reg_q1313 <= '1' when reg_fullgraph1 = "0100010001" else '0'; 
		reg_q1132 <= '1' when reg_fullgraph1 = "0100010010" else '0'; 
		reg_q2308 <= '1' when reg_fullgraph1 = "0100010011" else '0'; 
		reg_q702 <= '1' when reg_fullgraph1 = "0100010100" else '0'; 
		reg_q1081 <= '1' when reg_fullgraph1 = "0100010101" else '0'; 
		reg_q988 <= '1' when reg_fullgraph1 = "0100010110" else '0'; 
		reg_q1689 <= '1' when reg_fullgraph1 = "0100010111" else '0'; 
		reg_q1691 <= '1' when reg_fullgraph1 = "0100011000" else '0'; 
		reg_q2615 <= '1' when reg_fullgraph1 = "0100011001" else '0'; 
		reg_q1514 <= '1' when reg_fullgraph1 = "0100011010" else '0'; 
		reg_q1516 <= '1' when reg_fullgraph1 = "0100011011" else '0'; 
		reg_q740 <= '1' when reg_fullgraph1 = "0100011100" else '0'; 
		reg_q563 <= '1' when reg_fullgraph1 = "0100011101" else '0'; 
		reg_q994 <= '1' when reg_fullgraph1 = "0100011110" else '0'; 
		reg_q2002 <= '1' when reg_fullgraph1 = "0100011111" else '0'; 
		reg_q708 <= '1' when reg_fullgraph1 = "0100100000" else '0'; 
		reg_q710 <= '1' when reg_fullgraph1 = "0100100001" else '0'; 
		reg_q1185 <= '1' when reg_fullgraph1 = "0100100010" else '0'; 
		reg_q2357 <= '1' when reg_fullgraph1 = "0100100011" else '0'; 
		reg_q2359 <= '1' when reg_fullgraph1 = "0100100100" else '0'; 
		reg_q226 <= '1' when reg_fullgraph1 = "0100100101" else '0'; 
		reg_q228 <= '1' when reg_fullgraph1 = "0100100110" else '0'; 
		reg_q1339 <= '1' when reg_fullgraph1 = "0100100111" else '0'; 
		reg_q1341 <= '1' when reg_fullgraph1 = "0100101000" else '0'; 
		reg_q1124 <= '1' when reg_fullgraph1 = "0100101001" else '0'; 
		reg_q1317 <= '1' when reg_fullgraph1 = "0100101010" else '0'; 
		reg_q38 <= '1' when reg_fullgraph1 = "0100101011" else '0'; 
		reg_q673 <= '1' when reg_fullgraph1 = "0100101100" else '0'; 
		reg_q1349 <= '1' when reg_fullgraph1 = "0100101101" else '0'; 
		reg_q1351 <= '1' when reg_fullgraph1 = "0100101110" else '0'; 
		reg_q1494 <= '1' when reg_fullgraph1 = "0100101111" else '0'; 
		reg_q1496 <= '1' when reg_fullgraph1 = "0100110000" else '0'; 
		reg_q532 <= '1' when reg_fullgraph1 = "0100110001" else '0'; 
		reg_q534 <= '1' when reg_fullgraph1 = "0100110010" else '0'; 
		reg_q967 <= '1' when reg_fullgraph1 = "0100110011" else '0'; 
		reg_q955 <= '1' when reg_fullgraph1 = "0100110100" else '0'; 
		reg_q270 <= '1' when reg_fullgraph1 = "0100110101" else '0'; 
		reg_q272 <= '1' when reg_fullgraph1 = "0100110110" else '0'; 
		reg_q734 <= '1' when reg_fullgraph1 = "0100110111" else '0'; 
		reg_q736 <= '1' when reg_fullgraph1 = "0100111000" else '0'; 
		reg_q1004 <= '1' when reg_fullgraph1 = "0100111001" else '0'; 
		reg_q1006 <= '1' when reg_fullgraph1 = "0100111010" else '0'; 
		reg_q1077 <= '1' when reg_fullgraph1 = "0100111011" else '0'; 
		reg_q1079 <= '1' when reg_fullgraph1 = "0100111100" else '0'; 
		reg_q2268 <= '1' when reg_fullgraph1 = "0100111101" else '0'; 
		reg_q2270 <= '1' when reg_fullgraph1 = "0100111110" else '0'; 
		reg_q2298 <= '1' when reg_fullgraph1 = "0100111111" else '0'; 
		reg_q2300 <= '1' when reg_fullgraph1 = "0101000000" else '0'; 
		reg_q1905 <= '1' when reg_fullgraph1 = "0101000001" else '0'; 
		reg_q1163 <= '1' when reg_fullgraph1 = "0101000010" else '0'; 
		reg_q1812 <= '1' when reg_fullgraph1 = "0101000011" else '0'; 
		reg_q1814 <= '1' when reg_fullgraph1 = "0101000100" else '0'; 
		reg_q1000 <= '1' when reg_fullgraph1 = "0101000101" else '0'; 
		reg_q1069 <= '1' when reg_fullgraph1 = "0101000110" else '0'; 
		reg_q274 <= '1' when reg_fullgraph1 = "0101000111" else '0'; 
		reg_q1794 <= '1' when reg_fullgraph1 = "0101001000" else '0'; 
		reg_q1796 <= '1' when reg_fullgraph1 = "0101001001" else '0'; 
		reg_q280 <= '1' when reg_fullgraph1 = "0101001010" else '0'; 
		reg_q2347 <= '1' when reg_fullgraph1 = "0101001011" else '0'; 
		reg_q2349 <= '1' when reg_fullgraph1 = "0101001100" else '0'; 
		reg_q387 <= '1' when reg_fullgraph1 = "0101001101" else '0'; 
		reg_q389 <= '1' when reg_fullgraph1 = "0101001110" else '0'; 
		reg_q1343 <= '1' when reg_fullgraph1 = "0101001111" else '0'; 
		reg_q1729 <= '1' when reg_fullgraph1 = "0101010000" else '0'; 
		reg_q2522 <= '1' when reg_fullgraph1 = "0101010001" else '0'; 
		reg_q2722 <= '1' when reg_fullgraph1 = "0101010010" else '0'; 
		reg_q2724 <= '1' when reg_fullgraph1 = "0101010011" else '0'; 
		reg_q1776 <= '1' when reg_fullgraph1 = "0101010100" else '0'; 
		reg_q2286 <= '1' when reg_fullgraph1 = "0101010101" else '0'; 
		reg_q264 <= '1' when reg_fullgraph1 = "0101010110" else '0'; 
		reg_q2373 <= '1' when reg_fullgraph1 = "0101010111" else '0'; 
		reg_q2375 <= '1' when reg_fullgraph1 = "0101011000" else '0'; 
		reg_q2702 <= '1' when reg_fullgraph1 = "0101011001" else '0'; 
		reg_q276 <= '1' when reg_fullgraph1 = "0101011010" else '0'; 
		reg_q278 <= '1' when reg_fullgraph1 = "0101011011" else '0'; 
		reg_q383 <= '1' when reg_fullgraph1 = "0101011100" else '0'; 
		reg_q385 <= '1' when reg_fullgraph1 = "0101011101" else '0'; 
		reg_q679 <= '1' when reg_fullgraph1 = "0101011110" else '0'; 
		reg_q2284 <= '1' when reg_fullgraph1 = "0101011111" else '0'; 
		reg_q1008 <= '1' when reg_fullgraph1 = "0101100000" else '0'; 
		reg_q83 <= '1' when reg_fullgraph1 = "0101100001" else '0'; 
		reg_q85 <= '1' when reg_fullgraph1 = "0101100010" else '0'; 
		reg_q1181 <= '1' when reg_fullgraph1 = "0101100011" else '0'; 
		reg_q1345 <= '1' when reg_fullgraph1 = "0101100100" else '0'; 
		reg_q730 <= '1' when reg_fullgraph1 = "0101100101" else '0'; 
		reg_q2341 <= '1' when reg_fullgraph1 = "0101100110" else '0'; 
		reg_q2343 <= '1' when reg_fullgraph1 = "0101100111" else '0'; 
		reg_q669 <= '1' when reg_fullgraph1 = "0101101000" else '0'; 
		reg_q1518 <= '1' when reg_fullgraph1 = "0101101001" else '0'; 
		reg_q1112 <= '1' when reg_fullgraph1 = "0101101010" else '0'; 
		reg_q1114 <= '1' when reg_fullgraph1 = "0101101011" else '0'; 
		reg_q230 <= '1' when reg_fullgraph1 = "0101101100" else '0'; 
		reg_q1118 <= '1' when reg_fullgraph1 = "0101101101" else '0'; 
		reg_q1120 <= '1' when reg_fullgraph1 = "0101101110" else '0'; 
		reg_q14 <= '1' when reg_fullgraph1 = "0101101111" else '0'; 
		reg_q16 <= '1' when reg_fullgraph1 = "0101110000" else '0'; 
		reg_q1071 <= '1' when reg_fullgraph1 = "0101110001" else '0'; 
		reg_q2256 <= '1' when reg_fullgraph1 = "0101110010" else '0'; 
		reg_q2258 <= '1' when reg_fullgraph1 = "0101110011" else '0'; 
		reg_q1335 <= '1' when reg_fullgraph1 = "0101110100" else '0'; 
		reg_q681 <= '1' when reg_fullgraph1 = "0101110101" else '0'; 
		reg_q683 <= '1' when reg_fullgraph1 = "0101110110" else '0'; 
		reg_q1984 <= '1' when reg_fullgraph1 = "0101110111" else '0'; 
		reg_q1986 <= '1' when reg_fullgraph1 = "0101111000" else '0'; 
		reg_q26 <= '1' when reg_fullgraph1 = "0101111001" else '0'; 
		reg_q28 <= '1' when reg_fullgraph1 = "0101111010" else '0'; 
		reg_q22 <= '1' when reg_fullgraph1 = "0101111011" else '0'; 
		reg_q1699 <= '1' when reg_fullgraph1 = "0101111100" else '0'; 
		reg_q1175 <= '1' when reg_fullgraph1 = "0101111101" else '0'; 
		reg_q1177 <= '1' when reg_fullgraph1 = "0101111110" else '0'; 
		reg_q381 <= '1' when reg_fullgraph1 = "0101111111" else '0'; 
		reg_q2365 <= '1' when reg_fullgraph1 = "0110000000" else '0'; 
		reg_q2367 <= '1' when reg_fullgraph1 = "0110000001" else '0'; 
		reg_q192 <= '1' when reg_fullgraph1 = "0110000010" else '0'; 
		reg_q194 <= '1' when reg_fullgraph1 = "0110000011" else '0'; 
		reg_q1488 <= '1' when reg_fullgraph1 = "0110000100" else '0'; 
		reg_q1490 <= '1' when reg_fullgraph1 = "0110000101" else '0'; 
		reg_q1758 <= '1' when reg_fullgraph1 = "0110000110" else '0'; 
		reg_q1760 <= '1' when reg_fullgraph1 = "0110000111" else '0'; 
		reg_q2331 <= '1' when reg_fullgraph1 = "0110001000" else '0'; 
		reg_q2333 <= '1' when reg_fullgraph1 = "0110001001" else '0'; 
		reg_q163 <= '1' when reg_fullgraph1 = "0110001010" else '0'; 
		reg_q165 <= '1' when reg_fullgraph1 = "0110001011" else '0'; 
		reg_q2252 <= '1' when reg_fullgraph1 = "0110001100" else '0'; 
		reg_q2254 <= '1' when reg_fullgraph1 = "0110001101" else '0'; 
		reg_q1988 <= '1' when reg_fullgraph1 = "0110001110" else '0'; 
		reg_q553 <= '1' when reg_fullgraph1 = "0110001111" else '0'; 
		reg_q671 <= '1' when reg_fullgraph1 = "0110010000" else '0'; 
		reg_q2716 <= '1' when reg_fullgraph1 = "0110010001" else '0'; 
		reg_q2690 <= '1' when reg_fullgraph1 = "0110010010" else '0'; 
		reg_q2692 <= '1' when reg_fullgraph1 = "0110010011" else '0'; 
		reg_q1741 <= '1' when reg_fullgraph1 = "0110010100" else '0'; 
		reg_q1337 <= '1' when reg_fullgraph1 = "0110010101" else '0'; 
		reg_q75 <= '1' when reg_fullgraph1 = "0110010110" else '0'; 
		reg_q24 <= '1' when reg_fullgraph1 = "0110010111" else '0'; 
		reg_q1191 <= '1' when reg_fullgraph1 = "0110011000" else '0'; 
		reg_q2603 <= '1' when reg_fullgraph1 = "0110011001" else '0'; 
		reg_q2605 <= '1' when reg_fullgraph1 = "0110011010" else '0'; 
		reg_q1932 <= '1' when reg_fullgraph1 = "0110011011" else '0'; 
		reg_q950 <= '1' when reg_fullgraph1 = "0110011100" else '0'; 
		reg_q2710 <= '1' when reg_fullgraph1 = "0110011101" else '0'; 
		reg_q36 <= '1' when reg_fullgraph1 = "0110011110" else '0'; 
		reg_q1155 <= '1' when reg_fullgraph1 = "0110011111" else '0'; 
		reg_q1157 <= '1' when reg_fullgraph1 = "0110100000" else '0'; 
		reg_q153 <= '1' when reg_fullgraph1 = "0110100001" else '0'; 
		reg_q1169 <= '1' when reg_fullgraph1 = "0110100010" else '0'; 
		reg_q266 <= '1' when reg_fullgraph1 = "0110100011" else '0'; 
		reg_q507 <= '1' when reg_fullgraph1 = "0110100100" else '0'; 
		reg_q509 <= '1' when reg_fullgraph1 = "0110100101" else '0'; 
		reg_q2611 <= '1' when reg_fullgraph1 = "0110100110" else '0'; 
		reg_q2613 <= '1' when reg_fullgraph1 = "0110100111" else '0'; 
		reg_q2700 <= '1' when reg_fullgraph1 = "0110101000" else '0'; 
		reg_q196 <= '1' when reg_fullgraph1 = "0110101001" else '0'; 
		reg_q2708 <= '1' when reg_fullgraph1 = "0110101010" else '0'; 
		reg_q561 <= '1' when reg_fullgraph1 = "0110101011" else '0'; 
		reg_q161 <= '1' when reg_fullgraph1 = "0110101100" else '0'; 
		reg_q224 <= '1' when reg_fullgraph1 = "0110101101" else '0'; 
		reg_q232 <= '1' when reg_fullgraph1 = "0110101110" else '0'; 
		reg_q234 <= '1' when reg_fullgraph1 = "0110101111" else '0'; 
		reg_q2593 <= '1' when reg_fullgraph1 = "0110110000" else '0'; 
		reg_q2595 <= '1' when reg_fullgraph1 = "0110110001" else '0'; 
		reg_q594 <= '1' when reg_fullgraph1 = "0110110010" else '0'; 
		reg_q2698 <= '1' when reg_fullgraph1 = "0110110011" else '0'; 
		reg_q67 <= '1' when reg_fullgraph1 = "0110110100" else '0'; 
		reg_q2302 <= '1' when reg_fullgraph1 = "0110110101" else '0'; 
		reg_q2351 <= '1' when reg_fullgraph1 = "0110110110" else '0'; 
		reg_q2353 <= '1' when reg_fullgraph1 = "0110110111" else '0'; 
		reg_q1930 <= '1' when reg_fullgraph1 = "0110111000" else '0'; 
		reg_q1695 <= '1' when reg_fullgraph1 = "0110111001" else '0'; 
		reg_q1697 <= '1' when reg_fullgraph1 = "0110111010" else '0'; 
		reg_q268 <= '1' when reg_fullgraph1 = "0110111011" else '0'; 
		reg_q1085 <= '1' when reg_fullgraph1 = "0110111100" else '0'; 
		reg_q685 <= '1' when reg_fullgraph1 = "0110111101" else '0'; 
		reg_q1739 <= '1' when reg_fullgraph1 = "0110111110" else '0'; 
		reg_q2361 <= '1' when reg_fullgraph1 = "0110111111" else '0'; 
		reg_q262 <= '1' when reg_fullgraph1 = "0111000000" else '0'; 
		reg_q46 <= '1' when reg_fullgraph1 = "0111000001" else '0'; 
		reg_q1747 <= '1' when reg_fullgraph1 = "0111000010" else '0'; 
		reg_q2371 <= '1' when reg_fullgraph1 = "0111000011" else '0'; 
		reg_q2324 <= '1' when reg_fullgraph1 = "0111000100" else '0'; 
		reg_q1980 <= '1' when reg_fullgraph1 = "0111000101" else '0'; 
		reg_q2379 <= '1' when reg_fullgraph1 = "0111000110" else '0'; 
		reg_q139 <= '1' when reg_fullgraph1 = "0111000111" else '0'; 
		reg_q2377 <= '1' when reg_fullgraph1 = "0111001000" else '0'; 
		reg_q93 <= '1' when reg_fullgraph1 = "0111001001" else '0'; 
		reg_q95 <= '1' when reg_fullgraph1 = "0111001010" else '0'; 
		reg_q1798 <= '1' when reg_fullgraph1 = "0111001011" else '0'; 
		reg_q2730 <= '1' when reg_fullgraph1 = "0111001100" else '0'; 
		reg_q2732 <= '1' when reg_fullgraph1 = "0111001101" else '0'; 
		reg_q1329 <= '1' when reg_fullgraph1 = "0111001110" else '0'; 
		reg_q155 <= '1' when reg_fullgraph1 = "0111001111" else '0'; 
		reg_q157 <= '1' when reg_fullgraph1 = "0111010000" else '0'; 
		reg_q1784 <= '1' when reg_fullgraph1 = "0111010001" else '0'; 
		reg_q202 <= '1' when reg_fullgraph1 = "0111010010" else '0'; 
		reg_q1002 <= '1' when reg_fullgraph1 = "0111010011" else '0'; 
		reg_q2335 <= '1' when reg_fullgraph1 = "0111010100" else '0'; 
		reg_q1792 <= '1' when reg_fullgraph1 = "0111010101" else '0'; 
		reg_q1134 <= '1' when reg_fullgraph1 = "0111010110" else '0'; 
		reg_q677 <= '1' when reg_fullgraph1 = "0111010111" else '0'; 
		reg_q2734 <= '1' when reg_fullgraph1 = "0111011000" else '0'; 
		reg_q2322 <= '1' when reg_fullgraph1 = "0111011001" else '0'; 
		reg_q1140 <= '1' when reg_fullgraph1 = "0111011010" else '0'; 
		reg_q2403 <= '1' when reg_fullgraph1 = "0111011011" else '0'; 
		reg_q2405 <= '1' when reg_fullgraph1 = "0111011100" else '0'; 
		reg_q2320 <= '1' when reg_fullgraph1 = "0111011101" else '0'; 
		reg_q1153 <= '1' when reg_fullgraph1 = "0111011110" else '0'; 
		reg_q505 <= '1' when reg_fullgraph1 = "0111011111" else '0'; 
		reg_q1687 <= '1' when reg_fullgraph1 = "0111100000" else '0'; 
		reg_q65 <= '1' when reg_fullgraph1 = "0111100001" else '0'; 
		reg_q56 <= '1' when reg_fullgraph1 = "0111100010" else '0'; 
		reg_q687 <= '1' when reg_fullgraph1 = "0111100011" else '0'; 
		reg_q365 <= '1' when reg_fullgraph1 = "0111100100" else '0'; 
		reg_q367 <= '1' when reg_fullgraph1 = "0111100101" else '0'; 
		reg_q2260 <= '1' when reg_fullgraph1 = "0111100110" else '0'; 
		reg_q2262 <= '1' when reg_fullgraph1 = "0111100111" else '0'; 
		reg_q363 <= '1' when reg_fullgraph1 = "0111101000" else '0'; 
		reg_q1104 <= '1' when reg_fullgraph1 = "0111101001" else '0'; 
		reg_q1106 <= '1' when reg_fullgraph1 = "0111101010" else '0'; 
		reg_q728 <= '1' when reg_fullgraph1 = "0111101011" else '0'; 
		reg_q957 <= '1' when reg_fullgraph1 = "0111101100" else '0'; 
		reg_q1506 <= '1' when reg_fullgraph1 = "0111101101" else '0'; 
		reg_q137 <= '1' when reg_fullgraph1 = "0111101110" else '0'; 
		reg_q2337 <= '1' when reg_fullgraph1 = "0111101111" else '0'; 
		reg_q2339 <= '1' when reg_fullgraph1 = "0111110000" else '0'; 
		reg_q986 <= '1' when reg_fullgraph1 = "0111110001" else '0'; 
		reg_q738 <= '1' when reg_fullgraph1 = "0111110010" else '0'; 
		reg_q1116 <= '1' when reg_fullgraph1 = "0111110011" else '0'; 
		reg_q91 <= '1' when reg_fullgraph1 = "0111110100" else '0'; 
		reg_q1179 <= '1' when reg_fullgraph1 = "0111110101" else '0'; 
		reg_q1693 <= '1' when reg_fullgraph1 = "0111110110" else '0'; 
		reg_q2391 <= '1' when reg_fullgraph1 = "0111110111" else '0'; 
		reg_q2607 <= '1' when reg_fullgraph1 = "0111111000" else '0'; 
		reg_q2609 <= '1' when reg_fullgraph1 = "0111111001" else '0'; 
		reg_q1087 <= '1' when reg_fullgraph1 = "0111111010" else '0'; 
		reg_q1786 <= '1' when reg_fullgraph1 = "0111111011" else '0'; 
		reg_q1788 <= '1' when reg_fullgraph1 = "0111111100" else '0'; 
		reg_q1016 <= '1' when reg_fullgraph1 = "0111111101" else '0'; 
		reg_q706 <= '1' when reg_fullgraph1 = "0111111110" else '0'; 
		reg_q2355 <= '1' when reg_fullgraph1 = "0111111111" else '0'; 
		reg_q2688 <= '1' when reg_fullgraph1 = "1000000000" else '0'; 
		reg_q222 <= '1' when reg_fullgraph1 = "1000000001" else '0'; 
		reg_q248 <= '1' when reg_fullgraph1 = "1000000010" else '0'; 
		reg_q1353 <= '1' when reg_fullgraph1 = "1000000011" else '0'; 
		reg_q63 <= '1' when reg_fullgraph1 = "1000000100" else '0'; 
		reg_q984 <= '1' when reg_fullgraph1 = "1000000101" else '0'; 
		reg_q2748 <= '1' when reg_fullgraph1 = "1000000110" else '0'; 
		reg_q1018 <= '1' when reg_fullgraph1 = "1000000111" else '0'; 
		reg_q2411 <= '1' when reg_fullgraph1 = "1000001000" else '0'; 
		reg_q2589 <= '1' when reg_fullgraph1 = "1000001001" else '0'; 
		reg_q2591 <= '1' when reg_fullgraph1 = "1000001010" else '0'; 
		reg_q1982 <= '1' when reg_fullgraph1 = "1000001011" else '0'; 
		reg_q2401 <= '1' when reg_fullgraph1 = "1000001100" else '0'; 
		reg_q1319 <= '1' when reg_fullgraph1 = "1000001101" else '0'; 
		reg_q726 <= '1' when reg_fullgraph1 = "1000001110" else '0'; 
		reg_q1108 <= '1' when reg_fullgraph1 = "1000001111" else '0'; 
		reg_q1110 <= '1' when reg_fullgraph1 = "1000010000" else '0'; 
		reg_q1355 <= '1' when reg_fullgraph1 = "1000010001" else '0'; 
		reg_q704 <= '1' when reg_fullgraph1 = "1000010010" else '0'; 
		reg_q1122 <= '1' when reg_fullgraph1 = "1000010011" else '0'; 
		reg_q1749 <= '1' when reg_fullgraph1 = "1000010100" else '0'; 
		reg_q159 <= '1' when reg_fullgraph1 = "1000010101" else '0'; 
		reg_q2587 <= '1' when reg_fullgraph1 = "1000010110" else '0'; 
		reg_q2345 <= '1' when reg_fullgraph1 = "1000010111" else '0'; 
		reg_q2750 <= '1' when reg_fullgraph1 = "1000011000" else '0'; 
		reg_q1937 <= '1' when reg_fullgraph1 = "1000011001" else '0'; 
		reg_q1705 <= '1' when reg_fullgraph1 = "1000011010" else '0'; 
		reg_q748 <= '1' when reg_fullgraph1 = "1000011011" else '0'; 
		reg_q2369 <= '1' when reg_fullgraph1 = "1000011100" else '0'; 
		reg_q596 <= '1' when reg_fullgraph1 = "1000011101" else '0'; 
		reg_q598 <= '1' when reg_fullgraph1 = "1000011110" else '0'; 
		reg_q1321 <= '1' when reg_fullgraph1 = "1000011111" else '0'; 
		reg_q2318 <= '1' when reg_fullgraph1 = "1000100000" else '0'; 
		reg_q976 <= '1' when reg_fullgraph1 = "1000100001" else '0'; 
		reg_q1782 <= '1' when reg_fullgraph1 = "1000100010" else '0'; 
		reg_q7 <= '1' when reg_fullgraph1 = "1000100011" else '0'; 
		reg_q2248 <= '1' when reg_fullgraph1 = "1000100100" else '0'; 
		reg_q103 <= '1' when reg_fullgraph1 = "1000100101" else '0'; 
		reg_q513 <= '1' when reg_fullgraph1 = "1000100110" else '0'; 
		reg_q980 <= '1' when reg_fullgraph1 = "1000100111" else '0'; 
		reg_q982 <= '1' when reg_fullgraph1 = "1000101000" else '0'; 
		reg_q246 <= '1' when reg_fullgraph1 = "1000101001" else '0'; 
		reg_q965 <= '1' when reg_fullgraph1 = "1000101010" else '0'; 
		reg_q1508 <= '1' when reg_fullgraph1 = "1000101011" else '0'; 
		reg_q1067 <= '1' when reg_fullgraph1 = "1000101100" else '0'; 
		reg_q48 <= '1' when reg_fullgraph1 = "1000101101" else '0'; 
		reg_q1347 <= '1' when reg_fullgraph1 = "1000101110" else '0'; 
		reg_q1091 <= '1' when reg_fullgraph1 = "1000101111" else '0'; 
		reg_q1093 <= '1' when reg_fullgraph1 = "1000110000" else '0'; 
		reg_q1751 <= '1' when reg_fullgraph1 = "1000110001" else '0'; 
		reg_q1790 <= '1' when reg_fullgraph1 = "1000110010" else '0'; 
		reg_q750 <= '1' when reg_fullgraph1 = "1000110011" else '0'; 
		reg_q1492 <= '1' when reg_fullgraph1 = "1000110100" else '0'; 
		reg_q1928 <= '1' when reg_fullgraph1 = "1000110101" else '0'; 
		reg_q1089 <= '1' when reg_fullgraph1 = "1000110110" else '0'; 
		reg_q1197 <= '1' when reg_fullgraph1 = "1000110111" else '0'; 
		reg_q600 <= '1' when reg_fullgraph1 = "1000111000" else '0'; 
		reg_q602 <= '1' when reg_fullgraph1 = "1000111001" else '0'; 
		reg_q536 <= '1' when reg_fullgraph1 = "1000111010" else '0'; 
		reg_q538 <= '1' when reg_fullgraph1 = "1000111011" else '0'; 
		reg_q2250 <= '1' when reg_fullgraph1 = "1000111100" else '0'; 
		reg_q73 <= '1' when reg_fullgraph1 = "1000111101" else '0'; 
		reg_q978 <= '1' when reg_fullgraph1 = "1000111110" else '0'; 
		reg_q256 <= '1' when reg_fullgraph1 = "1000111111" else '0'; 
		reg_q128 <= '1' when reg_fullgraph1 = "1001000000" else '0'; 
		reg_q130 <= '1' when reg_fullgraph1 = "1001000001" else '0'; 
		reg_q959 <= '1' when reg_fullgraph1 = "1001000010" else '0'; 
		reg_q960 <= '1' when reg_fullgraph1 = "1001000011" else '0'; 
		reg_q2413 <= '1' when reg_fullgraph1 = "1001000100" else '0'; 
		reg_q752 <= '1' when reg_fullgraph1 = "1001000101" else '0'; 
		reg_q1216 <= '1' when reg_fullgraph1 = "1001000110" else '0'; 
		reg_q198 <= '1' when reg_fullgraph1 = "1001000111" else '0'; 
		reg_q1142 <= '1' when reg_fullgraph1 = "1001001000" else '0'; 
		reg_q2755 <= '1' when reg_fullgraph1 = "1001001001" else '0'; 
		reg_q689 <= '1' when reg_fullgraph1 = "1001001010" else '0'; 
		reg_q97 <= '1' when reg_fullgraph1 = "1001001011" else '0'; 
		reg_q754 <= '1' when reg_fullgraph1 = "1001001100" else '0'; 
		reg_q1753 <= '1' when reg_fullgraph1 = "1001001101" else '0'; 
		reg_q691 <= '1' when reg_fullgraph1 = "1001001110" else '0'; 
		reg_q200 <= '1' when reg_fullgraph1 = "1001001111" else '0'; 
		reg_q1020 <= '1' when reg_fullgraph1 = "1001010000" else '0'; 
--end decoder 

reg_q772_in <= (reg_q772 AND symb_decoder(16#ff#)) OR
 					(reg_q772 AND symb_decoder(16#81#)) OR
 					(reg_q772 AND symb_decoder(16#d7#)) OR
 					(reg_q772 AND symb_decoder(16#9e#)) OR
 					(reg_q772 AND symb_decoder(16#15#)) OR
 					(reg_q772 AND symb_decoder(16#56#)) OR
 					(reg_q772 AND symb_decoder(16#24#)) OR
 					(reg_q772 AND symb_decoder(16#7f#)) OR
 					(reg_q772 AND symb_decoder(16#84#)) OR
 					(reg_q772 AND symb_decoder(16#c7#)) OR
 					(reg_q772 AND symb_decoder(16#66#)) OR
 					(reg_q772 AND symb_decoder(16#20#)) OR
 					(reg_q772 AND symb_decoder(16#32#)) OR
 					(reg_q772 AND symb_decoder(16#48#)) OR
 					(reg_q772 AND symb_decoder(16#4d#)) OR
 					(reg_q772 AND symb_decoder(16#a2#)) OR
 					(reg_q772 AND symb_decoder(16#f1#)) OR
 					(reg_q772 AND symb_decoder(16#09#)) OR
 					(reg_q772 AND symb_decoder(16#8d#)) OR
 					(reg_q772 AND symb_decoder(16#c0#)) OR
 					(reg_q772 AND symb_decoder(16#69#)) OR
 					(reg_q772 AND symb_decoder(16#31#)) OR
 					(reg_q772 AND symb_decoder(16#9d#)) OR
 					(reg_q772 AND symb_decoder(16#87#)) OR
 					(reg_q772 AND symb_decoder(16#b6#)) OR
 					(reg_q772 AND symb_decoder(16#97#)) OR
 					(reg_q772 AND symb_decoder(16#cd#)) OR
 					(reg_q772 AND symb_decoder(16#5e#)) OR
 					(reg_q772 AND symb_decoder(16#ba#)) OR
 					(reg_q772 AND symb_decoder(16#bd#)) OR
 					(reg_q772 AND symb_decoder(16#93#)) OR
 					(reg_q772 AND symb_decoder(16#88#)) OR
 					(reg_q772 AND symb_decoder(16#52#)) OR
 					(reg_q772 AND symb_decoder(16#94#)) OR
 					(reg_q772 AND symb_decoder(16#0b#)) OR
 					(reg_q772 AND symb_decoder(16#47#)) OR
 					(reg_q772 AND symb_decoder(16#cc#)) OR
 					(reg_q772 AND symb_decoder(16#4e#)) OR
 					(reg_q772 AND symb_decoder(16#4c#)) OR
 					(reg_q772 AND symb_decoder(16#e5#)) OR
 					(reg_q772 AND symb_decoder(16#07#)) OR
 					(reg_q772 AND symb_decoder(16#e4#)) OR
 					(reg_q772 AND symb_decoder(16#08#)) OR
 					(reg_q772 AND symb_decoder(16#80#)) OR
 					(reg_q772 AND symb_decoder(16#13#)) OR
 					(reg_q772 AND symb_decoder(16#62#)) OR
 					(reg_q772 AND symb_decoder(16#e3#)) OR
 					(reg_q772 AND symb_decoder(16#76#)) OR
 					(reg_q772 AND symb_decoder(16#85#)) OR
 					(reg_q772 AND symb_decoder(16#fd#)) OR
 					(reg_q772 AND symb_decoder(16#ab#)) OR
 					(reg_q772 AND symb_decoder(16#2e#)) OR
 					(reg_q772 AND symb_decoder(16#50#)) OR
 					(reg_q772 AND symb_decoder(16#26#)) OR
 					(reg_q772 AND symb_decoder(16#03#)) OR
 					(reg_q772 AND symb_decoder(16#14#)) OR
 					(reg_q772 AND symb_decoder(16#7c#)) OR
 					(reg_q772 AND symb_decoder(16#d8#)) OR
 					(reg_q772 AND symb_decoder(16#c1#)) OR
 					(reg_q772 AND symb_decoder(16#60#)) OR
 					(reg_q772 AND symb_decoder(16#51#)) OR
 					(reg_q772 AND symb_decoder(16#99#)) OR
 					(reg_q772 AND symb_decoder(16#c4#)) OR
 					(reg_q772 AND symb_decoder(16#4a#)) OR
 					(reg_q772 AND symb_decoder(16#29#)) OR
 					(reg_q772 AND symb_decoder(16#da#)) OR
 					(reg_q772 AND symb_decoder(16#a5#)) OR
 					(reg_q772 AND symb_decoder(16#4f#)) OR
 					(reg_q772 AND symb_decoder(16#17#)) OR
 					(reg_q772 AND symb_decoder(16#53#)) OR
 					(reg_q772 AND symb_decoder(16#28#)) OR
 					(reg_q772 AND symb_decoder(16#8a#)) OR
 					(reg_q772 AND symb_decoder(16#64#)) OR
 					(reg_q772 AND symb_decoder(16#e0#)) OR
 					(reg_q772 AND symb_decoder(16#e8#)) OR
 					(reg_q772 AND symb_decoder(16#23#)) OR
 					(reg_q772 AND symb_decoder(16#bb#)) OR
 					(reg_q772 AND symb_decoder(16#5d#)) OR
 					(reg_q772 AND symb_decoder(16#7a#)) OR
 					(reg_q772 AND symb_decoder(16#5f#)) OR
 					(reg_q772 AND symb_decoder(16#df#)) OR
 					(reg_q772 AND symb_decoder(16#d0#)) OR
 					(reg_q772 AND symb_decoder(16#2c#)) OR
 					(reg_q772 AND symb_decoder(16#b0#)) OR
 					(reg_q772 AND symb_decoder(16#8f#)) OR
 					(reg_q772 AND symb_decoder(16#55#)) OR
 					(reg_q772 AND symb_decoder(16#c2#)) OR
 					(reg_q772 AND symb_decoder(16#f7#)) OR
 					(reg_q772 AND symb_decoder(16#d9#)) OR
 					(reg_q772 AND symb_decoder(16#5b#)) OR
 					(reg_q772 AND symb_decoder(16#ac#)) OR
 					(reg_q772 AND symb_decoder(16#2b#)) OR
 					(reg_q772 AND symb_decoder(16#40#)) OR
 					(reg_q772 AND symb_decoder(16#4b#)) OR
 					(reg_q772 AND symb_decoder(16#34#)) OR
 					(reg_q772 AND symb_decoder(16#89#)) OR
 					(reg_q772 AND symb_decoder(16#45#)) OR
 					(reg_q772 AND symb_decoder(16#c9#)) OR
 					(reg_q772 AND symb_decoder(16#ad#)) OR
 					(reg_q772 AND symb_decoder(16#ef#)) OR
 					(reg_q772 AND symb_decoder(16#5a#)) OR
 					(reg_q772 AND symb_decoder(16#83#)) OR
 					(reg_q772 AND symb_decoder(16#8e#)) OR
 					(reg_q772 AND symb_decoder(16#00#)) OR
 					(reg_q772 AND symb_decoder(16#16#)) OR
 					(reg_q772 AND symb_decoder(16#72#)) OR
 					(reg_q772 AND symb_decoder(16#a0#)) OR
 					(reg_q772 AND symb_decoder(16#9c#)) OR
 					(reg_q772 AND symb_decoder(16#ed#)) OR
 					(reg_q772 AND symb_decoder(16#2f#)) OR
 					(reg_q772 AND symb_decoder(16#39#)) OR
 					(reg_q772 AND symb_decoder(16#2d#)) OR
 					(reg_q772 AND symb_decoder(16#19#)) OR
 					(reg_q772 AND symb_decoder(16#21#)) OR
 					(reg_q772 AND symb_decoder(16#77#)) OR
 					(reg_q772 AND symb_decoder(16#04#)) OR
 					(reg_q772 AND symb_decoder(16#e9#)) OR
 					(reg_q772 AND symb_decoder(16#ca#)) OR
 					(reg_q772 AND symb_decoder(16#3f#)) OR
 					(reg_q772 AND symb_decoder(16#90#)) OR
 					(reg_q772 AND symb_decoder(16#33#)) OR
 					(reg_q772 AND symb_decoder(16#bf#)) OR
 					(reg_q772 AND symb_decoder(16#57#)) OR
 					(reg_q772 AND symb_decoder(16#8b#)) OR
 					(reg_q772 AND symb_decoder(16#d1#)) OR
 					(reg_q772 AND symb_decoder(16#e6#)) OR
 					(reg_q772 AND symb_decoder(16#fa#)) OR
 					(reg_q772 AND symb_decoder(16#01#)) OR
 					(reg_q772 AND symb_decoder(16#c8#)) OR
 					(reg_q772 AND symb_decoder(16#b4#)) OR
 					(reg_q772 AND symb_decoder(16#49#)) OR
 					(reg_q772 AND symb_decoder(16#1e#)) OR
 					(reg_q772 AND symb_decoder(16#eb#)) OR
 					(reg_q772 AND symb_decoder(16#f9#)) OR
 					(reg_q772 AND symb_decoder(16#79#)) OR
 					(reg_q772 AND symb_decoder(16#dc#)) OR
 					(reg_q772 AND symb_decoder(16#c6#)) OR
 					(reg_q772 AND symb_decoder(16#e7#)) OR
 					(reg_q772 AND symb_decoder(16#0a#)) OR
 					(reg_q772 AND symb_decoder(16#5c#)) OR
 					(reg_q772 AND symb_decoder(16#38#)) OR
 					(reg_q772 AND symb_decoder(16#f4#)) OR
 					(reg_q772 AND symb_decoder(16#0e#)) OR
 					(reg_q772 AND symb_decoder(16#1a#)) OR
 					(reg_q772 AND symb_decoder(16#82#)) OR
 					(reg_q772 AND symb_decoder(16#25#)) OR
 					(reg_q772 AND symb_decoder(16#6c#)) OR
 					(reg_q772 AND symb_decoder(16#7d#)) OR
 					(reg_q772 AND symb_decoder(16#61#)) OR
 					(reg_q772 AND symb_decoder(16#6a#)) OR
 					(reg_q772 AND symb_decoder(16#6f#)) OR
 					(reg_q772 AND symb_decoder(16#a9#)) OR
 					(reg_q772 AND symb_decoder(16#a4#)) OR
 					(reg_q772 AND symb_decoder(16#67#)) OR
 					(reg_q772 AND symb_decoder(16#58#)) OR
 					(reg_q772 AND symb_decoder(16#cb#)) OR
 					(reg_q772 AND symb_decoder(16#af#)) OR
 					(reg_q772 AND symb_decoder(16#63#)) OR
 					(reg_q772 AND symb_decoder(16#3d#)) OR
 					(reg_q772 AND symb_decoder(16#0c#)) OR
 					(reg_q772 AND symb_decoder(16#e1#)) OR
 					(reg_q772 AND symb_decoder(16#10#)) OR
 					(reg_q772 AND symb_decoder(16#f8#)) OR
 					(reg_q772 AND symb_decoder(16#02#)) OR
 					(reg_q772 AND symb_decoder(16#46#)) OR
 					(reg_q772 AND symb_decoder(16#12#)) OR
 					(reg_q772 AND symb_decoder(16#11#)) OR
 					(reg_q772 AND symb_decoder(16#d5#)) OR
 					(reg_q772 AND symb_decoder(16#b9#)) OR
 					(reg_q772 AND symb_decoder(16#0f#)) OR
 					(reg_q772 AND symb_decoder(16#8c#)) OR
 					(reg_q772 AND symb_decoder(16#cf#)) OR
 					(reg_q772 AND symb_decoder(16#ea#)) OR
 					(reg_q772 AND symb_decoder(16#44#)) OR
 					(reg_q772 AND symb_decoder(16#f0#)) OR
 					(reg_q772 AND symb_decoder(16#1f#)) OR
 					(reg_q772 AND symb_decoder(16#d2#)) OR
 					(reg_q772 AND symb_decoder(16#7b#)) OR
 					(reg_q772 AND symb_decoder(16#35#)) OR
 					(reg_q772 AND symb_decoder(16#73#)) OR
 					(reg_q772 AND symb_decoder(16#70#)) OR
 					(reg_q772 AND symb_decoder(16#a7#)) OR
 					(reg_q772 AND symb_decoder(16#de#)) OR
 					(reg_q772 AND symb_decoder(16#98#)) OR
 					(reg_q772 AND symb_decoder(16#3b#)) OR
 					(reg_q772 AND symb_decoder(16#9f#)) OR
 					(reg_q772 AND symb_decoder(16#9b#)) OR
 					(reg_q772 AND symb_decoder(16#41#)) OR
 					(reg_q772 AND symb_decoder(16#74#)) OR
 					(reg_q772 AND symb_decoder(16#43#)) OR
 					(reg_q772 AND symb_decoder(16#22#)) OR
 					(reg_q772 AND symb_decoder(16#f2#)) OR
 					(reg_q772 AND symb_decoder(16#a8#)) OR
 					(reg_q772 AND symb_decoder(16#b8#)) OR
 					(reg_q772 AND symb_decoder(16#30#)) OR
 					(reg_q772 AND symb_decoder(16#9a#)) OR
 					(reg_q772 AND symb_decoder(16#aa#)) OR
 					(reg_q772 AND symb_decoder(16#96#)) OR
 					(reg_q772 AND symb_decoder(16#ce#)) OR
 					(reg_q772 AND symb_decoder(16#dd#)) OR
 					(reg_q772 AND symb_decoder(16#c3#)) OR
 					(reg_q772 AND symb_decoder(16#bc#)) OR
 					(reg_q772 AND symb_decoder(16#7e#)) OR
 					(reg_q772 AND symb_decoder(16#0d#)) OR
 					(reg_q772 AND symb_decoder(16#d4#)) OR
 					(reg_q772 AND symb_decoder(16#ee#)) OR
 					(reg_q772 AND symb_decoder(16#b3#)) OR
 					(reg_q772 AND symb_decoder(16#37#)) OR
 					(reg_q772 AND symb_decoder(16#95#)) OR
 					(reg_q772 AND symb_decoder(16#b2#)) OR
 					(reg_q772 AND symb_decoder(16#18#)) OR
 					(reg_q772 AND symb_decoder(16#6e#)) OR
 					(reg_q772 AND symb_decoder(16#b7#)) OR
 					(reg_q772 AND symb_decoder(16#db#)) OR
 					(reg_q772 AND symb_decoder(16#65#)) OR
 					(reg_q772 AND symb_decoder(16#ec#)) OR
 					(reg_q772 AND symb_decoder(16#a6#)) OR
 					(reg_q772 AND symb_decoder(16#b5#)) OR
 					(reg_q772 AND symb_decoder(16#36#)) OR
 					(reg_q772 AND symb_decoder(16#68#)) OR
 					(reg_q772 AND symb_decoder(16#2a#)) OR
 					(reg_q772 AND symb_decoder(16#c5#)) OR
 					(reg_q772 AND symb_decoder(16#fe#)) OR
 					(reg_q772 AND symb_decoder(16#06#)) OR
 					(reg_q772 AND symb_decoder(16#3a#)) OR
 					(reg_q772 AND symb_decoder(16#d3#)) OR
 					(reg_q772 AND symb_decoder(16#3c#)) OR
 					(reg_q772 AND symb_decoder(16#91#)) OR
 					(reg_q772 AND symb_decoder(16#3e#)) OR
 					(reg_q772 AND symb_decoder(16#f5#)) OR
 					(reg_q772 AND symb_decoder(16#e2#)) OR
 					(reg_q772 AND symb_decoder(16#1c#)) OR
 					(reg_q772 AND symb_decoder(16#86#)) OR
 					(reg_q772 AND symb_decoder(16#d6#)) OR
 					(reg_q772 AND symb_decoder(16#be#)) OR
 					(reg_q772 AND symb_decoder(16#f3#)) OR
 					(reg_q772 AND symb_decoder(16#ae#)) OR
 					(reg_q772 AND symb_decoder(16#a3#)) OR
 					(reg_q772 AND symb_decoder(16#1d#)) OR
 					(reg_q772 AND symb_decoder(16#f6#)) OR
 					(reg_q772 AND symb_decoder(16#fb#)) OR
 					(reg_q772 AND symb_decoder(16#92#)) OR
 					(reg_q772 AND symb_decoder(16#78#)) OR
 					(reg_q772 AND symb_decoder(16#59#)) OR
 					(reg_q772 AND symb_decoder(16#1b#)) OR
 					(reg_q772 AND symb_decoder(16#a1#)) OR
 					(reg_q772 AND symb_decoder(16#6b#)) OR
 					(reg_q772 AND symb_decoder(16#fc#)) OR
 					(reg_q772 AND symb_decoder(16#05#)) OR
 					(reg_q772 AND symb_decoder(16#6d#)) OR
 					(reg_q772 AND symb_decoder(16#42#)) OR
 					(reg_q772 AND symb_decoder(16#54#)) OR
 					(reg_q772 AND symb_decoder(16#71#)) OR
 					(reg_q772 AND symb_decoder(16#b1#)) OR
 					(reg_q772 AND symb_decoder(16#75#)) OR
 					(reg_q772 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#));
reg_q772_init <= '0' ;
	p_reg_q772: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q772 <= reg_q772_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q772 <= reg_q772_init;
        else
          reg_q772 <= reg_q772_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q590_in <= (reg_q590 AND symb_decoder(16#a7#)) OR
 					(reg_q590 AND symb_decoder(16#7e#)) OR
 					(reg_q590 AND symb_decoder(16#1f#)) OR
 					(reg_q590 AND symb_decoder(16#86#)) OR
 					(reg_q590 AND symb_decoder(16#1c#)) OR
 					(reg_q590 AND symb_decoder(16#14#)) OR
 					(reg_q590 AND symb_decoder(16#7a#)) OR
 					(reg_q590 AND symb_decoder(16#8f#)) OR
 					(reg_q590 AND symb_decoder(16#2a#)) OR
 					(reg_q590 AND symb_decoder(16#97#)) OR
 					(reg_q590 AND symb_decoder(16#1b#)) OR
 					(reg_q590 AND symb_decoder(16#e3#)) OR
 					(reg_q590 AND symb_decoder(16#5f#)) OR
 					(reg_q590 AND symb_decoder(16#9c#)) OR
 					(reg_q590 AND symb_decoder(16#58#)) OR
 					(reg_q590 AND symb_decoder(16#e0#)) OR
 					(reg_q590 AND symb_decoder(16#71#)) OR
 					(reg_q590 AND symb_decoder(16#8d#)) OR
 					(reg_q590 AND symb_decoder(16#20#)) OR
 					(reg_q590 AND symb_decoder(16#3b#)) OR
 					(reg_q590 AND symb_decoder(16#32#)) OR
 					(reg_q590 AND symb_decoder(16#ed#)) OR
 					(reg_q590 AND symb_decoder(16#bd#)) OR
 					(reg_q590 AND symb_decoder(16#1a#)) OR
 					(reg_q590 AND symb_decoder(16#4a#)) OR
 					(reg_q590 AND symb_decoder(16#ac#)) OR
 					(reg_q590 AND symb_decoder(16#6e#)) OR
 					(reg_q590 AND symb_decoder(16#e8#)) OR
 					(reg_q590 AND symb_decoder(16#74#)) OR
 					(reg_q590 AND symb_decoder(16#f5#)) OR
 					(reg_q590 AND symb_decoder(16#2f#)) OR
 					(reg_q590 AND symb_decoder(16#02#)) OR
 					(reg_q590 AND symb_decoder(16#67#)) OR
 					(reg_q590 AND symb_decoder(16#17#)) OR
 					(reg_q590 AND symb_decoder(16#91#)) OR
 					(reg_q590 AND symb_decoder(16#fe#)) OR
 					(reg_q590 AND symb_decoder(16#77#)) OR
 					(reg_q590 AND symb_decoder(16#0c#)) OR
 					(reg_q590 AND symb_decoder(16#72#)) OR
 					(reg_q590 AND symb_decoder(16#69#)) OR
 					(reg_q590 AND symb_decoder(16#90#)) OR
 					(reg_q590 AND symb_decoder(16#46#)) OR
 					(reg_q590 AND symb_decoder(16#6d#)) OR
 					(reg_q590 AND symb_decoder(16#82#)) OR
 					(reg_q590 AND symb_decoder(16#fd#)) OR
 					(reg_q590 AND symb_decoder(16#16#)) OR
 					(reg_q590 AND symb_decoder(16#6b#)) OR
 					(reg_q590 AND symb_decoder(16#ce#)) OR
 					(reg_q590 AND symb_decoder(16#88#)) OR
 					(reg_q590 AND symb_decoder(16#0f#)) OR
 					(reg_q590 AND symb_decoder(16#d1#)) OR
 					(reg_q590 AND symb_decoder(16#b7#)) OR
 					(reg_q590 AND symb_decoder(16#03#)) OR
 					(reg_q590 AND symb_decoder(16#e6#)) OR
 					(reg_q590 AND symb_decoder(16#c8#)) OR
 					(reg_q590 AND symb_decoder(16#54#)) OR
 					(reg_q590 AND symb_decoder(16#2c#)) OR
 					(reg_q590 AND symb_decoder(16#4d#)) OR
 					(reg_q590 AND symb_decoder(16#3d#)) OR
 					(reg_q590 AND symb_decoder(16#c1#)) OR
 					(reg_q590 AND symb_decoder(16#ec#)) OR
 					(reg_q590 AND symb_decoder(16#6f#)) OR
 					(reg_q590 AND symb_decoder(16#a3#)) OR
 					(reg_q590 AND symb_decoder(16#4f#)) OR
 					(reg_q590 AND symb_decoder(16#76#)) OR
 					(reg_q590 AND symb_decoder(16#ea#)) OR
 					(reg_q590 AND symb_decoder(16#8e#)) OR
 					(reg_q590 AND symb_decoder(16#95#)) OR
 					(reg_q590 AND symb_decoder(16#3e#)) OR
 					(reg_q590 AND symb_decoder(16#65#)) OR
 					(reg_q590 AND symb_decoder(16#e7#)) OR
 					(reg_q590 AND symb_decoder(16#62#)) OR
 					(reg_q590 AND symb_decoder(16#9d#)) OR
 					(reg_q590 AND symb_decoder(16#e9#)) OR
 					(reg_q590 AND symb_decoder(16#fc#)) OR
 					(reg_q590 AND symb_decoder(16#96#)) OR
 					(reg_q590 AND symb_decoder(16#48#)) OR
 					(reg_q590 AND symb_decoder(16#49#)) OR
 					(reg_q590 AND symb_decoder(16#b5#)) OR
 					(reg_q590 AND symb_decoder(16#9b#)) OR
 					(reg_q590 AND symb_decoder(16#05#)) OR
 					(reg_q590 AND symb_decoder(16#c7#)) OR
 					(reg_q590 AND symb_decoder(16#73#)) OR
 					(reg_q590 AND symb_decoder(16#d5#)) OR
 					(reg_q590 AND symb_decoder(16#a4#)) OR
 					(reg_q590 AND symb_decoder(16#26#)) OR
 					(reg_q590 AND symb_decoder(16#22#)) OR
 					(reg_q590 AND symb_decoder(16#61#)) OR
 					(reg_q590 AND symb_decoder(16#ef#)) OR
 					(reg_q590 AND symb_decoder(16#b0#)) OR
 					(reg_q590 AND symb_decoder(16#5d#)) OR
 					(reg_q590 AND symb_decoder(16#ae#)) OR
 					(reg_q590 AND symb_decoder(16#9f#)) OR
 					(reg_q590 AND symb_decoder(16#37#)) OR
 					(reg_q590 AND symb_decoder(16#09#)) OR
 					(reg_q590 AND symb_decoder(16#83#)) OR
 					(reg_q590 AND symb_decoder(16#ab#)) OR
 					(reg_q590 AND symb_decoder(16#af#)) OR
 					(reg_q590 AND symb_decoder(16#34#)) OR
 					(reg_q590 AND symb_decoder(16#60#)) OR
 					(reg_q590 AND symb_decoder(16#d9#)) OR
 					(reg_q590 AND symb_decoder(16#be#)) OR
 					(reg_q590 AND symb_decoder(16#93#)) OR
 					(reg_q590 AND symb_decoder(16#41#)) OR
 					(reg_q590 AND symb_decoder(16#2d#)) OR
 					(reg_q590 AND symb_decoder(16#c6#)) OR
 					(reg_q590 AND symb_decoder(16#92#)) OR
 					(reg_q590 AND symb_decoder(16#75#)) OR
 					(reg_q590 AND symb_decoder(16#a1#)) OR
 					(reg_q590 AND symb_decoder(16#fa#)) OR
 					(reg_q590 AND symb_decoder(16#ff#)) OR
 					(reg_q590 AND symb_decoder(16#25#)) OR
 					(reg_q590 AND symb_decoder(16#b4#)) OR
 					(reg_q590 AND symb_decoder(16#cb#)) OR
 					(reg_q590 AND symb_decoder(16#5a#)) OR
 					(reg_q590 AND symb_decoder(16#31#)) OR
 					(reg_q590 AND symb_decoder(16#44#)) OR
 					(reg_q590 AND symb_decoder(16#45#)) OR
 					(reg_q590 AND symb_decoder(16#1e#)) OR
 					(reg_q590 AND symb_decoder(16#9e#)) OR
 					(reg_q590 AND symb_decoder(16#79#)) OR
 					(reg_q590 AND symb_decoder(16#f8#)) OR
 					(reg_q590 AND symb_decoder(16#43#)) OR
 					(reg_q590 AND symb_decoder(16#00#)) OR
 					(reg_q590 AND symb_decoder(16#55#)) OR
 					(reg_q590 AND symb_decoder(16#66#)) OR
 					(reg_q590 AND symb_decoder(16#f6#)) OR
 					(reg_q590 AND symb_decoder(16#f2#)) OR
 					(reg_q590 AND symb_decoder(16#11#)) OR
 					(reg_q590 AND symb_decoder(16#db#)) OR
 					(reg_q590 AND symb_decoder(16#52#)) OR
 					(reg_q590 AND symb_decoder(16#d8#)) OR
 					(reg_q590 AND symb_decoder(16#2b#)) OR
 					(reg_q590 AND symb_decoder(16#e4#)) OR
 					(reg_q590 AND symb_decoder(16#b2#)) OR
 					(reg_q590 AND symb_decoder(16#50#)) OR
 					(reg_q590 AND symb_decoder(16#5c#)) OR
 					(reg_q590 AND symb_decoder(16#0e#)) OR
 					(reg_q590 AND symb_decoder(16#c0#)) OR
 					(reg_q590 AND symb_decoder(16#d7#)) OR
 					(reg_q590 AND symb_decoder(16#ba#)) OR
 					(reg_q590 AND symb_decoder(16#cc#)) OR
 					(reg_q590 AND symb_decoder(16#f9#)) OR
 					(reg_q590 AND symb_decoder(16#94#)) OR
 					(reg_q590 AND symb_decoder(16#5e#)) OR
 					(reg_q590 AND symb_decoder(16#aa#)) OR
 					(reg_q590 AND symb_decoder(16#0a#)) OR
 					(reg_q590 AND symb_decoder(16#8b#)) OR
 					(reg_q590 AND symb_decoder(16#8a#)) OR
 					(reg_q590 AND symb_decoder(16#3a#)) OR
 					(reg_q590 AND symb_decoder(16#63#)) OR
 					(reg_q590 AND symb_decoder(16#15#)) OR
 					(reg_q590 AND symb_decoder(16#bc#)) OR
 					(reg_q590 AND symb_decoder(16#a6#)) OR
 					(reg_q590 AND symb_decoder(16#d0#)) OR
 					(reg_q590 AND symb_decoder(16#a2#)) OR
 					(reg_q590 AND symb_decoder(16#a0#)) OR
 					(reg_q590 AND symb_decoder(16#78#)) OR
 					(reg_q590 AND symb_decoder(16#57#)) OR
 					(reg_q590 AND symb_decoder(16#dc#)) OR
 					(reg_q590 AND symb_decoder(16#c3#)) OR
 					(reg_q590 AND symb_decoder(16#cd#)) OR
 					(reg_q590 AND symb_decoder(16#81#)) OR
 					(reg_q590 AND symb_decoder(16#b3#)) OR
 					(reg_q590 AND symb_decoder(16#de#)) OR
 					(reg_q590 AND symb_decoder(16#0d#)) OR
 					(reg_q590 AND symb_decoder(16#51#)) OR
 					(reg_q590 AND symb_decoder(16#4e#)) OR
 					(reg_q590 AND symb_decoder(16#df#)) OR
 					(reg_q590 AND symb_decoder(16#68#)) OR
 					(reg_q590 AND symb_decoder(16#ad#)) OR
 					(reg_q590 AND symb_decoder(16#0b#)) OR
 					(reg_q590 AND symb_decoder(16#7d#)) OR
 					(reg_q590 AND symb_decoder(16#98#)) OR
 					(reg_q590 AND symb_decoder(16#19#)) OR
 					(reg_q590 AND symb_decoder(16#47#)) OR
 					(reg_q590 AND symb_decoder(16#bf#)) OR
 					(reg_q590 AND symb_decoder(16#40#)) OR
 					(reg_q590 AND symb_decoder(16#a8#)) OR
 					(reg_q590 AND symb_decoder(16#21#)) OR
 					(reg_q590 AND symb_decoder(16#13#)) OR
 					(reg_q590 AND symb_decoder(16#64#)) OR
 					(reg_q590 AND symb_decoder(16#85#)) OR
 					(reg_q590 AND symb_decoder(16#35#)) OR
 					(reg_q590 AND symb_decoder(16#e1#)) OR
 					(reg_q590 AND symb_decoder(16#3c#)) OR
 					(reg_q590 AND symb_decoder(16#b8#)) OR
 					(reg_q590 AND symb_decoder(16#b9#)) OR
 					(reg_q590 AND symb_decoder(16#8c#)) OR
 					(reg_q590 AND symb_decoder(16#c4#)) OR
 					(reg_q590 AND symb_decoder(16#c2#)) OR
 					(reg_q590 AND symb_decoder(16#5b#)) OR
 					(reg_q590 AND symb_decoder(16#53#)) OR
 					(reg_q590 AND symb_decoder(16#c5#)) OR
 					(reg_q590 AND symb_decoder(16#08#)) OR
 					(reg_q590 AND symb_decoder(16#6c#)) OR
 					(reg_q590 AND symb_decoder(16#27#)) OR
 					(reg_q590 AND symb_decoder(16#06#)) OR
 					(reg_q590 AND symb_decoder(16#99#)) OR
 					(reg_q590 AND symb_decoder(16#84#)) OR
 					(reg_q590 AND symb_decoder(16#39#)) OR
 					(reg_q590 AND symb_decoder(16#f7#)) OR
 					(reg_q590 AND symb_decoder(16#3f#)) OR
 					(reg_q590 AND symb_decoder(16#b1#)) OR
 					(reg_q590 AND symb_decoder(16#f1#)) OR
 					(reg_q590 AND symb_decoder(16#2e#)) OR
 					(reg_q590 AND symb_decoder(16#70#)) OR
 					(reg_q590 AND symb_decoder(16#12#)) OR
 					(reg_q590 AND symb_decoder(16#07#)) OR
 					(reg_q590 AND symb_decoder(16#e5#)) OR
 					(reg_q590 AND symb_decoder(16#7f#)) OR
 					(reg_q590 AND symb_decoder(16#24#)) OR
 					(reg_q590 AND symb_decoder(16#f4#)) OR
 					(reg_q590 AND symb_decoder(16#d3#)) OR
 					(reg_q590 AND symb_decoder(16#33#)) OR
 					(reg_q590 AND symb_decoder(16#bb#)) OR
 					(reg_q590 AND symb_decoder(16#04#)) OR
 					(reg_q590 AND symb_decoder(16#f3#)) OR
 					(reg_q590 AND symb_decoder(16#23#)) OR
 					(reg_q590 AND symb_decoder(16#fb#)) OR
 					(reg_q590 AND symb_decoder(16#d6#)) OR
 					(reg_q590 AND symb_decoder(16#f0#)) OR
 					(reg_q590 AND symb_decoder(16#89#)) OR
 					(reg_q590 AND symb_decoder(16#56#)) OR
 					(reg_q590 AND symb_decoder(16#dd#)) OR
 					(reg_q590 AND symb_decoder(16#ee#)) OR
 					(reg_q590 AND symb_decoder(16#eb#)) OR
 					(reg_q590 AND symb_decoder(16#ca#)) OR
 					(reg_q590 AND symb_decoder(16#01#)) OR
 					(reg_q590 AND symb_decoder(16#d4#)) OR
 					(reg_q590 AND symb_decoder(16#10#)) OR
 					(reg_q590 AND symb_decoder(16#7c#)) OR
 					(reg_q590 AND symb_decoder(16#42#)) OR
 					(reg_q590 AND symb_decoder(16#28#)) OR
 					(reg_q590 AND symb_decoder(16#e2#)) OR
 					(reg_q590 AND symb_decoder(16#29#)) OR
 					(reg_q590 AND symb_decoder(16#80#)) OR
 					(reg_q590 AND symb_decoder(16#cf#)) OR
 					(reg_q590 AND symb_decoder(16#9a#)) OR
 					(reg_q590 AND symb_decoder(16#18#)) OR
 					(reg_q590 AND symb_decoder(16#36#)) OR
 					(reg_q590 AND symb_decoder(16#4b#)) OR
 					(reg_q590 AND symb_decoder(16#4c#)) OR
 					(reg_q590 AND symb_decoder(16#1d#)) OR
 					(reg_q590 AND symb_decoder(16#d2#)) OR
 					(reg_q590 AND symb_decoder(16#7b#)) OR
 					(reg_q590 AND symb_decoder(16#a5#)) OR
 					(reg_q590 AND symb_decoder(16#c9#)) OR
 					(reg_q590 AND symb_decoder(16#6a#)) OR
 					(reg_q590 AND symb_decoder(16#a9#)) OR
 					(reg_q590 AND symb_decoder(16#b6#)) OR
 					(reg_q590 AND symb_decoder(16#59#)) OR
 					(reg_q590 AND symb_decoder(16#da#)) OR
 					(reg_q590 AND symb_decoder(16#38#)) OR
 					(reg_q590 AND symb_decoder(16#87#)) OR
 					(reg_q590 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#));
reg_q590_init <= '0' ;
	p_reg_q590: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q590 <= reg_q590_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q590 <= reg_q590_init;
        else
          reg_q590 <= reg_q590_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q545_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q545 AND symb_decoder(16#93#)) OR
 					(reg_q545 AND symb_decoder(16#d3#)) OR
 					(reg_q545 AND symb_decoder(16#8a#)) OR
 					(reg_q545 AND symb_decoder(16#b2#)) OR
 					(reg_q545 AND symb_decoder(16#ad#)) OR
 					(reg_q545 AND symb_decoder(16#69#)) OR
 					(reg_q545 AND symb_decoder(16#0c#)) OR
 					(reg_q545 AND symb_decoder(16#64#)) OR
 					(reg_q545 AND symb_decoder(16#00#)) OR
 					(reg_q545 AND symb_decoder(16#e4#)) OR
 					(reg_q545 AND symb_decoder(16#dd#)) OR
 					(reg_q545 AND symb_decoder(16#7b#)) OR
 					(reg_q545 AND symb_decoder(16#ca#)) OR
 					(reg_q545 AND symb_decoder(16#89#)) OR
 					(reg_q545 AND symb_decoder(16#24#)) OR
 					(reg_q545 AND symb_decoder(16#7c#)) OR
 					(reg_q545 AND symb_decoder(16#60#)) OR
 					(reg_q545 AND symb_decoder(16#0d#)) OR
 					(reg_q545 AND symb_decoder(16#c1#)) OR
 					(reg_q545 AND symb_decoder(16#de#)) OR
 					(reg_q545 AND symb_decoder(16#95#)) OR
 					(reg_q545 AND symb_decoder(16#8b#)) OR
 					(reg_q545 AND symb_decoder(16#c0#)) OR
 					(reg_q545 AND symb_decoder(16#81#)) OR
 					(reg_q545 AND symb_decoder(16#aa#)) OR
 					(reg_q545 AND symb_decoder(16#a1#)) OR
 					(reg_q545 AND symb_decoder(16#91#)) OR
 					(reg_q545 AND symb_decoder(16#d6#)) OR
 					(reg_q545 AND symb_decoder(16#a4#)) OR
 					(reg_q545 AND symb_decoder(16#fe#)) OR
 					(reg_q545 AND symb_decoder(16#18#)) OR
 					(reg_q545 AND symb_decoder(16#67#)) OR
 					(reg_q545 AND symb_decoder(16#dc#)) OR
 					(reg_q545 AND symb_decoder(16#40#)) OR
 					(reg_q545 AND symb_decoder(16#b8#)) OR
 					(reg_q545 AND symb_decoder(16#0f#)) OR
 					(reg_q545 AND symb_decoder(16#e0#)) OR
 					(reg_q545 AND symb_decoder(16#c7#)) OR
 					(reg_q545 AND symb_decoder(16#30#)) OR
 					(reg_q545 AND symb_decoder(16#29#)) OR
 					(reg_q545 AND symb_decoder(16#cc#)) OR
 					(reg_q545 AND symb_decoder(16#88#)) OR
 					(reg_q545 AND symb_decoder(16#96#)) OR
 					(reg_q545 AND symb_decoder(16#0e#)) OR
 					(reg_q545 AND symb_decoder(16#7f#)) OR
 					(reg_q545 AND symb_decoder(16#5d#)) OR
 					(reg_q545 AND symb_decoder(16#f1#)) OR
 					(reg_q545 AND symb_decoder(16#63#)) OR
 					(reg_q545 AND symb_decoder(16#d1#)) OR
 					(reg_q545 AND symb_decoder(16#ec#)) OR
 					(reg_q545 AND symb_decoder(16#56#)) OR
 					(reg_q545 AND symb_decoder(16#66#)) OR
 					(reg_q545 AND symb_decoder(16#84#)) OR
 					(reg_q545 AND symb_decoder(16#31#)) OR
 					(reg_q545 AND symb_decoder(16#e5#)) OR
 					(reg_q545 AND symb_decoder(16#45#)) OR
 					(reg_q545 AND symb_decoder(16#b0#)) OR
 					(reg_q545 AND symb_decoder(16#a6#)) OR
 					(reg_q545 AND symb_decoder(16#8c#)) OR
 					(reg_q545 AND symb_decoder(16#b4#)) OR
 					(reg_q545 AND symb_decoder(16#ee#)) OR
 					(reg_q545 AND symb_decoder(16#3b#)) OR
 					(reg_q545 AND symb_decoder(16#ff#)) OR
 					(reg_q545 AND symb_decoder(16#61#)) OR
 					(reg_q545 AND symb_decoder(16#80#)) OR
 					(reg_q545 AND symb_decoder(16#ae#)) OR
 					(reg_q545 AND symb_decoder(16#11#)) OR
 					(reg_q545 AND symb_decoder(16#0b#)) OR
 					(reg_q545 AND symb_decoder(16#be#)) OR
 					(reg_q545 AND symb_decoder(16#1f#)) OR
 					(reg_q545 AND symb_decoder(16#49#)) OR
 					(reg_q545 AND symb_decoder(16#d7#)) OR
 					(reg_q545 AND symb_decoder(16#3c#)) OR
 					(reg_q545 AND symb_decoder(16#e2#)) OR
 					(reg_q545 AND symb_decoder(16#85#)) OR
 					(reg_q545 AND symb_decoder(16#1d#)) OR
 					(reg_q545 AND symb_decoder(16#52#)) OR
 					(reg_q545 AND symb_decoder(16#fb#)) OR
 					(reg_q545 AND symb_decoder(16#c4#)) OR
 					(reg_q545 AND symb_decoder(16#87#)) OR
 					(reg_q545 AND symb_decoder(16#bb#)) OR
 					(reg_q545 AND symb_decoder(16#1b#)) OR
 					(reg_q545 AND symb_decoder(16#44#)) OR
 					(reg_q545 AND symb_decoder(16#f4#)) OR
 					(reg_q545 AND symb_decoder(16#15#)) OR
 					(reg_q545 AND symb_decoder(16#5f#)) OR
 					(reg_q545 AND symb_decoder(16#c2#)) OR
 					(reg_q545 AND symb_decoder(16#6b#)) OR
 					(reg_q545 AND symb_decoder(16#6f#)) OR
 					(reg_q545 AND symb_decoder(16#eb#)) OR
 					(reg_q545 AND symb_decoder(16#26#)) OR
 					(reg_q545 AND symb_decoder(16#9d#)) OR
 					(reg_q545 AND symb_decoder(16#75#)) OR
 					(reg_q545 AND symb_decoder(16#99#)) OR
 					(reg_q545 AND symb_decoder(16#f0#)) OR
 					(reg_q545 AND symb_decoder(16#51#)) OR
 					(reg_q545 AND symb_decoder(16#ea#)) OR
 					(reg_q545 AND symb_decoder(16#cb#)) OR
 					(reg_q545 AND symb_decoder(16#05#)) OR
 					(reg_q545 AND symb_decoder(16#07#)) OR
 					(reg_q545 AND symb_decoder(16#b6#)) OR
 					(reg_q545 AND symb_decoder(16#d2#)) OR
 					(reg_q545 AND symb_decoder(16#53#)) OR
 					(reg_q545 AND symb_decoder(16#50#)) OR
 					(reg_q545 AND symb_decoder(16#f6#)) OR
 					(reg_q545 AND symb_decoder(16#65#)) OR
 					(reg_q545 AND symb_decoder(16#2b#)) OR
 					(reg_q545 AND symb_decoder(16#34#)) OR
 					(reg_q545 AND symb_decoder(16#a7#)) OR
 					(reg_q545 AND symb_decoder(16#3d#)) OR
 					(reg_q545 AND symb_decoder(16#6a#)) OR
 					(reg_q545 AND symb_decoder(16#6c#)) OR
 					(reg_q545 AND symb_decoder(16#5e#)) OR
 					(reg_q545 AND symb_decoder(16#21#)) OR
 					(reg_q545 AND symb_decoder(16#b3#)) OR
 					(reg_q545 AND symb_decoder(16#02#)) OR
 					(reg_q545 AND symb_decoder(16#0a#)) OR
 					(reg_q545 AND symb_decoder(16#94#)) OR
 					(reg_q545 AND symb_decoder(16#f5#)) OR
 					(reg_q545 AND symb_decoder(16#b5#)) OR
 					(reg_q545 AND symb_decoder(16#d4#)) OR
 					(reg_q545 AND symb_decoder(16#17#)) OR
 					(reg_q545 AND symb_decoder(16#82#)) OR
 					(reg_q545 AND symb_decoder(16#22#)) OR
 					(reg_q545 AND symb_decoder(16#47#)) OR
 					(reg_q545 AND symb_decoder(16#58#)) OR
 					(reg_q545 AND symb_decoder(16#f2#)) OR
 					(reg_q545 AND symb_decoder(16#16#)) OR
 					(reg_q545 AND symb_decoder(16#71#)) OR
 					(reg_q545 AND symb_decoder(16#10#)) OR
 					(reg_q545 AND symb_decoder(16#b1#)) OR
 					(reg_q545 AND symb_decoder(16#3f#)) OR
 					(reg_q545 AND symb_decoder(16#6d#)) OR
 					(reg_q545 AND symb_decoder(16#a2#)) OR
 					(reg_q545 AND symb_decoder(16#12#)) OR
 					(reg_q545 AND symb_decoder(16#9b#)) OR
 					(reg_q545 AND symb_decoder(16#3a#)) OR
 					(reg_q545 AND symb_decoder(16#5a#)) OR
 					(reg_q545 AND symb_decoder(16#59#)) OR
 					(reg_q545 AND symb_decoder(16#38#)) OR
 					(reg_q545 AND symb_decoder(16#28#)) OR
 					(reg_q545 AND symb_decoder(16#33#)) OR
 					(reg_q545 AND symb_decoder(16#08#)) OR
 					(reg_q545 AND symb_decoder(16#70#)) OR
 					(reg_q545 AND symb_decoder(16#2c#)) OR
 					(reg_q545 AND symb_decoder(16#43#)) OR
 					(reg_q545 AND symb_decoder(16#03#)) OR
 					(reg_q545 AND symb_decoder(16#4f#)) OR
 					(reg_q545 AND symb_decoder(16#4c#)) OR
 					(reg_q545 AND symb_decoder(16#4b#)) OR
 					(reg_q545 AND symb_decoder(16#1e#)) OR
 					(reg_q545 AND symb_decoder(16#c5#)) OR
 					(reg_q545 AND symb_decoder(16#a3#)) OR
 					(reg_q545 AND symb_decoder(16#09#)) OR
 					(reg_q545 AND symb_decoder(16#8e#)) OR
 					(reg_q545 AND symb_decoder(16#c9#)) OR
 					(reg_q545 AND symb_decoder(16#cf#)) OR
 					(reg_q545 AND symb_decoder(16#cd#)) OR
 					(reg_q545 AND symb_decoder(16#f8#)) OR
 					(reg_q545 AND symb_decoder(16#f7#)) OR
 					(reg_q545 AND symb_decoder(16#d8#)) OR
 					(reg_q545 AND symb_decoder(16#79#)) OR
 					(reg_q545 AND symb_decoder(16#57#)) OR
 					(reg_q545 AND symb_decoder(16#bc#)) OR
 					(reg_q545 AND symb_decoder(16#2e#)) OR
 					(reg_q545 AND symb_decoder(16#ed#)) OR
 					(reg_q545 AND symb_decoder(16#72#)) OR
 					(reg_q545 AND symb_decoder(16#83#)) OR
 					(reg_q545 AND symb_decoder(16#73#)) OR
 					(reg_q545 AND symb_decoder(16#d5#)) OR
 					(reg_q545 AND symb_decoder(16#8d#)) OR
 					(reg_q545 AND symb_decoder(16#41#)) OR
 					(reg_q545 AND symb_decoder(16#5c#)) OR
 					(reg_q545 AND symb_decoder(16#01#)) OR
 					(reg_q545 AND symb_decoder(16#14#)) OR
 					(reg_q545 AND symb_decoder(16#6e#)) OR
 					(reg_q545 AND symb_decoder(16#7e#)) OR
 					(reg_q545 AND symb_decoder(16#d9#)) OR
 					(reg_q545 AND symb_decoder(16#19#)) OR
 					(reg_q545 AND symb_decoder(16#a0#)) OR
 					(reg_q545 AND symb_decoder(16#04#)) OR
 					(reg_q545 AND symb_decoder(16#86#)) OR
 					(reg_q545 AND symb_decoder(16#68#)) OR
 					(reg_q545 AND symb_decoder(16#54#)) OR
 					(reg_q545 AND symb_decoder(16#da#)) OR
 					(reg_q545 AND symb_decoder(16#f3#)) OR
 					(reg_q545 AND symb_decoder(16#2f#)) OR
 					(reg_q545 AND symb_decoder(16#13#)) OR
 					(reg_q545 AND symb_decoder(16#ab#)) OR
 					(reg_q545 AND symb_decoder(16#4a#)) OR
 					(reg_q545 AND symb_decoder(16#e6#)) OR
 					(reg_q545 AND symb_decoder(16#1a#)) OR
 					(reg_q545 AND symb_decoder(16#35#)) OR
 					(reg_q545 AND symb_decoder(16#ce#)) OR
 					(reg_q545 AND symb_decoder(16#2d#)) OR
 					(reg_q545 AND symb_decoder(16#55#)) OR
 					(reg_q545 AND symb_decoder(16#af#)) OR
 					(reg_q545 AND symb_decoder(16#db#)) OR
 					(reg_q545 AND symb_decoder(16#9a#)) OR
 					(reg_q545 AND symb_decoder(16#98#)) OR
 					(reg_q545 AND symb_decoder(16#4d#)) OR
 					(reg_q545 AND symb_decoder(16#ac#)) OR
 					(reg_q545 AND symb_decoder(16#74#)) OR
 					(reg_q545 AND symb_decoder(16#20#)) OR
 					(reg_q545 AND symb_decoder(16#a8#)) OR
 					(reg_q545 AND symb_decoder(16#b7#)) OR
 					(reg_q545 AND symb_decoder(16#f9#)) OR
 					(reg_q545 AND symb_decoder(16#4e#)) OR
 					(reg_q545 AND symb_decoder(16#7a#)) OR
 					(reg_q545 AND symb_decoder(16#2a#)) OR
 					(reg_q545 AND symb_decoder(16#b9#)) OR
 					(reg_q545 AND symb_decoder(16#c8#)) OR
 					(reg_q545 AND symb_decoder(16#8f#)) OR
 					(reg_q545 AND symb_decoder(16#ef#)) OR
 					(reg_q545 AND symb_decoder(16#97#)) OR
 					(reg_q545 AND symb_decoder(16#c6#)) OR
 					(reg_q545 AND symb_decoder(16#42#)) OR
 					(reg_q545 AND symb_decoder(16#9e#)) OR
 					(reg_q545 AND symb_decoder(16#a5#)) OR
 					(reg_q545 AND symb_decoder(16#df#)) OR
 					(reg_q545 AND symb_decoder(16#1c#)) OR
 					(reg_q545 AND symb_decoder(16#78#)) OR
 					(reg_q545 AND symb_decoder(16#ba#)) OR
 					(reg_q545 AND symb_decoder(16#fa#)) OR
 					(reg_q545 AND symb_decoder(16#46#)) OR
 					(reg_q545 AND symb_decoder(16#5b#)) OR
 					(reg_q545 AND symb_decoder(16#32#)) OR
 					(reg_q545 AND symb_decoder(16#23#)) OR
 					(reg_q545 AND symb_decoder(16#e1#)) OR
 					(reg_q545 AND symb_decoder(16#c3#)) OR
 					(reg_q545 AND symb_decoder(16#3e#)) OR
 					(reg_q545 AND symb_decoder(16#76#)) OR
 					(reg_q545 AND symb_decoder(16#39#)) OR
 					(reg_q545 AND symb_decoder(16#9f#)) OR
 					(reg_q545 AND symb_decoder(16#06#)) OR
 					(reg_q545 AND symb_decoder(16#25#)) OR
 					(reg_q545 AND symb_decoder(16#77#)) OR
 					(reg_q545 AND symb_decoder(16#7d#)) OR
 					(reg_q545 AND symb_decoder(16#e7#)) OR
 					(reg_q545 AND symb_decoder(16#a9#)) OR
 					(reg_q545 AND symb_decoder(16#e9#)) OR
 					(reg_q545 AND symb_decoder(16#36#)) OR
 					(reg_q545 AND symb_decoder(16#fd#)) OR
 					(reg_q545 AND symb_decoder(16#9c#)) OR
 					(reg_q545 AND symb_decoder(16#37#)) OR
 					(reg_q545 AND symb_decoder(16#90#)) OR
 					(reg_q545 AND symb_decoder(16#fc#)) OR
 					(reg_q545 AND symb_decoder(16#92#)) OR
 					(reg_q545 AND symb_decoder(16#bd#)) OR
 					(reg_q545 AND symb_decoder(16#e8#)) OR
 					(reg_q545 AND symb_decoder(16#d0#)) OR
 					(reg_q545 AND symb_decoder(16#bf#)) OR
 					(reg_q545 AND symb_decoder(16#27#)) OR
 					(reg_q545 AND symb_decoder(16#e3#)) OR
 					(reg_q545 AND symb_decoder(16#48#)) OR
 					(reg_q545 AND symb_decoder(16#62#));
reg_q545_init <= '0' ;
	p_reg_q545: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q545 <= reg_q545_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q545 <= reg_q545_init;
        else
          reg_q545 <= reg_q545_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph5

reg_q2231_in <= (reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2229 AND symb_decoder(16#2f#));
reg_q2233_in <= (reg_q2231 AND symb_decoder(16#67#)) OR
 					(reg_q2231 AND symb_decoder(16#47#));
reg_q1961_in <= (reg_q1959 AND symb_decoder(16#7c#));
reg_q1672_in <= (reg_q1670 AND symb_decoder(16#3f#));
reg_q2429_in <= (reg_q2427 AND symb_decoder(16#3e#));
reg_q1602_in <= (reg_q1600 AND symb_decoder(16#65#)) OR
 					(reg_q1600 AND symb_decoder(16#45#));
reg_q1604_in <= (reg_q1602 AND symb_decoder(16#45#)) OR
 					(reg_q1602 AND symb_decoder(16#65#));
reg_q308_in <= (reg_q308 AND symb_decoder(16#0c#)) OR
 					(reg_q308 AND symb_decoder(16#09#)) OR
 					(reg_q308 AND symb_decoder(16#0a#)) OR
 					(reg_q308 AND symb_decoder(16#20#)) OR
 					(reg_q308 AND symb_decoder(16#0d#)) OR
 					(reg_q306 AND symb_decoder(16#0a#)) OR
 					(reg_q306 AND symb_decoder(16#09#)) OR
 					(reg_q306 AND symb_decoder(16#20#)) OR
 					(reg_q306 AND symb_decoder(16#0d#)) OR
 					(reg_q306 AND symb_decoder(16#0c#));
reg_q2651_in <= (reg_q2649 AND symb_decoder(16#7c#));
reg_q1443_in <= (reg_q1441 AND symb_decoder(16#6e#)) OR
 					(reg_q1441 AND symb_decoder(16#4e#));
reg_q644_in <= (reg_q642 AND symb_decoder(16#65#)) OR
 					(reg_q642 AND symb_decoder(16#45#));
reg_q646_in <= (reg_q644 AND symb_decoder(16#0d#)) OR
 					(reg_q644 AND symb_decoder(16#20#)) OR
 					(reg_q644 AND symb_decoder(16#09#)) OR
 					(reg_q644 AND symb_decoder(16#0c#)) OR
 					(reg_q644 AND symb_decoder(16#0a#)) OR
 					(reg_q646 AND symb_decoder(16#09#)) OR
 					(reg_q646 AND symb_decoder(16#0d#)) OR
 					(reg_q646 AND symb_decoder(16#20#)) OR
 					(reg_q646 AND symb_decoder(16#0a#)) OR
 					(reg_q646 AND symb_decoder(16#0c#));
reg_q179_in <= (reg_q179 AND symb_decoder(16#38#)) OR
 					(reg_q179 AND symb_decoder(16#34#)) OR
 					(reg_q179 AND symb_decoder(16#32#)) OR
 					(reg_q179 AND symb_decoder(16#39#)) OR
 					(reg_q179 AND symb_decoder(16#33#)) OR
 					(reg_q179 AND symb_decoder(16#30#)) OR
 					(reg_q179 AND symb_decoder(16#31#)) OR
 					(reg_q179 AND symb_decoder(16#35#)) OR
 					(reg_q179 AND symb_decoder(16#36#)) OR
 					(reg_q179 AND symb_decoder(16#37#)) OR
 					(reg_q177 AND symb_decoder(16#34#)) OR
 					(reg_q177 AND symb_decoder(16#37#)) OR
 					(reg_q177 AND symb_decoder(16#35#)) OR
 					(reg_q177 AND symb_decoder(16#32#)) OR
 					(reg_q177 AND symb_decoder(16#39#)) OR
 					(reg_q177 AND symb_decoder(16#33#)) OR
 					(reg_q177 AND symb_decoder(16#31#)) OR
 					(reg_q177 AND symb_decoder(16#36#)) OR
 					(reg_q177 AND symb_decoder(16#30#)) OR
 					(reg_q177 AND symb_decoder(16#38#));
reg_q634_in <= (reg_q632 AND symb_decoder(16#73#)) OR
 					(reg_q632 AND symb_decoder(16#53#));
reg_q636_in <= (reg_q634 AND symb_decoder(16#0c#)) OR
 					(reg_q634 AND symb_decoder(16#0a#)) OR
 					(reg_q634 AND symb_decoder(16#09#)) OR
 					(reg_q634 AND symb_decoder(16#20#)) OR
 					(reg_q634 AND symb_decoder(16#0d#)) OR
 					(reg_q636 AND symb_decoder(16#0a#)) OR
 					(reg_q636 AND symb_decoder(16#0d#)) OR
 					(reg_q636 AND symb_decoder(16#20#)) OR
 					(reg_q636 AND symb_decoder(16#0c#)) OR
 					(reg_q636 AND symb_decoder(16#09#));
reg_q2570_in <= (reg_q2570 AND symb_decoder(16#0a#)) OR
 					(reg_q2570 AND symb_decoder(16#0d#)) OR
 					(reg_q2570 AND symb_decoder(16#09#)) OR
 					(reg_q2570 AND symb_decoder(16#0c#)) OR
 					(reg_q2570 AND symb_decoder(16#20#)) OR
 					(reg_q2568 AND symb_decoder(16#20#)) OR
 					(reg_q2568 AND symb_decoder(16#09#)) OR
 					(reg_q2568 AND symb_decoder(16#0a#)) OR
 					(reg_q2568 AND symb_decoder(16#0c#)) OR
 					(reg_q2568 AND symb_decoder(16#0d#));
reg_q2572_in <= (reg_q2570 AND symb_decoder(16#4c#)) OR
 					(reg_q2570 AND symb_decoder(16#6c#));
reg_q2451_in <= (reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2449 AND symb_decoder(16#3c#));
reg_q2453_in <= (reg_q2451 AND symb_decoder(16#54#)) OR
 					(reg_q2451 AND symb_decoder(16#74#));
reg_q819_in <= (reg_q817 AND symb_decoder(16#3a#));
reg_q1377_in <= (reg_q1375 AND symb_decoder(16#6c#)) OR
 					(reg_q1375 AND symb_decoder(16#4c#));
reg_q1379_in <= (reg_q1377 AND symb_decoder(16#0c#)) OR
 					(reg_q1377 AND symb_decoder(16#09#)) OR
 					(reg_q1377 AND symb_decoder(16#0d#)) OR
 					(reg_q1377 AND symb_decoder(16#20#)) OR
 					(reg_q1377 AND symb_decoder(16#0a#)) OR
 					(reg_q1379 AND symb_decoder(16#0a#)) OR
 					(reg_q1379 AND symb_decoder(16#0c#)) OR
 					(reg_q1379 AND symb_decoder(16#20#)) OR
 					(reg_q1379 AND symb_decoder(16#0d#)) OR
 					(reg_q1379 AND symb_decoder(16#09#));
reg_q2534_in <= (reg_q2532 AND symb_decoder(16#5c#));
reg_q1890_in <= (reg_q1888 AND symb_decoder(16#33#));
reg_q1892_in <= (reg_q1890 AND symb_decoder(16#23#));
reg_q2082_in <= (reg_q2080 AND symb_decoder(16#45#)) OR
 					(reg_q2080 AND symb_decoder(16#65#));
reg_q2627_in <= (reg_q2625 AND symb_decoder(16#33#)) OR
 					(reg_q2625 AND symb_decoder(16#32#)) OR
 					(reg_q2625 AND symb_decoder(16#36#)) OR
 					(reg_q2625 AND symb_decoder(16#35#)) OR
 					(reg_q2625 AND symb_decoder(16#38#)) OR
 					(reg_q2625 AND symb_decoder(16#39#)) OR
 					(reg_q2625 AND symb_decoder(16#30#)) OR
 					(reg_q2625 AND symb_decoder(16#31#)) OR
 					(reg_q2625 AND symb_decoder(16#34#)) OR
 					(reg_q2625 AND symb_decoder(16#37#)) OR
 					(reg_q2627 AND symb_decoder(16#37#)) OR
 					(reg_q2627 AND symb_decoder(16#39#)) OR
 					(reg_q2627 AND symb_decoder(16#34#)) OR
 					(reg_q2627 AND symb_decoder(16#33#)) OR
 					(reg_q2627 AND symb_decoder(16#32#)) OR
 					(reg_q2627 AND symb_decoder(16#30#)) OR
 					(reg_q2627 AND symb_decoder(16#35#)) OR
 					(reg_q2627 AND symb_decoder(16#36#)) OR
 					(reg_q2627 AND symb_decoder(16#31#)) OR
 					(reg_q2627 AND symb_decoder(16#38#));
reg_q2150_in <= (reg_q2148 AND symb_decoder(16#54#)) OR
 					(reg_q2148 AND symb_decoder(16#74#));
reg_q316_in <= (reg_q314 AND symb_decoder(16#76#)) OR
 					(reg_q314 AND symb_decoder(16#56#));
reg_q318_in <= (reg_q316 AND symb_decoder(16#69#)) OR
 					(reg_q316 AND symb_decoder(16#49#));
reg_q620_in <= (reg_q618 AND symb_decoder(16#46#)) OR
 					(reg_q618 AND symb_decoder(16#66#));
reg_q622_in <= (reg_q620 AND symb_decoder(16#65#)) OR
 					(reg_q620 AND symb_decoder(16#45#));
reg_q1616_in <= (reg_q1614 AND symb_decoder(16#3f#));
reg_q2112_in <= (reg_q2110 AND symb_decoder(16#3f#));
reg_q2439_in <= (reg_q2437 AND symb_decoder(16#68#)) OR
 					(reg_q2437 AND symb_decoder(16#48#));
reg_q2441_in <= (reg_q2439 AND symb_decoder(16#61#)) OR
 					(reg_q2439 AND symb_decoder(16#41#));
reg_q2192_in <= (reg_q2190 AND symb_decoder(16#2d#));
reg_q2194_in <= (reg_q2192 AND symb_decoder(16#4e#)) OR
 					(reg_q2192 AND symb_decoder(16#6e#));
reg_q1524_in <= (reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q1522 AND symb_decoder(16#77#)) OR
 					(reg_q1522 AND symb_decoder(16#57#));
reg_q2092_in <= (reg_q2090 AND symb_decoder(16#5f#));
reg_q2094_in <= (reg_q2092 AND symb_decoder(16#54#)) OR
 					(reg_q2092 AND symb_decoder(16#74#));
reg_q439_in <= (reg_q437 AND symb_decoder(16#42#)) OR
 					(reg_q437 AND symb_decoder(16#62#));
reg_q441_in <= (reg_q439 AND symb_decoder(16#0c#)) OR
 					(reg_q439 AND symb_decoder(16#0d#)) OR
 					(reg_q439 AND symb_decoder(16#09#)) OR
 					(reg_q439 AND symb_decoder(16#0a#)) OR
 					(reg_q439 AND symb_decoder(16#20#)) OR
 					(reg_q441 AND symb_decoder(16#09#)) OR
 					(reg_q441 AND symb_decoder(16#0d#)) OR
 					(reg_q441 AND symb_decoder(16#0c#)) OR
 					(reg_q441 AND symb_decoder(16#0a#)) OR
 					(reg_q441 AND symb_decoder(16#20#));
reg_q488_in <= (reg_q486 AND symb_decoder(16#3a#));
reg_q490_in <= (reg_q488 AND symb_decoder(16#39#)) OR
 					(reg_q488 AND symb_decoder(16#30#)) OR
 					(reg_q488 AND symb_decoder(16#37#)) OR
 					(reg_q488 AND symb_decoder(16#33#)) OR
 					(reg_q488 AND symb_decoder(16#35#)) OR
 					(reg_q488 AND symb_decoder(16#38#)) OR
 					(reg_q488 AND symb_decoder(16#31#)) OR
 					(reg_q488 AND symb_decoder(16#32#)) OR
 					(reg_q488 AND symb_decoder(16#34#)) OR
 					(reg_q488 AND symb_decoder(16#36#)) OR
 					(reg_q490 AND symb_decoder(16#36#)) OR
 					(reg_q490 AND symb_decoder(16#30#)) OR
 					(reg_q490 AND symb_decoder(16#33#)) OR
 					(reg_q490 AND symb_decoder(16#32#)) OR
 					(reg_q490 AND symb_decoder(16#35#)) OR
 					(reg_q490 AND symb_decoder(16#31#)) OR
 					(reg_q490 AND symb_decoder(16#37#)) OR
 					(reg_q490 AND symb_decoder(16#39#)) OR
 					(reg_q490 AND symb_decoder(16#38#)) OR
 					(reg_q490 AND symb_decoder(16#34#));
reg_q173_in <= (reg_q173 AND symb_decoder(16#39#)) OR
 					(reg_q173 AND symb_decoder(16#36#)) OR
 					(reg_q173 AND symb_decoder(16#33#)) OR
 					(reg_q173 AND symb_decoder(16#32#)) OR
 					(reg_q173 AND symb_decoder(16#30#)) OR
 					(reg_q173 AND symb_decoder(16#35#)) OR
 					(reg_q173 AND symb_decoder(16#31#)) OR
 					(reg_q173 AND symb_decoder(16#37#)) OR
 					(reg_q173 AND symb_decoder(16#38#)) OR
 					(reg_q173 AND symb_decoder(16#34#)) OR
 					(reg_q171 AND symb_decoder(16#38#)) OR
 					(reg_q171 AND symb_decoder(16#35#)) OR
 					(reg_q171 AND symb_decoder(16#31#)) OR
 					(reg_q171 AND symb_decoder(16#39#)) OR
 					(reg_q171 AND symb_decoder(16#36#)) OR
 					(reg_q171 AND symb_decoder(16#32#)) OR
 					(reg_q171 AND symb_decoder(16#37#)) OR
 					(reg_q171 AND symb_decoder(16#30#)) OR
 					(reg_q171 AND symb_decoder(16#34#)) OR
 					(reg_q171 AND symb_decoder(16#33#));
reg_q2576_in <= (reg_q2574 AND symb_decoder(16#53#)) OR
 					(reg_q2574 AND symb_decoder(16#73#));
reg_q2578_in <= (reg_q2576 AND symb_decoder(16#74#)) OR
 					(reg_q2576 AND symb_decoder(16#54#));
reg_q1042_in <= (reg_q1040 AND symb_decoder(16#50#));
reg_q1044_in <= (reg_q1042 AND symb_decoder(16#0a#)) OR
 					(reg_q1042 AND symb_decoder(16#09#)) OR
 					(reg_q1042 AND symb_decoder(16#0c#)) OR
 					(reg_q1042 AND symb_decoder(16#0d#)) OR
 					(reg_q1042 AND symb_decoder(16#20#)) OR
 					(reg_q1044 AND symb_decoder(16#0c#)) OR
 					(reg_q1044 AND symb_decoder(16#20#)) OR
 					(reg_q1044 AND symb_decoder(16#09#)) OR
 					(reg_q1044 AND symb_decoder(16#0d#)) OR
 					(reg_q1044 AND symb_decoder(16#0a#));
reg_q2235_in <= (reg_q2233 AND symb_decoder(16#72#)) OR
 					(reg_q2233 AND symb_decoder(16#52#));
reg_q608_in <= (reg_q606 AND symb_decoder(16#52#)) OR
 					(reg_q606 AND symb_decoder(16#72#));
reg_q1658_in <= (reg_q1656 AND symb_decoder(16#65#)) OR
 					(reg_q1656 AND symb_decoder(16#45#));
reg_q1660_in <= (reg_q1658 AND symb_decoder(16#6d#)) OR
 					(reg_q1658 AND symb_decoder(16#4d#));
reg_q792_in <= (reg_q788 AND symb_decoder(16#32#)) OR
 					(reg_q800 AND symb_decoder(16#32#));
reg_q794_in <= (reg_q792 AND symb_decoder(16#2e#));
reg_q1606_in <= (reg_q1604 AND symb_decoder(16#64#)) OR
 					(reg_q1604 AND symb_decoder(16#44#));
reg_q312_in <= (reg_q310 AND symb_decoder(16#45#)) OR
 					(reg_q310 AND symb_decoder(16#65#));
reg_q314_in <= (reg_q312 AND symb_decoder(16#52#)) OR
 					(reg_q312 AND symb_decoder(16#72#));
reg_q2479_in <= (reg_q2479 AND symb_decoder(16#20#)) OR
 					(reg_q2479 AND symb_decoder(16#0c#)) OR
 					(reg_q2479 AND symb_decoder(16#0d#)) OR
 					(reg_q2479 AND symb_decoder(16#0a#)) OR
 					(reg_q2479 AND symb_decoder(16#09#)) OR
 					(reg_q2477 AND symb_decoder(16#0d#)) OR
 					(reg_q2477 AND symb_decoder(16#0c#)) OR
 					(reg_q2477 AND symb_decoder(16#0a#)) OR
 					(reg_q2477 AND symb_decoder(16#09#)) OR
 					(reg_q2477 AND symb_decoder(16#20#));
reg_q1526_in <= (reg_q1524 AND symb_decoder(16#49#)) OR
 					(reg_q1524 AND symb_decoder(16#69#));
reg_q1528_in <= (reg_q1526 AND symb_decoder(16#4e#)) OR
 					(reg_q1526 AND symb_decoder(16#6e#));
reg_q1844_in <= (reg_q1844 AND symb_decoder(16#0d#)) OR
 					(reg_q1844 AND symb_decoder(16#20#)) OR
 					(reg_q1844 AND symb_decoder(16#0a#)) OR
 					(reg_q1844 AND symb_decoder(16#0c#)) OR
 					(reg_q1844 AND symb_decoder(16#09#)) OR
 					(reg_q1842 AND symb_decoder(16#0a#)) OR
 					(reg_q1842 AND symb_decoder(16#09#)) OR
 					(reg_q1842 AND symb_decoder(16#0c#)) OR
 					(reg_q1842 AND symb_decoder(16#20#)) OR
 					(reg_q1842 AND symb_decoder(16#0d#));
reg_q890_in <= (reg_q888 AND symb_decoder(16#53#)) OR
 					(reg_q888 AND symb_decoder(16#73#));
reg_q892_in <= (reg_q890 AND symb_decoder(16#0a#)) OR
 					(reg_q890 AND symb_decoder(16#09#)) OR
 					(reg_q890 AND symb_decoder(16#0c#)) OR
 					(reg_q890 AND symb_decoder(16#20#)) OR
 					(reg_q890 AND symb_decoder(16#0d#)) OR
 					(reg_q892 AND symb_decoder(16#09#)) OR
 					(reg_q892 AND symb_decoder(16#0c#)) OR
 					(reg_q892 AND symb_decoder(16#0d#)) OR
 					(reg_q892 AND symb_decoder(16#0a#)) OR
 					(reg_q892 AND symb_decoder(16#20#));
reg_q183_in <= (reg_q183 AND symb_decoder(16#33#)) OR
 					(reg_q183 AND symb_decoder(16#32#)) OR
 					(reg_q183 AND symb_decoder(16#30#)) OR
 					(reg_q183 AND symb_decoder(16#37#)) OR
 					(reg_q183 AND symb_decoder(16#34#)) OR
 					(reg_q183 AND symb_decoder(16#38#)) OR
 					(reg_q183 AND symb_decoder(16#36#)) OR
 					(reg_q183 AND symb_decoder(16#31#)) OR
 					(reg_q183 AND symb_decoder(16#35#)) OR
 					(reg_q183 AND symb_decoder(16#39#)) OR
 					(reg_q181 AND symb_decoder(16#36#)) OR
 					(reg_q181 AND symb_decoder(16#30#)) OR
 					(reg_q181 AND symb_decoder(16#31#)) OR
 					(reg_q181 AND symb_decoder(16#38#)) OR
 					(reg_q181 AND symb_decoder(16#33#)) OR
 					(reg_q181 AND symb_decoder(16#37#)) OR
 					(reg_q181 AND symb_decoder(16#32#)) OR
 					(reg_q181 AND symb_decoder(16#39#)) OR
 					(reg_q181 AND symb_decoder(16#34#)) OR
 					(reg_q181 AND symb_decoder(16#35#));
reg_q2509_in <= (reg_q2507 AND symb_decoder(16#69#)) OR
 					(reg_q2507 AND symb_decoder(16#49#));
reg_q2511_in <= (reg_q2509 AND symb_decoder(16#74#)) OR
 					(reg_q2509 AND symb_decoder(16#54#));
reg_q1858_in <= (reg_q1856 AND symb_decoder(16#41#)) OR
 					(reg_q1856 AND symb_decoder(16#61#));
reg_q1860_in <= (reg_q1858 AND symb_decoder(16#09#)) OR
 					(reg_q1858 AND symb_decoder(16#0a#)) OR
 					(reg_q1858 AND symb_decoder(16#0c#)) OR
 					(reg_q1858 AND symb_decoder(16#20#)) OR
 					(reg_q1858 AND symb_decoder(16#0d#)) OR
 					(reg_q1860 AND symb_decoder(16#0c#)) OR
 					(reg_q1860 AND symb_decoder(16#0a#)) OR
 					(reg_q1860 AND symb_decoder(16#0d#)) OR
 					(reg_q1860 AND symb_decoder(16#20#)) OR
 					(reg_q1860 AND symb_decoder(16#09#));
reg_q290_in <= (reg_q288 AND symb_decoder(16#43#)) OR
 					(reg_q288 AND symb_decoder(16#63#));
reg_q292_in <= (reg_q290 AND symb_decoder(16#68#)) OR
 					(reg_q290 AND symb_decoder(16#48#));
reg_q2437_in <= (reg_q2435 AND symb_decoder(16#63#)) OR
 					(reg_q2435 AND symb_decoder(16#43#));
reg_q1473_in <= (reg_q1471 AND symb_decoder(16#6d#)) OR
 					(reg_q1471 AND symb_decoder(16#4d#));
reg_q1475_in <= (reg_q1473 AND symb_decoder(16#4f#)) OR
 					(reg_q1473 AND symb_decoder(16#6f#));
reg_q1260_in <= (reg_q1258 AND symb_decoder(16#75#)) OR
 					(reg_q1258 AND symb_decoder(16#55#));
reg_q1262_in <= (reg_q1260 AND symb_decoder(16#41#)) OR
 					(reg_q1260 AND symb_decoder(16#61#));
reg_q575_in <= (reg_q575 AND symb_decoder(16#38#)) OR
 					(reg_q575 AND symb_decoder(16#33#)) OR
 					(reg_q575 AND symb_decoder(16#31#)) OR
 					(reg_q575 AND symb_decoder(16#39#)) OR
 					(reg_q575 AND symb_decoder(16#32#)) OR
 					(reg_q575 AND symb_decoder(16#30#)) OR
 					(reg_q575 AND symb_decoder(16#36#)) OR
 					(reg_q575 AND symb_decoder(16#34#)) OR
 					(reg_q575 AND symb_decoder(16#37#)) OR
 					(reg_q575 AND symb_decoder(16#35#)) OR
 					(reg_q573 AND symb_decoder(16#32#)) OR
 					(reg_q573 AND symb_decoder(16#35#)) OR
 					(reg_q573 AND symb_decoder(16#38#)) OR
 					(reg_q573 AND symb_decoder(16#33#)) OR
 					(reg_q573 AND symb_decoder(16#37#)) OR
 					(reg_q573 AND symb_decoder(16#31#)) OR
 					(reg_q573 AND symb_decoder(16#30#)) OR
 					(reg_q573 AND symb_decoder(16#36#)) OR
 					(reg_q573 AND symb_decoder(16#39#)) OR
 					(reg_q573 AND symb_decoder(16#34#));
reg_q1427_in <= (reg_q1425 AND symb_decoder(16#41#)) OR
 					(reg_q1425 AND symb_decoder(16#61#));
reg_q1429_in <= (reg_q1427 AND symb_decoder(16#54#)) OR
 					(reg_q1427 AND symb_decoder(16#74#));
reg_q904_in <= (reg_q902 AND symb_decoder(16#72#)) OR
 					(reg_q902 AND symb_decoder(16#52#));
reg_q906_in <= (reg_q904 AND symb_decoder(16#09#)) OR
 					(reg_q904 AND symb_decoder(16#0c#)) OR
 					(reg_q904 AND symb_decoder(16#0d#)) OR
 					(reg_q904 AND symb_decoder(16#20#)) OR
 					(reg_q904 AND symb_decoder(16#0a#)) OR
 					(reg_q906 AND symb_decoder(16#09#)) OR
 					(reg_q906 AND symb_decoder(16#0c#)) OR
 					(reg_q906 AND symb_decoder(16#0a#)) OR
 					(reg_q906 AND symb_decoder(16#20#)) OR
 					(reg_q906 AND symb_decoder(16#0d#));
reg_q862_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q861 AND symb_decoder(16#53#)) OR
 					(reg_q861 AND symb_decoder(16#73#));
reg_q1832_in <= (reg_q1830 AND symb_decoder(16#70#)) OR
 					(reg_q1830 AND symb_decoder(16#50#));
reg_q1834_in <= (reg_q1832 AND symb_decoder(16#72#)) OR
 					(reg_q1832 AND symb_decoder(16#52#));
reg_q1610_in <= (reg_q1608 AND symb_decoder(16#50#)) OR
 					(reg_q1608 AND symb_decoder(16#70#));
reg_q1612_in <= (reg_q1610 AND symb_decoder(16#68#)) OR
 					(reg_q1610 AND symb_decoder(16#48#));
reg_q767_in <= (reg_q765 AND symb_decoder(16#54#)) OR
 					(reg_q765 AND symb_decoder(16#74#));
reg_q1546_in <= (reg_q1544 AND symb_decoder(16#45#)) OR
 					(reg_q1544 AND symb_decoder(16#65#));
reg_q1548_in <= (reg_q1546 AND symb_decoder(16#63#)) OR
 					(reg_q1546 AND symb_decoder(16#43#));
reg_q1854_in <= (reg_q1852 AND symb_decoder(16#53#)) OR
 					(reg_q1852 AND symb_decoder(16#73#));
reg_q1856_in <= (reg_q1854 AND symb_decoder(16#54#)) OR
 					(reg_q1854 AND symb_decoder(16#74#));
reg_q437_in <= (reg_q435 AND symb_decoder(16#65#)) OR
 					(reg_q435 AND symb_decoder(16#45#));
reg_q328_in <= (reg_q328 AND symb_decoder(16#0d#)) OR
 					(reg_q328 AND symb_decoder(16#0a#)) OR
 					(reg_q328 AND symb_decoder(16#09#)) OR
 					(reg_q328 AND symb_decoder(16#0c#)) OR
 					(reg_q328 AND symb_decoder(16#20#)) OR
 					(reg_q326 AND symb_decoder(16#0d#)) OR
 					(reg_q326 AND symb_decoder(16#09#)) OR
 					(reg_q326 AND symb_decoder(16#0a#)) OR
 					(reg_q326 AND symb_decoder(16#0c#)) OR
 					(reg_q326 AND symb_decoder(16#20#));
reg_q330_in <= (reg_q328 AND symb_decoder(16#70#)) OR
 					(reg_q328 AND symb_decoder(16#50#));
reg_q2190_in <= (reg_q2188 AND symb_decoder(16#41#)) OR
 					(reg_q2188 AND symb_decoder(16#61#));
reg_q1600_in <= (reg_q1598 AND symb_decoder(16#66#)) OR
 					(reg_q1598 AND symb_decoder(16#46#));
reg_q2560_in <= (reg_q2558 AND symb_decoder(16#64#)) OR
 					(reg_q2558 AND symb_decoder(16#44#));
reg_q2562_in <= (reg_q2560 AND symb_decoder(16#72#)) OR
 					(reg_q2560 AND symb_decoder(16#52#));
reg_q2168_in <= (reg_q2166 AND symb_decoder(16#4e#)) OR
 					(reg_q2166 AND symb_decoder(16#6e#));
reg_q2170_in <= (reg_q2168 AND symb_decoder(16#69#)) OR
 					(reg_q2168 AND symb_decoder(16#49#));
reg_q583_in <= (reg_q583 AND symb_decoder(16#33#)) OR
 					(reg_q583 AND symb_decoder(16#31#)) OR
 					(reg_q583 AND symb_decoder(16#38#)) OR
 					(reg_q583 AND symb_decoder(16#35#)) OR
 					(reg_q583 AND symb_decoder(16#36#)) OR
 					(reg_q583 AND symb_decoder(16#34#)) OR
 					(reg_q583 AND symb_decoder(16#39#)) OR
 					(reg_q583 AND symb_decoder(16#32#)) OR
 					(reg_q583 AND symb_decoder(16#30#)) OR
 					(reg_q583 AND symb_decoder(16#37#)) OR
 					(reg_q581 AND symb_decoder(16#38#)) OR
 					(reg_q581 AND symb_decoder(16#35#)) OR
 					(reg_q581 AND symb_decoder(16#39#)) OR
 					(reg_q581 AND symb_decoder(16#30#)) OR
 					(reg_q581 AND symb_decoder(16#33#)) OR
 					(reg_q581 AND symb_decoder(16#36#)) OR
 					(reg_q581 AND symb_decoder(16#37#)) OR
 					(reg_q581 AND symb_decoder(16#34#)) OR
 					(reg_q581 AND symb_decoder(16#31#)) OR
 					(reg_q581 AND symb_decoder(16#32#));
reg_q2568_in <= (reg_q2566 AND symb_decoder(16#45#)) OR
 					(reg_q2566 AND symb_decoder(16#65#));
reg_q1431_in <= (reg_q1429 AND symb_decoder(16#0c#)) OR
 					(reg_q1429 AND symb_decoder(16#0a#)) OR
 					(reg_q1429 AND symb_decoder(16#0d#)) OR
 					(reg_q1429 AND symb_decoder(16#09#)) OR
 					(reg_q1429 AND symb_decoder(16#20#)) OR
 					(reg_q1431 AND symb_decoder(16#09#)) OR
 					(reg_q1431 AND symb_decoder(16#0c#)) OR
 					(reg_q1431 AND symb_decoder(16#0a#)) OR
 					(reg_q1431 AND symb_decoder(16#20#)) OR
 					(reg_q1431 AND symb_decoder(16#0d#));
reg_q419_in <= (reg_q419 AND symb_decoder(16#20#)) OR
 					(reg_q419 AND symb_decoder(16#0a#)) OR
 					(reg_q419 AND symb_decoder(16#09#)) OR
 					(reg_q419 AND symb_decoder(16#0d#)) OR
 					(reg_q419 AND symb_decoder(16#0c#)) OR
 					(reg_q417 AND symb_decoder(16#20#)) OR
 					(reg_q417 AND symb_decoder(16#0c#)) OR
 					(reg_q417 AND symb_decoder(16#0d#)) OR
 					(reg_q417 AND symb_decoder(16#0a#)) OR
 					(reg_q417 AND symb_decoder(16#09#));
reg_q415_in <= (reg_q413 AND symb_decoder(16#45#)) OR
 					(reg_q413 AND symb_decoder(16#65#));
reg_q417_in <= (reg_q415 AND symb_decoder(16#54#)) OR
 					(reg_q415 AND symb_decoder(16#74#));
reg_q1266_in <= (reg_q1266 AND symb_decoder(16#0c#)) OR
 					(reg_q1266 AND symb_decoder(16#0d#)) OR
 					(reg_q1266 AND symb_decoder(16#0a#)) OR
 					(reg_q1266 AND symb_decoder(16#09#)) OR
 					(reg_q1266 AND symb_decoder(16#20#)) OR
 					(reg_q1264 AND symb_decoder(16#20#)) OR
 					(reg_q1264 AND symb_decoder(16#09#)) OR
 					(reg_q1264 AND symb_decoder(16#0a#)) OR
 					(reg_q1264 AND symb_decoder(16#0c#)) OR
 					(reg_q1264 AND symb_decoder(16#0d#));
reg_q2108_in <= (reg_q2106 AND symb_decoder(16#6f#)) OR
 					(reg_q2106 AND symb_decoder(16#4f#));
reg_q2110_in <= (reg_q2108 AND symb_decoder(16#75#)) OR
 					(reg_q2108 AND symb_decoder(16#55#));
reg_q1371_in <= (reg_q1369 AND symb_decoder(16#4f#)) OR
 					(reg_q1369 AND symb_decoder(16#6f#));
reg_q1373_in <= (reg_q1371 AND symb_decoder(16#6e#)) OR
 					(reg_q1371 AND symb_decoder(16#4e#));
reg_q786_in <= (reg_q784 AND symb_decoder(16#54#)) OR
 					(reg_q784 AND symb_decoder(16#74#));
reg_q2659_in <= (reg_q2657 AND symb_decoder(16#55#)) OR
 					(reg_q2657 AND symb_decoder(16#75#));
reg_q2661_in <= (reg_q2659 AND symb_decoder(16#52#)) OR
 					(reg_q2659 AND symb_decoder(16#72#));
reg_q1274_in <= (reg_q1272 AND symb_decoder(16#65#)) OR
 					(reg_q1272 AND symb_decoder(16#45#));
reg_q1276_in <= (reg_q1274 AND symb_decoder(16#0c#)) OR
 					(reg_q1274 AND symb_decoder(16#20#)) OR
 					(reg_q1274 AND symb_decoder(16#09#)) OR
 					(reg_q1274 AND symb_decoder(16#0d#)) OR
 					(reg_q1274 AND symb_decoder(16#0a#)) OR
 					(reg_q1276 AND symb_decoder(16#0d#)) OR
 					(reg_q1276 AND symb_decoder(16#0a#)) OR
 					(reg_q1276 AND symb_decoder(16#0c#)) OR
 					(reg_q1276 AND symb_decoder(16#09#)) OR
 					(reg_q1276 AND symb_decoder(16#20#));
reg_q2493_in <= (reg_q2493 AND symb_decoder(16#0c#)) OR
 					(reg_q2493 AND symb_decoder(16#0d#)) OR
 					(reg_q2493 AND symb_decoder(16#09#)) OR
 					(reg_q2493 AND symb_decoder(16#20#)) OR
 					(reg_q2493 AND symb_decoder(16#0a#)) OR
 					(reg_q2491 AND symb_decoder(16#09#)) OR
 					(reg_q2491 AND symb_decoder(16#0a#)) OR
 					(reg_q2491 AND symb_decoder(16#0c#)) OR
 					(reg_q2491 AND symb_decoder(16#0d#)) OR
 					(reg_q2491 AND symb_decoder(16#20#));
reg_q1375_in <= (reg_q1373 AND symb_decoder(16#61#)) OR
 					(reg_q1373 AND symb_decoder(16#41#));
reg_q1405_in <= (reg_q1403 AND symb_decoder(16#6f#)) OR
 					(reg_q1403 AND symb_decoder(16#4f#));
reg_q1407_in <= (reg_q1405 AND symb_decoder(16#54#)) OR
 					(reg_q1405 AND symb_decoder(16#74#));
reg_q916_in <= (reg_q914 AND symb_decoder(16#70#)) OR
 					(reg_q914 AND symb_decoder(16#50#));
reg_q918_in <= (reg_q916 AND symb_decoder(16#0d#)) OR
 					(reg_q916 AND symb_decoder(16#0c#)) OR
 					(reg_q916 AND symb_decoder(16#09#)) OR
 					(reg_q916 AND symb_decoder(16#20#)) OR
 					(reg_q916 AND symb_decoder(16#0a#)) OR
 					(reg_q918 AND symb_decoder(16#0d#)) OR
 					(reg_q918 AND symb_decoder(16#0a#)) OR
 					(reg_q918 AND symb_decoder(16#0c#)) OR
 					(reg_q918 AND symb_decoder(16#20#)) OR
 					(reg_q918 AND symb_decoder(16#09#));
reg_q2467_in <= (reg_q2465 AND symb_decoder(16#72#)) OR
 					(reg_q2465 AND symb_decoder(16#52#));
reg_q2469_in <= (reg_q2467 AND symb_decoder(16#6f#)) OR
 					(reg_q2467 AND symb_decoder(16#4f#));
reg_q1943_in <= (reg_q1941 AND symb_decoder(16#54#));
reg_q1232_in <= (reg_q1230 AND symb_decoder(16#45#)) OR
 					(reg_q1230 AND symb_decoder(16#65#));
reg_q1234_in <= (reg_q1232 AND symb_decoder(16#09#)) OR
 					(reg_q1232 AND symb_decoder(16#0c#)) OR
 					(reg_q1232 AND symb_decoder(16#0a#)) OR
 					(reg_q1232 AND symb_decoder(16#20#)) OR
 					(reg_q1232 AND symb_decoder(16#0d#)) OR
 					(reg_q1234 AND symb_decoder(16#0a#)) OR
 					(reg_q1234 AND symb_decoder(16#20#)) OR
 					(reg_q1234 AND symb_decoder(16#0d#)) OR
 					(reg_q1234 AND symb_decoder(16#0c#)) OR
 					(reg_q1234 AND symb_decoder(16#09#));
reg_q1477_in <= (reg_q1475 AND symb_decoder(16#4e#)) OR
 					(reg_q1475 AND symb_decoder(16#6e#));
reg_q1230_in <= (reg_q1228 AND symb_decoder(16#4d#)) OR
 					(reg_q1228 AND symb_decoder(16#6d#));
reg_q1250_in <= (reg_q1248 AND symb_decoder(16#4f#)) OR
 					(reg_q1248 AND symb_decoder(16#6f#));
reg_q1252_in <= (reg_q1250 AND symb_decoder(16#6d#)) OR
 					(reg_q1250 AND symb_decoder(16#4d#));
reg_q1423_in <= (reg_q1421 AND symb_decoder(16#52#)) OR
 					(reg_q1421 AND symb_decoder(16#72#));
reg_q1425_in <= (reg_q1423 AND symb_decoder(16#45#)) OR
 					(reg_q1423 AND symb_decoder(16#65#));
reg_q2212_in <= (reg_q2210 AND symb_decoder(16#7a#)) OR
 					(reg_q2210 AND symb_decoder(16#5a#));
reg_q2214_in <= (reg_q2212 AND symb_decoder(16#74#)) OR
 					(reg_q2212 AND symb_decoder(16#54#));
reg_q1288_in <= (reg_q1286 AND symb_decoder(16#66#)) OR
 					(reg_q1286 AND symb_decoder(16#46#));
reg_q1290_in <= (reg_q1288 AND symb_decoder(16#45#)) OR
 					(reg_q1288 AND symb_decoder(16#65#));
reg_q340_in <= (reg_q340 AND symb_decoder(16#20#)) OR
 					(reg_q340 AND symb_decoder(16#0d#)) OR
 					(reg_q340 AND symb_decoder(16#0a#)) OR
 					(reg_q340 AND symb_decoder(16#0c#)) OR
 					(reg_q340 AND symb_decoder(16#09#)) OR
 					(reg_q338 AND symb_decoder(16#20#)) OR
 					(reg_q338 AND symb_decoder(16#09#)) OR
 					(reg_q338 AND symb_decoder(16#0c#)) OR
 					(reg_q338 AND symb_decoder(16#0d#)) OR
 					(reg_q338 AND symb_decoder(16#0a#));
reg_q1622_in <= (reg_q1620 AND symb_decoder(16#78#)) OR
 					(reg_q1620 AND symb_decoder(16#58#));
reg_q624_in <= (reg_q622 AND symb_decoder(16#61#)) OR
 					(reg_q622 AND symb_decoder(16#41#));
reg_q423_in <= (reg_q421 AND symb_decoder(16#65#)) OR
 					(reg_q421 AND symb_decoder(16#45#));
reg_q425_in <= (reg_q423 AND symb_decoder(16#6d#)) OR
 					(reg_q423 AND symb_decoder(16#4d#));
reg_q1588_in <= (reg_q1586 AND symb_decoder(16#4c#)) OR
 					(reg_q1586 AND symb_decoder(16#6c#));
reg_q1590_in <= (reg_q1588 AND symb_decoder(16#75#)) OR
 					(reg_q1588 AND symb_decoder(16#55#));
reg_q332_in <= (reg_q330 AND symb_decoder(16#6f#)) OR
 					(reg_q330 AND symb_decoder(16#4f#));
reg_q2076_in <= (reg_q2074 AND symb_decoder(16#69#)) OR
 					(reg_q2074 AND symb_decoder(16#49#));
reg_q2078_in <= (reg_q2076 AND symb_decoder(16#70#)) OR
 					(reg_q2076 AND symb_decoder(16#50#));
reg_q1248_in <= (reg_q1248 AND symb_decoder(16#0d#)) OR
 					(reg_q1248 AND symb_decoder(16#20#)) OR
 					(reg_q1248 AND symb_decoder(16#0a#)) OR
 					(reg_q1248 AND symb_decoder(16#09#)) OR
 					(reg_q1248 AND symb_decoder(16#0c#)) OR
 					(reg_q1246 AND symb_decoder(16#0d#)) OR
 					(reg_q1246 AND symb_decoder(16#20#)) OR
 					(reg_q1246 AND symb_decoder(16#0a#)) OR
 					(reg_q1246 AND symb_decoder(16#09#)) OR
 					(reg_q1246 AND symb_decoder(16#0c#));
reg_q181_in <= (reg_q179 AND symb_decoder(16#2e#));
reg_q585_in <= (reg_q583 AND symb_decoder(16#23#));
reg_q334_in <= (reg_q332 AND symb_decoder(16#52#)) OR
 					(reg_q332 AND symb_decoder(16#72#));
reg_q2124_in <= (reg_q2122 AND symb_decoder(16#5f#));
reg_q2126_in <= (reg_q2124 AND symb_decoder(16#4e#)) OR
 					(reg_q2124 AND symb_decoder(16#6e#));
reg_q2558_in <= (reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2556 AND symb_decoder(16#5b#));
reg_q1449_in <= (reg_q1447 AND symb_decoder(16#69#)) OR
 					(reg_q1447 AND symb_decoder(16#49#));
reg_q1451_in <= (reg_q1449 AND symb_decoder(16#43#)) OR
 					(reg_q1449 AND symb_decoder(16#63#));
reg_q835_in <= (reg_q833 AND symb_decoder(16#49#)) OR
 					(reg_q833 AND symb_decoder(16#69#));
reg_q837_in <= (reg_q835 AND symb_decoder(16#6e#)) OR
 					(reg_q835 AND symb_decoder(16#4e#));
reg_q626_in <= (reg_q624 AND symb_decoder(16#72#)) OR
 					(reg_q624 AND symb_decoder(16#52#));
reg_q628_in <= (reg_q626 AND symb_decoder(16#6c#)) OR
 					(reg_q626 AND symb_decoder(16#4c#));
reg_q1258_in <= (reg_q1256 AND symb_decoder(16#71#)) OR
 					(reg_q1256 AND symb_decoder(16#51#));
reg_q1558_in <= (reg_q1558 AND symb_decoder(16#0a#)) OR
 					(reg_q1558 AND symb_decoder(16#0c#)) OR
 					(reg_q1558 AND symb_decoder(16#09#)) OR
 					(reg_q1558 AND symb_decoder(16#0d#)) OR
 					(reg_q1558 AND symb_decoder(16#20#)) OR
 					(reg_q1556 AND symb_decoder(16#09#)) OR
 					(reg_q1556 AND symb_decoder(16#0c#)) OR
 					(reg_q1556 AND symb_decoder(16#20#)) OR
 					(reg_q1556 AND symb_decoder(16#0d#)) OR
 					(reg_q1556 AND symb_decoder(16#0a#));
reg_q1668_in <= (reg_q1666 AND symb_decoder(16#68#)) OR
 					(reg_q1666 AND symb_decoder(16#48#));
reg_q1670_in <= (reg_q1668 AND symb_decoder(16#70#)) OR
 					(reg_q1668 AND symb_decoder(16#50#));
reg_q1570_in <= (reg_q1568 AND symb_decoder(16#45#)) OR
 					(reg_q1568 AND symb_decoder(16#65#));
reg_q1572_in <= (reg_q1570 AND symb_decoder(16#64#)) OR
 					(reg_q1570 AND symb_decoder(16#44#));
reg_q1580_in <= (reg_q1578 AND symb_decoder(16#2d#));
reg_q1582_in <= (reg_q1580 AND symb_decoder(16#69#)) OR
 					(reg_q1580 AND symb_decoder(16#49#));
reg_q841_in <= (reg_q841 AND symb_decoder(16#09#)) OR
 					(reg_q841 AND symb_decoder(16#0d#)) OR
 					(reg_q841 AND symb_decoder(16#0c#)) OR
 					(reg_q841 AND symb_decoder(16#0a#)) OR
 					(reg_q841 AND symb_decoder(16#20#)) OR
 					(reg_q839 AND symb_decoder(16#20#)) OR
 					(reg_q839 AND symb_decoder(16#0a#)) OR
 					(reg_q839 AND symb_decoder(16#09#)) OR
 					(reg_q839 AND symb_decoder(16#0d#)) OR
 					(reg_q839 AND symb_decoder(16#0c#));
reg_q652_in <= (reg_q650 AND symb_decoder(16#52#)) OR
 					(reg_q650 AND symb_decoder(16#72#));
reg_q654_in <= (reg_q652 AND symb_decoder(16#76#)) OR
 					(reg_q652 AND symb_decoder(16#56#));
reg_q1409_in <= (reg_q1407 AND symb_decoder(16#09#)) OR
 					(reg_q1407 AND symb_decoder(16#0d#)) OR
 					(reg_q1407 AND symb_decoder(16#20#)) OR
 					(reg_q1407 AND symb_decoder(16#0c#)) OR
 					(reg_q1407 AND symb_decoder(16#0a#)) OR
 					(reg_q1409 AND symb_decoder(16#20#)) OR
 					(reg_q1409 AND symb_decoder(16#0c#)) OR
 					(reg_q1409 AND symb_decoder(16#09#)) OR
 					(reg_q1409 AND symb_decoder(16#0d#)) OR
 					(reg_q1409 AND symb_decoder(16#0a#));
reg_q839_in <= (reg_q837 AND symb_decoder(16#45#)) OR
 					(reg_q837 AND symb_decoder(16#65#));
reg_q1421_in <= (reg_q1419 AND symb_decoder(16#67#)) OR
 					(reg_q1419 AND symb_decoder(16#47#));
reg_q912_in <= (reg_q912 AND symb_decoder(16#0a#)) OR
 					(reg_q912 AND symb_decoder(16#20#)) OR
 					(reg_q912 AND symb_decoder(16#0c#)) OR
 					(reg_q912 AND symb_decoder(16#0d#)) OR
 					(reg_q912 AND symb_decoder(16#09#)) OR
 					(reg_q910 AND symb_decoder(16#0a#)) OR
 					(reg_q910 AND symb_decoder(16#0c#)) OR
 					(reg_q910 AND symb_decoder(16#0d#)) OR
 					(reg_q910 AND symb_decoder(16#09#)) OR
 					(reg_q910 AND symb_decoder(16#20#));
reg_q1272_in <= (reg_q1270 AND symb_decoder(16#6c#)) OR
 					(reg_q1270 AND symb_decoder(16#4c#));
reg_q1614_in <= (reg_q1612 AND symb_decoder(16#50#)) OR
 					(reg_q1612 AND symb_decoder(16#70#));
reg_q2530_in <= (reg_q2526 AND symb_decoder(16#3b#)) OR
 					(reg_q2554 AND symb_decoder(16#3b#));
reg_q2532_in <= (reg_q2530 AND symb_decoder(16#5c#));
reg_q928_in <= (reg_q926 AND symb_decoder(16#52#)) OR
 					(reg_q926 AND symb_decoder(16#72#));
reg_q930_in <= (reg_q928 AND symb_decoder(16#75#)) OR
 					(reg_q928 AND symb_decoder(16#55#));
reg_q2198_in <= (reg_q2196 AND symb_decoder(16#74#)) OR
 					(reg_q2196 AND symb_decoder(16#54#));
reg_q2200_in <= (reg_q2198 AND symb_decoder(16#69#)) OR
 					(reg_q2198 AND symb_decoder(16#49#));
reg_q503_in <= (reg_q501 AND symb_decoder(16#4e#)) OR
 					(reg_q501 AND symb_decoder(16#6e#));
reg_q2146_in <= (reg_q2144 AND symb_decoder(16#45#)) OR
 					(reg_q2144 AND symb_decoder(16#65#));
reg_q2148_in <= (reg_q2146 AND symb_decoder(16#73#)) OR
 					(reg_q2146 AND symb_decoder(16#53#));
reg_q926_in <= (reg_q926 AND symb_decoder(16#0d#)) OR
 					(reg_q926 AND symb_decoder(16#0c#)) OR
 					(reg_q926 AND symb_decoder(16#20#)) OR
 					(reg_q926 AND symb_decoder(16#0a#)) OR
 					(reg_q926 AND symb_decoder(16#09#)) OR
 					(reg_q924 AND symb_decoder(16#0d#)) OR
 					(reg_q924 AND symb_decoder(16#0c#)) OR
 					(reg_q924 AND symb_decoder(16#20#)) OR
 					(reg_q924 AND symb_decoder(16#0a#)) OR
 					(reg_q924 AND symb_decoder(16#09#));
reg_q1325_in <= (reg_q1323 AND symb_decoder(16#74#)) OR
 					(reg_q1323 AND symb_decoder(16#54#));
reg_q549_in <= (reg_q547 AND symb_decoder(16#49#)) OR
 					(reg_q547 AND symb_decoder(16#69#));
reg_q403_in <= (reg_q401 AND symb_decoder(16#68#)) OR
 					(reg_q401 AND symb_decoder(16#48#));
reg_q2188_in <= (reg_q2186 AND symb_decoder(16#49#)) OR
 					(reg_q2186 AND symb_decoder(16#69#));
reg_q898_in <= (reg_q896 AND symb_decoder(16#52#)) OR
 					(reg_q896 AND symb_decoder(16#72#));
reg_q900_in <= (reg_q898 AND symb_decoder(16#56#)) OR
 					(reg_q898 AND symb_decoder(16#76#));
reg_q630_in <= (reg_q628 AND symb_decoder(16#65#)) OR
 					(reg_q628 AND symb_decoder(16#45#));
reg_q632_in <= (reg_q630 AND symb_decoder(16#73#)) OR
 					(reg_q630 AND symb_decoder(16#53#));
reg_q1455_in <= (reg_q1453 AND symb_decoder(16#69#)) OR
 					(reg_q1453 AND symb_decoder(16#49#));
reg_q1254_in <= (reg_q1252 AND symb_decoder(16#4e#)) OR
 					(reg_q1252 AND symb_decoder(16#6e#));
reg_q1256_in <= (reg_q1254 AND symb_decoder(16#49#)) OR
 					(reg_q1254 AND symb_decoder(16#69#));
reg_q1138_in <= (reg_q1136 AND symb_decoder(16#54#)) OR
 					(reg_q1136 AND symb_decoder(16#74#));
reg_q1278_in <= (reg_q1276 AND symb_decoder(16#54#)) OR
 					(reg_q1276 AND symb_decoder(16#74#));
reg_q1280_in <= (reg_q1278 AND symb_decoder(16#52#)) OR
 					(reg_q1278 AND symb_decoder(16#72#));
reg_q656_in <= (reg_q654 AND symb_decoder(16#45#)) OR
 					(reg_q654 AND symb_decoder(16#65#));
reg_q2540_in <= (reg_q2538 AND symb_decoder(16#53#)) OR
 					(reg_q2538 AND symb_decoder(16#73#));
reg_q2542_in <= (reg_q2540 AND symb_decoder(16#76#)) OR
 					(reg_q2540 AND symb_decoder(16#56#));
reg_q910_in <= (reg_q908 AND symb_decoder(16#53#)) OR
 					(reg_q908 AND symb_decoder(16#73#));
reg_q2176_in <= (reg_q2174 AND symb_decoder(16#6e#)) OR
 					(reg_q2174 AND symb_decoder(16#4e#));
reg_q2178_in <= (reg_q2176 AND symb_decoder(16#61#)) OR
 					(reg_q2176 AND symb_decoder(16#41#));
reg_q2070_in <= (reg_q2068 AND symb_decoder(16#64#)) OR
 					(reg_q2068 AND symb_decoder(16#44#));
reg_q2072_in <= (reg_q2070 AND symb_decoder(16#73#)) OR
 					(reg_q2070 AND symb_decoder(16#53#));
reg_q1242_in <= (reg_q1240 AND symb_decoder(16#74#)) OR
 					(reg_q1240 AND symb_decoder(16#54#));
reg_q1244_in <= (reg_q1242 AND symb_decoder(16#68#)) OR
 					(reg_q1242 AND symb_decoder(16#48#));
reg_q2156_in <= (reg_q2154 AND symb_decoder(16#52#)) OR
 					(reg_q2154 AND symb_decoder(16#72#));
reg_q2158_in <= (reg_q2156 AND symb_decoder(16#49#)) OR
 					(reg_q2156 AND symb_decoder(16#69#));
reg_q2465_in <= (reg_q2463 AND symb_decoder(16#74#)) OR
 					(reg_q2463 AND symb_decoder(16#54#));
reg_q924_in <= (reg_q922 AND symb_decoder(16#64#)) OR
 					(reg_q922 AND symb_decoder(16#44#));
reg_q2088_in <= (reg_q2086 AND symb_decoder(16#49#)) OR
 					(reg_q2086 AND symb_decoder(16#69#));
reg_q2090_in <= (reg_q2088 AND symb_decoder(16#6c#)) OR
 					(reg_q2088 AND symb_decoder(16#4c#));
reg_q2066_in <= (reg_q2064 AND symb_decoder(16#45#)) OR
 					(reg_q2064 AND symb_decoder(16#65#));
reg_q870_in <= (reg_q868 AND symb_decoder(16#45#)) OR
 					(reg_q868 AND symb_decoder(16#65#));
reg_q2184_in <= (reg_q2182 AND symb_decoder(16#3d#));
reg_q2186_in <= (reg_q2184 AND symb_decoder(16#63#)) OR
 					(reg_q2184 AND symb_decoder(16#43#));
reg_q864_in <= (reg_q862 AND symb_decoder(16#75#)) OR
 					(reg_q862 AND symb_decoder(16#55#));
reg_q866_in <= (reg_q864 AND symb_decoder(16#62#)) OR
 					(reg_q864 AND symb_decoder(16#42#));
reg_q2497_in <= (reg_q2495 AND symb_decoder(16#6f#)) OR
 					(reg_q2495 AND symb_decoder(16#4f#));
reg_q433_in <= (reg_q433 AND symb_decoder(16#09#)) OR
 					(reg_q433 AND symb_decoder(16#0d#)) OR
 					(reg_q433 AND symb_decoder(16#0c#)) OR
 					(reg_q433 AND symb_decoder(16#0a#)) OR
 					(reg_q433 AND symb_decoder(16#20#)) OR
 					(reg_q431 AND symb_decoder(16#0a#)) OR
 					(reg_q431 AND symb_decoder(16#0c#)) OR
 					(reg_q431 AND symb_decoder(16#0d#)) OR
 					(reg_q431 AND symb_decoder(16#09#)) OR
 					(reg_q431 AND symb_decoder(16#20#));
reg_q1822_in <= (reg_q1820 AND symb_decoder(16#23#));
reg_q1662_in <= (reg_q1660 AND symb_decoder(16#45#)) OR
 					(reg_q1660 AND symb_decoder(16#65#));
reg_q2120_in <= (reg_q2118 AND symb_decoder(16#63#)) OR
 					(reg_q2118 AND symb_decoder(16#43#));
reg_q1236_in <= (reg_q1234 AND symb_decoder(16#54#)) OR
 					(reg_q1234 AND symb_decoder(16#74#));
reg_q1036_in <= (reg_q1034 AND symb_decoder(16#0d#)) OR
 					(reg_q1034 AND symb_decoder(16#20#)) OR
 					(reg_q1034 AND symb_decoder(16#0a#)) OR
 					(reg_q1034 AND symb_decoder(16#09#)) OR
 					(reg_q1034 AND symb_decoder(16#0c#)) OR
 					(reg_q1036 AND symb_decoder(16#09#)) OR
 					(reg_q1036 AND symb_decoder(16#20#)) OR
 					(reg_q1036 AND symb_decoder(16#0c#)) OR
 					(reg_q1036 AND symb_decoder(16#0a#)) OR
 					(reg_q1036 AND symb_decoder(16#0d#));
reg_q1538_in <= (reg_q1538 AND symb_decoder(16#20#)) OR
 					(reg_q1538 AND symb_decoder(16#0d#)) OR
 					(reg_q1538 AND symb_decoder(16#0c#)) OR
 					(reg_q1538 AND symb_decoder(16#0a#)) OR
 					(reg_q1538 AND symb_decoder(16#09#)) OR
 					(reg_q1536 AND symb_decoder(16#0d#)) OR
 					(reg_q1536 AND symb_decoder(16#0a#)) OR
 					(reg_q1536 AND symb_decoder(16#09#)) OR
 					(reg_q1536 AND symb_decoder(16#0c#)) OR
 					(reg_q1536 AND symb_decoder(16#20#));
reg_q1540_in <= (reg_q1538 AND symb_decoder(16#64#)) OR
 					(reg_q1538 AND symb_decoder(16#44#));
reg_q1550_in <= (reg_q1548 AND symb_decoder(16#74#)) OR
 					(reg_q1548 AND symb_decoder(16#54#));
reg_q1552_in <= (reg_q1550 AND symb_decoder(16#4f#)) OR
 					(reg_q1550 AND symb_decoder(16#6f#));
reg_q742_in <= (reg_q740 AND symb_decoder(16#65#)) OR
 					(reg_q740 AND symb_decoder(16#45#));
reg_q2671_in <= (reg_q2669 AND symb_decoder(16#2e#));
reg_q1284_in <= (reg_q1282 AND symb_decoder(16#6e#)) OR
 					(reg_q1282 AND symb_decoder(16#4e#));
reg_q1286_in <= (reg_q1284 AND symb_decoder(16#73#)) OR
 					(reg_q1284 AND symb_decoder(16#53#));
reg_q1850_in <= (reg_q1850 AND symb_decoder(16#20#)) OR
 					(reg_q1850 AND symb_decoder(16#0c#)) OR
 					(reg_q1850 AND symb_decoder(16#09#)) OR
 					(reg_q1850 AND symb_decoder(16#0d#)) OR
 					(reg_q1850 AND symb_decoder(16#0a#)) OR
 					(reg_q1848 AND symb_decoder(16#0c#)) OR
 					(reg_q1848 AND symb_decoder(16#20#)) OR
 					(reg_q1848 AND symb_decoder(16#0d#)) OR
 					(reg_q1848 AND symb_decoder(16#09#)) OR
 					(reg_q1848 AND symb_decoder(16#0a#));
reg_q1852_in <= (reg_q1850 AND symb_decoder(16#45#)) OR
 					(reg_q1850 AND symb_decoder(16#65#));
reg_q1731_in <= (reg_q1729 AND symb_decoder(16#45#)) OR
 					(reg_q1729 AND symb_decoder(16#65#));
reg_q1733_in <= (reg_q1731 AND symb_decoder(16#72#)) OR
 					(reg_q1731 AND symb_decoder(16#52#));
reg_q612_in <= (reg_q610 AND symb_decoder(16#49#)) OR
 					(reg_q610 AND symb_decoder(16#69#));
reg_q614_in <= (reg_q612 AND symb_decoder(16#4e#)) OR
 					(reg_q612 AND symb_decoder(16#6e#));
reg_q825_in <= (reg_q823 AND symb_decoder(16#6d#)) OR
 					(reg_q823 AND symb_decoder(16#4d#));
reg_q2206_in <= (reg_q2204 AND symb_decoder(16#2d#));
reg_q2208_in <= (reg_q2206 AND symb_decoder(16#74#)) OR
 					(reg_q2206 AND symb_decoder(16#54#));
reg_q1648_in <= (reg_q1646 AND symb_decoder(16#65#)) OR
 					(reg_q1646 AND symb_decoder(16#45#));
reg_q1650_in <= (reg_q1648 AND symb_decoder(16#53#)) OR
 					(reg_q1648 AND symb_decoder(16#73#));
reg_q1401_in <= (reg_q1401 AND symb_decoder(16#0a#)) OR
 					(reg_q1401 AND symb_decoder(16#20#)) OR
 					(reg_q1401 AND symb_decoder(16#09#)) OR
 					(reg_q1401 AND symb_decoder(16#0d#)) OR
 					(reg_q1401 AND symb_decoder(16#0c#)) OR
 					(reg_q1399 AND symb_decoder(16#0d#)) OR
 					(reg_q1399 AND symb_decoder(16#20#)) OR
 					(reg_q1399 AND symb_decoder(16#09#)) OR
 					(reg_q1399 AND symb_decoder(16#0c#)) OR
 					(reg_q1399 AND symb_decoder(16#0a#));
reg_q1888_in <= (reg_q1886 AND symb_decoder(16#23#));
reg_q2471_in <= (reg_q2469 AND symb_decoder(16#79#)) OR
 					(reg_q2469 AND symb_decoder(16#59#));
reg_q2473_in <= (reg_q2471 AND symb_decoder(16#61#)) OR
 					(reg_q2471 AND symb_decoder(16#41#));
reg_q326_in <= (reg_q324 AND symb_decoder(16#2e#));
reg_q1471_in <= (reg_q1469 AND symb_decoder(16#45#)) OR
 					(reg_q1469 AND symb_decoder(16#65#));
reg_q1246_in <= (reg_q1244 AND symb_decoder(16#45#)) OR
 					(reg_q1244 AND symb_decoder(16#65#));
reg_q2742_in <= (reg_q2740 AND symb_decoder(16#61#)) OR
 					(reg_q2740 AND symb_decoder(16#41#));
reg_q2421_in <= (reg_q2419 AND symb_decoder(16#63#)) OR
 					(reg_q2419 AND symb_decoder(16#43#));
reg_q2423_in <= (reg_q2421 AND symb_decoder(16#68#)) OR
 					(reg_q2421 AND symb_decoder(16#48#));
reg_q579_in <= (reg_q579 AND symb_decoder(16#31#)) OR
 					(reg_q579 AND symb_decoder(16#33#)) OR
 					(reg_q579 AND symb_decoder(16#30#)) OR
 					(reg_q579 AND symb_decoder(16#39#)) OR
 					(reg_q579 AND symb_decoder(16#36#)) OR
 					(reg_q579 AND symb_decoder(16#37#)) OR
 					(reg_q579 AND symb_decoder(16#38#)) OR
 					(reg_q579 AND symb_decoder(16#32#)) OR
 					(reg_q579 AND symb_decoder(16#34#)) OR
 					(reg_q579 AND symb_decoder(16#35#)) OR
 					(reg_q577 AND symb_decoder(16#34#)) OR
 					(reg_q577 AND symb_decoder(16#37#)) OR
 					(reg_q577 AND symb_decoder(16#33#)) OR
 					(reg_q577 AND symb_decoder(16#30#)) OR
 					(reg_q577 AND symb_decoder(16#38#)) OR
 					(reg_q577 AND symb_decoder(16#36#)) OR
 					(reg_q577 AND symb_decoder(16#35#)) OR
 					(reg_q577 AND symb_decoder(16#31#)) OR
 					(reg_q577 AND symb_decoder(16#32#)) OR
 					(reg_q577 AND symb_decoder(16#39#));
reg_q932_in <= (reg_q930 AND symb_decoder(16#4e#)) OR
 					(reg_q930 AND symb_decoder(16#6e#));
reg_q934_in <= (reg_q932 AND symb_decoder(16#4e#)) OR
 					(reg_q932 AND symb_decoder(16#6e#));
reg_q1907_in <= (reg_q1905 AND symb_decoder(16#52#));
reg_q1367_in <= (reg_q1365 AND symb_decoder(16#54#)) OR
 					(reg_q1365 AND symb_decoder(16#74#));
reg_q2665_in <= (reg_q2665 AND symb_decoder(16#20#)) OR
 					(reg_q2665 AND symb_decoder(16#0a#)) OR
 					(reg_q2665 AND symb_decoder(16#0c#)) OR
 					(reg_q2665 AND symb_decoder(16#09#)) OR
 					(reg_q2665 AND symb_decoder(16#0d#)) OR
 					(reg_q2663 AND symb_decoder(16#0c#)) OR
 					(reg_q2663 AND symb_decoder(16#0a#)) OR
 					(reg_q2663 AND symb_decoder(16#09#)) OR
 					(reg_q2663 AND symb_decoder(16#20#)) OR
 					(reg_q2663 AND symb_decoder(16#0d#));
reg_q2667_in <= (reg_q2665 AND symb_decoder(16#56#)) OR
 					(reg_q2665 AND symb_decoder(16#76#));
reg_q1638_in <= (reg_q1636 AND symb_decoder(16#6e#)) OR
 					(reg_q1636 AND symb_decoder(16#4e#));
reg_q1967_in <= (reg_q1965 AND symb_decoder(16#2d#));
reg_q1866_in <= (reg_q1864 AND symb_decoder(16#6e#)) OR
 					(reg_q1864 AND symb_decoder(16#4e#));
reg_q1868_in <= (reg_q1866 AND symb_decoder(16#45#)) OR
 					(reg_q1866 AND symb_decoder(16#65#));
reg_q1304_in <= (reg_q1302 AND symb_decoder(16#65#)) OR
 					(reg_q1302 AND symb_decoder(16#45#));
reg_q1306_in <= (reg_q1304 AND symb_decoder(16#52#)) OR
 					(reg_q1304 AND symb_decoder(16#72#));
reg_q2513_in <= (reg_q2511 AND symb_decoder(16#4c#)) OR
 					(reg_q2511 AND symb_decoder(16#6c#));
reg_q1870_in <= (reg_q1868 AND symb_decoder(16#63#)) OR
 					(reg_q1868 AND symb_decoder(16#43#));
reg_q1872_in <= (reg_q1870 AND symb_decoder(16#74#)) OR
 					(reg_q1870 AND symb_decoder(16#54#));
reg_q1969_in <= (reg_q1967 AND symb_decoder(16#2d#));
reg_q1971_in <= (reg_q1969 AND symb_decoder(16#2d#));
reg_q577_in <= (reg_q575 AND symb_decoder(16#2e#));
reg_q413_in <= (reg_q411 AND symb_decoder(16#6e#)) OR
 					(reg_q411 AND symb_decoder(16#4e#));
reg_q405_in <= (reg_q403 AND symb_decoder(16#61#)) OR
 					(reg_q403 AND symb_decoder(16#41#));
reg_q407_in <= (reg_q405 AND symb_decoder(16#44#)) OR
 					(reg_q405 AND symb_decoder(16#64#));
reg_q2564_in <= (reg_q2562 AND symb_decoder(16#49#)) OR
 					(reg_q2562 AND symb_decoder(16#69#));
reg_q2740_in <= (reg_q2738 AND symb_decoder(16#54#)) OR
 					(reg_q2738 AND symb_decoder(16#74#));
reg_q2477_in <= (reg_q2475 AND symb_decoder(16#2d#));
reg_q1632_in <= (reg_q1630 AND symb_decoder(16#70#)) OR
 					(reg_q1630 AND symb_decoder(16#50#));
reg_q306_in <= (reg_q304 AND symb_decoder(16#52#)) OR
 					(reg_q304 AND symb_decoder(16#72#));
reg_q2174_in <= (reg_q2172 AND symb_decoder(16#6b#)) OR
 					(reg_q2172 AND symb_decoder(16#4b#));
reg_q1282_in <= (reg_q1280 AND symb_decoder(16#61#)) OR
 					(reg_q1280 AND symb_decoder(16#41#));
reg_q2084_in <= (reg_q2082 AND symb_decoder(16#6d#)) OR
 					(reg_q2082 AND symb_decoder(16#4d#));
reg_q1955_in <= (reg_q1953 AND symb_decoder(16#2d#));
reg_q1957_in <= (reg_q1955 AND symb_decoder(16#2d#));
reg_q1238_in <= (reg_q1236 AND symb_decoder(16#4f#)) OR
 					(reg_q1236 AND symb_decoder(16#6f#));
reg_q922_in <= (reg_q920 AND symb_decoder(16#4e#)) OR
 					(reg_q920 AND symb_decoder(16#6e#));
reg_q2457_in <= (reg_q2455 AND symb_decoder(16#54#)) OR
 					(reg_q2455 AND symb_decoder(16#74#));
reg_q2459_in <= (reg_q2457 AND symb_decoder(16#6c#)) OR
 					(reg_q2457 AND symb_decoder(16#4c#));
reg_q463_in <= (reg_q461 AND symb_decoder(16#41#)) OR
 					(reg_q461 AND symb_decoder(16#61#));
reg_q465_in <= (reg_q463 AND symb_decoder(16#72#)) OR
 					(reg_q463 AND symb_decoder(16#52#));
reg_q320_in <= (reg_q318 AND symb_decoder(16#44#)) OR
 					(reg_q318 AND symb_decoder(16#64#));
reg_q322_in <= (reg_q320 AND symb_decoder(16#6f#)) OR
 					(reg_q320 AND symb_decoder(16#4f#));
reg_q2475_in <= (reg_q2473 AND symb_decoder(16#20#)) OR
 					(reg_q2473 AND symb_decoder(16#0c#)) OR
 					(reg_q2473 AND symb_decoder(16#0d#)) OR
 					(reg_q2473 AND symb_decoder(16#09#)) OR
 					(reg_q2473 AND symb_decoder(16#0a#)) OR
 					(reg_q2475 AND symb_decoder(16#0c#)) OR
 					(reg_q2475 AND symb_decoder(16#0a#)) OR
 					(reg_q2475 AND symb_decoder(16#09#)) OR
 					(reg_q2475 AND symb_decoder(16#20#)) OR
 					(reg_q2475 AND symb_decoder(16#0d#));
reg_q1901_in <= (reg_q2757 AND symb_decoder(16#2a#));
reg_q457_in <= (reg_q455 AND symb_decoder(16#50#)) OR
 					(reg_q455 AND symb_decoder(16#70#));
reg_q459_in <= (reg_q457 AND symb_decoder(16#59#)) OR
 					(reg_q457 AND symb_decoder(16#79#));
reg_q1560_in <= (reg_q1558 AND symb_decoder(16#46#)) OR
 					(reg_q1558 AND symb_decoder(16#66#));
reg_q1562_in <= (reg_q1560 AND symb_decoder(16#4c#)) OR
 					(reg_q1560 AND symb_decoder(16#6c#));
reg_q336_in <= (reg_q334 AND symb_decoder(16#54#)) OR
 					(reg_q334 AND symb_decoder(16#74#));
reg_q338_in <= (reg_q336 AND symb_decoder(16#41#)) OR
 					(reg_q336 AND symb_decoder(16#61#));
reg_q300_in <= (reg_q298 AND symb_decoder(16#64#)) OR
 					(reg_q298 AND symb_decoder(16#44#));
reg_q573_in <= (reg_q571 AND symb_decoder(16#2e#));
reg_q765_in <= (reg_q763 AND symb_decoder(16#72#)) OR
 					(reg_q763 AND symb_decoder(16#52#));
reg_q1264_in <= (reg_q1262 AND symb_decoder(16#64#)) OR
 					(reg_q1262 AND symb_decoder(16#44#));
reg_q610_in <= (reg_q608 AND symb_decoder(16#56#)) OR
 					(reg_q608 AND symb_decoder(16#76#));
reg_q1512_in <= (reg_q1510 AND symb_decoder(16#72#)) OR
 					(reg_q1510 AND symb_decoder(16#52#));
reg_q453_in <= (reg_q453 AND symb_decoder(16#0d#)) OR
 					(reg_q453 AND symb_decoder(16#20#)) OR
 					(reg_q453 AND symb_decoder(16#0a#)) OR
 					(reg_q453 AND symb_decoder(16#09#)) OR
 					(reg_q453 AND symb_decoder(16#0c#)) OR
 					(reg_q451 AND symb_decoder(16#20#)) OR
 					(reg_q451 AND symb_decoder(16#0a#)) OR
 					(reg_q451 AND symb_decoder(16#0c#)) OR
 					(reg_q451 AND symb_decoder(16#09#)) OR
 					(reg_q451 AND symb_decoder(16#0d#));
reg_q2491_in <= (reg_q2489 AND symb_decoder(16#41#)) OR
 					(reg_q2489 AND symb_decoder(16#61#));
reg_q1536_in <= (reg_q1534 AND symb_decoder(16#73#)) OR
 					(reg_q1534 AND symb_decoder(16#53#));
reg_q2202_in <= (reg_q2200 AND symb_decoder(16#46#)) OR
 					(reg_q2200 AND symb_decoder(16#66#));
reg_q2204_in <= (reg_q2202 AND symb_decoder(16#59#)) OR
 					(reg_q2202 AND symb_decoder(16#79#));
reg_q2663_in <= (reg_q2661 AND symb_decoder(16#69#)) OR
 					(reg_q2661 AND symb_decoder(16#49#));
reg_q2566_in <= (reg_q2564 AND symb_decoder(16#56#)) OR
 					(reg_q2564 AND symb_decoder(16#76#));
reg_q2580_in <= (reg_q2578 AND symb_decoder(16#5d#));
reg_q1959_in <= (reg_q1957 AND symb_decoder(16#2d#));
reg_q920_in <= (reg_q918 AND symb_decoder(16#41#)) OR
 					(reg_q918 AND symb_decoder(16#61#));
reg_q1654_in <= (reg_q1652 AND symb_decoder(16#74#)) OR
 					(reg_q1652 AND symb_decoder(16#54#));
reg_q1656_in <= (reg_q1654 AND symb_decoder(16#68#)) OR
 					(reg_q1654 AND symb_decoder(16#48#));
reg_q1224_in <= (reg_q1222 AND symb_decoder(16#6c#)) OR
 					(reg_q1222 AND symb_decoder(16#4c#));
reg_q2106_in <= (reg_q2104 AND symb_decoder(16#79#)) OR
 					(reg_q2104 AND symb_decoder(16#59#));
reg_q2182_in <= (reg_q2180 AND symb_decoder(16#45#)) OR
 					(reg_q2180 AND symb_decoder(16#65#));
reg_q1864_in <= (reg_q1862 AND symb_decoder(16#4f#)) OR
 					(reg_q1862 AND symb_decoder(16#6f#));
reg_q1586_in <= (reg_q1584 AND symb_decoder(16#63#)) OR
 					(reg_q1584 AND symb_decoder(16#43#));
reg_q2455_in <= (reg_q2453 AND symb_decoder(16#49#)) OR
 					(reg_q2453 AND symb_decoder(16#69#));
reg_q914_in <= (reg_q912 AND symb_decoder(16#75#)) OR
 					(reg_q912 AND symb_decoder(16#55#));
reg_q451_in <= (reg_q449 AND symb_decoder(16#64#)) OR
 					(reg_q449 AND symb_decoder(16#44#));
reg_q1556_in <= (reg_q1554 AND symb_decoder(16#59#)) OR
 					(reg_q1554 AND symb_decoder(16#79#));
reg_q2132_in <= (reg_q2130 AND symb_decoder(16#45#)) OR
 					(reg_q2130 AND symb_decoder(16#65#));
reg_q2134_in <= (reg_q2132 AND symb_decoder(16#3d#));
reg_q1417_in <= (reg_q1415 AND symb_decoder(16#53#)) OR
 					(reg_q1415 AND symb_decoder(16#73#));
reg_q1419_in <= (reg_q1417 AND symb_decoder(16#20#)) OR
 					(reg_q1417 AND symb_decoder(16#0c#)) OR
 					(reg_q1417 AND symb_decoder(16#0d#)) OR
 					(reg_q1417 AND symb_decoder(16#09#)) OR
 					(reg_q1417 AND symb_decoder(16#0a#)) OR
 					(reg_q1419 AND symb_decoder(16#0d#)) OR
 					(reg_q1419 AND symb_decoder(16#09#)) OR
 					(reg_q1419 AND symb_decoder(16#0a#)) OR
 					(reg_q1419 AND symb_decoder(16#20#)) OR
 					(reg_q1419 AND symb_decoder(16#0c#));
reg_q872_in <= (reg_q870 AND symb_decoder(16#63#)) OR
 					(reg_q870 AND symb_decoder(16#43#));
reg_q638_in <= (reg_q636 AND symb_decoder(16#6c#)) OR
 					(reg_q636 AND symb_decoder(16#4c#));
reg_q640_in <= (reg_q638 AND symb_decoder(16#69#)) OR
 					(reg_q638 AND symb_decoder(16#49#));
reg_q431_in <= (reg_q429 AND symb_decoder(16#45#)) OR
 					(reg_q429 AND symb_decoder(16#65#));
reg_q1646_in <= (reg_q1644 AND symb_decoder(16#44#)) OR
 					(reg_q1644 AND symb_decoder(16#64#));
reg_q1532_in <= (reg_q1530 AND symb_decoder(16#4f#)) OR
 					(reg_q1530 AND symb_decoder(16#6f#));
reg_q1624_in <= (reg_q1622 AND symb_decoder(16#3d#));
reg_q1292_in <= (reg_q1290 AND symb_decoder(16#52#)) OR
 					(reg_q1290 AND symb_decoder(16#72#));
reg_q1298_in <= (reg_q1296 AND symb_decoder(16#45#)) OR
 					(reg_q1296 AND symb_decoder(16#65#));
reg_q2196_in <= (reg_q2194 AND symb_decoder(16#4f#)) OR
 					(reg_q2194 AND symb_decoder(16#6f#));
reg_q936_in <= (reg_q934 AND symb_decoder(16#69#)) OR
 					(reg_q934 AND symb_decoder(16#49#));
reg_q938_in <= (reg_q936 AND symb_decoder(16#6e#)) OR
 					(reg_q936 AND symb_decoder(16#4e#));
reg_q1083_in <= (reg_q1081 AND symb_decoder(16#54#)) OR
 					(reg_q1081 AND symb_decoder(16#74#));
reg_q1403_in <= (reg_q1401 AND symb_decoder(16#47#)) OR
 					(reg_q1401 AND symb_decoder(16#67#));
reg_q2140_in <= (reg_q2138 AND symb_decoder(16#61#)) OR
 					(reg_q2138 AND symb_decoder(16#41#));
reg_q2142_in <= (reg_q2140 AND symb_decoder(16#2d#));
reg_q1886_in <= (reg_q1884 AND symb_decoder(16#23#));
reg_q1828_in <= (reg_q1826 AND symb_decoder(16#4f#)) OR
 					(reg_q1826 AND symb_decoder(16#6f#));
reg_q1830_in <= (reg_q1828 AND symb_decoder(16#4d#)) OR
 					(reg_q1828 AND symb_decoder(16#6d#));
reg_q2515_in <= (reg_q2513 AND symb_decoder(16#45#)) OR
 					(reg_q2513 AND symb_decoder(16#65#));
reg_q1381_in <= (reg_q1379 AND symb_decoder(16#44#)) OR
 					(reg_q1379 AND symb_decoder(16#64#));
reg_q1383_in <= (reg_q1381 AND symb_decoder(16#61#)) OR
 					(reg_q1381 AND symb_decoder(16#41#));
reg_q2489_in <= (reg_q2487 AND symb_decoder(16#6d#)) OR
 					(reg_q2487 AND symb_decoder(16#4d#));
reg_q650_in <= (reg_q648 AND symb_decoder(16#65#)) OR
 					(reg_q648 AND symb_decoder(16#45#));
reg_q744_in <= (reg_q742 AND symb_decoder(16#72#)) OR
 					(reg_q742 AND symb_decoder(16#52#));
reg_q1953_in <= (reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q1951 AND symb_decoder(16#2b#));
reg_q581_in <= (reg_q579 AND symb_decoder(16#2e#));
reg_q1542_in <= (reg_q1540 AND symb_decoder(16#69#)) OR
 					(reg_q1540 AND symb_decoder(16#49#));
reg_q1544_in <= (reg_q1542 AND symb_decoder(16#72#)) OR
 					(reg_q1542 AND symb_decoder(16#52#));
reg_q1842_in <= (reg_q1840 AND symb_decoder(16#52#)) OR
 					(reg_q1840 AND symb_decoder(16#72#));
reg_q2443_in <= (reg_q2441 AND symb_decoder(16#74#)) OR
 					(reg_q2441 AND symb_decoder(16#54#));
reg_q618_in <= (reg_q616 AND symb_decoder(16#6f#)) OR
 					(reg_q616 AND symb_decoder(16#4f#));
reg_q1413_in <= (reg_q1411 AND symb_decoder(16#68#)) OR
 					(reg_q1411 AND symb_decoder(16#48#));
reg_q1415_in <= (reg_q1413 AND symb_decoder(16#49#)) OR
 					(reg_q1413 AND symb_decoder(16#69#));
reg_q2548_in <= (reg_q2546 AND symb_decoder(16#3e#));
reg_q1040_in <= (reg_q1038 AND symb_decoder(16#54#));
reg_q2096_in <= (reg_q2094 AND symb_decoder(16#48#)) OR
 					(reg_q2094 AND symb_decoder(16#68#));
reg_q2098_in <= (reg_q2096 AND symb_decoder(16#41#)) OR
 					(reg_q2096 AND symb_decoder(16#61#));
reg_q827_in <= (reg_q825 AND symb_decoder(16#0c#)) OR
 					(reg_q825 AND symb_decoder(16#20#)) OR
 					(reg_q825 AND symb_decoder(16#0a#)) OR
 					(reg_q825 AND symb_decoder(16#0d#)) OR
 					(reg_q825 AND symb_decoder(16#09#)) OR
 					(reg_q827 AND symb_decoder(16#0c#)) OR
 					(reg_q827 AND symb_decoder(16#09#)) OR
 					(reg_q827 AND symb_decoder(16#0d#)) OR
 					(reg_q827 AND symb_decoder(16#0a#)) OR
 					(reg_q827 AND symb_decoder(16#20#));
reg_q1151_in <= (reg_q1149 AND symb_decoder(16#52#)) OR
 					(reg_q1149 AND symb_decoder(16#72#));
reg_q2144_in <= (reg_q2142 AND symb_decoder(16#54#)) OR
 					(reg_q2142 AND symb_decoder(16#74#));
reg_q888_in <= (reg_q886 AND symb_decoder(16#75#)) OR
 					(reg_q886 AND symb_decoder(16#55#));
reg_q616_in <= (reg_q614 AND symb_decoder(16#46#)) OR
 					(reg_q614 AND symb_decoder(16#66#));
reg_q1608_in <= (reg_q1606 AND symb_decoder(16#2e#));
reg_q1294_in <= (reg_q1292 AND symb_decoder(16#0c#)) OR
 					(reg_q1292 AND symb_decoder(16#20#)) OR
 					(reg_q1292 AND symb_decoder(16#0a#)) OR
 					(reg_q1292 AND symb_decoder(16#0d#)) OR
 					(reg_q1292 AND symb_decoder(16#09#)) OR
 					(reg_q1294 AND symb_decoder(16#0a#)) OR
 					(reg_q1294 AND symb_decoder(16#0d#)) OR
 					(reg_q1294 AND symb_decoder(16#0c#)) OR
 					(reg_q1294 AND symb_decoder(16#20#)) OR
 					(reg_q1294 AND symb_decoder(16#09#));
reg_q1240_in <= (reg_q1238 AND symb_decoder(16#0a#)) OR
 					(reg_q1238 AND symb_decoder(16#09#)) OR
 					(reg_q1238 AND symb_decoder(16#20#)) OR
 					(reg_q1238 AND symb_decoder(16#0d#)) OR
 					(reg_q1238 AND symb_decoder(16#0c#)) OR
 					(reg_q1240 AND symb_decoder(16#0a#)) OR
 					(reg_q1240 AND symb_decoder(16#0d#)) OR
 					(reg_q1240 AND symb_decoder(16#20#)) OR
 					(reg_q1240 AND symb_decoder(16#0c#)) OR
 					(reg_q1240 AND symb_decoder(16#09#));
reg_q658_in <= (reg_q656 AND symb_decoder(16#52#)) OR
 					(reg_q656 AND symb_decoder(16#72#));
reg_q886_in <= (reg_q884 AND symb_decoder(16#42#)) OR
 					(reg_q884 AND symb_decoder(16#62#));
reg_q1894_in <= (reg_q1892 AND symb_decoder(16#23#));
reg_q2445_in <= (reg_q2443 AND symb_decoder(16#3e#));
reg_q2138_in <= (reg_q2136 AND symb_decoder(16#49#)) OR
 					(reg_q2136 AND symb_decoder(16#69#));
reg_q2485_in <= (reg_q2485 AND symb_decoder(16#0a#)) OR
 					(reg_q2485 AND symb_decoder(16#09#)) OR
 					(reg_q2485 AND symb_decoder(16#0c#)) OR
 					(reg_q2485 AND symb_decoder(16#20#)) OR
 					(reg_q2485 AND symb_decoder(16#0d#)) OR
 					(reg_q2483 AND symb_decoder(16#0d#)) OR
 					(reg_q2483 AND symb_decoder(16#20#)) OR
 					(reg_q2483 AND symb_decoder(16#0c#)) OR
 					(reg_q2483 AND symb_decoder(16#0a#)) OR
 					(reg_q2483 AND symb_decoder(16#09#));
reg_q1564_in <= (reg_q1562 AND symb_decoder(16#6f#)) OR
 					(reg_q1562 AND symb_decoder(16#4f#));
reg_q1566_in <= (reg_q1564 AND symb_decoder(16#6f#)) OR
 					(reg_q1564 AND symb_decoder(16#4f#));
reg_q1862_in <= (reg_q1860 AND symb_decoder(16#63#)) OR
 					(reg_q1860 AND symb_decoder(16#43#));
reg_q443_in <= (reg_q441 AND symb_decoder(16#42#)) OR
 					(reg_q441 AND symb_decoder(16#62#));
reg_q2210_in <= (reg_q2208 AND symb_decoder(16#45#)) OR
 					(reg_q2208 AND symb_decoder(16#65#));
reg_q447_in <= (reg_q445 AND symb_decoder(16#73#)) OR
 					(reg_q445 AND symb_decoder(16#53#));
reg_q449_in <= (reg_q447 AND symb_decoder(16#45#)) OR
 					(reg_q447 AND symb_decoder(16#65#));
reg_q1840_in <= (reg_q1838 AND symb_decoder(16#41#)) OR
 					(reg_q1838 AND symb_decoder(16#61#));
reg_q1824_in <= (reg_q1822 AND symb_decoder(16#41#)) OR
 					(reg_q1822 AND symb_decoder(16#61#));
reg_q1774_in <= (reg_q1772 AND symb_decoder(16#65#)) OR
 					(reg_q1772 AND symb_decoder(16#45#));
reg_q720_in <= (reg_q718 AND symb_decoder(16#54#)) OR
 					(reg_q718 AND symb_decoder(16#74#));
reg_q2483_in <= (reg_q2481 AND symb_decoder(16#59#)) OR
 					(reg_q2481 AND symb_decoder(16#79#));
reg_q2481_in <= (reg_q2479 AND symb_decoder(16#42#)) OR
 					(reg_q2479 AND symb_decoder(16#62#));
reg_q1568_in <= (reg_q1566 AND symb_decoder(16#64#)) OR
 					(reg_q1566 AND symb_decoder(16#44#));
reg_q2128_in <= (reg_q2126 AND symb_decoder(16#61#)) OR
 					(reg_q2126 AND symb_decoder(16#41#));
reg_q1666_in <= (reg_q1664 AND symb_decoder(16#70#)) OR
 					(reg_q1664 AND symb_decoder(16#50#));
reg_q2517_in <= (reg_q2515 AND symb_decoder(16#3e#));
reg_q391_in <= (reg_q389 AND symb_decoder(16#72#)) OR
 					(reg_q389 AND symb_decoder(16#52#));
reg_q796_in <= (reg_q794 AND symb_decoder(16#34#));
reg_q798_in <= (reg_q796 AND symb_decoder(16#31#));
reg_q1878_in <= (reg_q1876 AND symb_decoder(16#4f#)) OR
 					(reg_q1876 AND symb_decoder(16#6f#));
reg_q1880_in <= (reg_q1878 AND symb_decoder(16#61#)) OR
 					(reg_q1878 AND symb_decoder(16#41#));
reg_q2499_in <= (reg_q2497 AND symb_decoder(16#66#)) OR
 					(reg_q2497 AND symb_decoder(16#46#));
reg_q2086_in <= (reg_q2084 AND symb_decoder(16#61#)) OR
 					(reg_q2084 AND symb_decoder(16#41#));
reg_q2180_in <= (reg_q2178 AND symb_decoder(16#6d#)) OR
 					(reg_q2178 AND symb_decoder(16#4d#));
reg_q421_in <= (reg_q419 AND symb_decoder(16#72#)) OR
 					(reg_q419 AND symb_decoder(16#52#));
reg_q2136_in <= (reg_q2134 AND symb_decoder(16#43#)) OR
 					(reg_q2134 AND symb_decoder(16#63#));
reg_q2507_in <= (reg_q2505 AND symb_decoder(16#74#)) OR
 					(reg_q2505 AND symb_decoder(16#54#));
reg_q2399_in <= (reg_q2361 AND symb_decoder(16#61#)) OR
 					(reg_q2361 AND symb_decoder(16#41#));
reg_q2501_in <= (reg_q2499 AND symb_decoder(16#74#)) OR
 					(reg_q2499 AND symb_decoder(16#54#));
reg_q304_in <= (reg_q302 AND symb_decoder(16#65#)) OR
 					(reg_q302 AND symb_decoder(16#45#));
reg_q2100_in <= (reg_q2098 AND symb_decoder(16#6e#)) OR
 					(reg_q2098 AND symb_decoder(16#4e#));
reg_q1664_in <= (reg_q1662 AND symb_decoder(16#2e#));
reg_q896_in <= (reg_q894 AND symb_decoder(16#45#)) OR
 					(reg_q894 AND symb_decoder(16#65#));
reg_q2675_in <= (reg_q2673 AND symb_decoder(16#7c#));
reg_q429_in <= (reg_q427 AND symb_decoder(16#74#)) OR
 					(reg_q427 AND symb_decoder(16#54#));
reg_q2657_in <= (reg_q2655 AND symb_decoder(16#59#)) OR
 					(reg_q2655 AND symb_decoder(16#79#));
reg_q2461_in <= (reg_q2459 AND symb_decoder(16#45#)) OR
 					(reg_q2459 AND symb_decoder(16#65#));
reg_q1226_in <= (reg_q1224 AND symb_decoder(16#63#)) OR
 					(reg_q1224 AND symb_decoder(16#43#));
reg_q1228_in <= (reg_q1226 AND symb_decoder(16#4f#)) OR
 					(reg_q1226 AND symb_decoder(16#6f#));
reg_q642_in <= (reg_q640 AND symb_decoder(16#74#)) OR
 					(reg_q640 AND symb_decoder(16#54#));
reg_q302_in <= (reg_q300 AND symb_decoder(16#6c#)) OR
 					(reg_q300 AND symb_decoder(16#4c#));
reg_q1939_in <= (reg_q1937 AND symb_decoder(16#4f#));
reg_q2425_in <= (reg_q2423 AND symb_decoder(16#41#)) OR
 					(reg_q2423 AND symb_decoder(16#61#));
reg_q2427_in <= (reg_q2425 AND symb_decoder(16#54#)) OR
 					(reg_q2425 AND symb_decoder(16#74#));
reg_q1054_in <= (reg_q1052 AND symb_decoder(16#65#));
reg_q1056_in <= (reg_q1054 AND symb_decoder(16#72#));
reg_q1826_in <= (reg_q1824 AND symb_decoder(16#43#)) OR
 					(reg_q1824 AND symb_decoder(16#63#));
reg_q1302_in <= (reg_q1300 AND symb_decoder(16#76#)) OR
 					(reg_q1300 AND symb_decoder(16#56#));
reg_q1268_in <= (reg_q1266 AND symb_decoder(16#66#)) OR
 					(reg_q1266 AND symb_decoder(16#46#));
reg_q1874_in <= (reg_q1872 AND symb_decoder(16#61#)) OR
 					(reg_q1872 AND symb_decoder(16#41#));
reg_q2574_in <= (reg_q2572 AND symb_decoder(16#69#)) OR
 					(reg_q2572 AND symb_decoder(16#49#));
reg_q467_in <= (reg_q465 AND symb_decoder(16#45#)) OR
 					(reg_q465 AND symb_decoder(16#65#));
reg_q1510_in <= (reg_q1508 AND symb_decoder(16#45#)) OR
 					(reg_q1508 AND symb_decoder(16#65#));
reg_q1199_in <= (reg_q1197 AND symb_decoder(16#45#)) OR
 					(reg_q1197 AND symb_decoder(16#65#));
reg_q1201_in <= (reg_q1199 AND symb_decoder(16#52#)) OR
 					(reg_q1199 AND symb_decoder(16#72#));
reg_q1876_in <= (reg_q1874 AND symb_decoder(16#44#)) OR
 					(reg_q1874 AND symb_decoder(16#64#));
reg_q1435_in <= (reg_q1433 AND symb_decoder(16#41#)) OR
 					(reg_q1433 AND symb_decoder(16#61#));
reg_q1437_in <= (reg_q1435 AND symb_decoder(16#45#)) OR
 					(reg_q1435 AND symb_decoder(16#65#));
reg_q833_in <= (reg_q831 AND symb_decoder(16#6c#)) OR
 					(reg_q831 AND symb_decoder(16#4c#));
reg_q445_in <= (reg_q443 AND symb_decoder(16#41#)) OR
 					(reg_q443 AND symb_decoder(16#61#));
reg_q780_in <= (reg_q778 AND symb_decoder(16#6a#)) OR
 					(reg_q778 AND symb_decoder(16#4a#));
reg_q2463_in <= (reg_q2461 AND symb_decoder(16#3e#));
reg_q409_in <= (reg_q407 AND symb_decoder(16#4f#)) OR
 					(reg_q407 AND symb_decoder(16#6f#));
reg_q1920_in <= (reg_q1918 AND symb_decoder(16#50#));
reg_q829_in <= (reg_q827 AND symb_decoder(16#6f#)) OR
 					(reg_q827 AND symb_decoder(16#4f#));
reg_q831_in <= (reg_q829 AND symb_decoder(16#6e#)) OR
 					(reg_q829 AND symb_decoder(16#4e#));
reg_q1439_in <= (reg_q1437 AND symb_decoder(16#4d#)) OR
 					(reg_q1437 AND symb_decoder(16#6d#));
reg_q1441_in <= (reg_q1439 AND symb_decoder(16#6f#)) OR
 					(reg_q1439 AND symb_decoder(16#4f#));
reg_q1678_in <= (reg_q1676 AND symb_decoder(16#7a#)) OR
 					(reg_q1676 AND symb_decoder(16#5a#));
reg_q1038_in <= (reg_q1036 AND symb_decoder(16#46#));
reg_q2068_in <= (reg_q2066 AND symb_decoder(16#6e#)) OR
 					(reg_q2066 AND symb_decoder(16#4e#));
reg_q1048_in <= (reg_q1046 AND symb_decoder(16#65#));
reg_q1050_in <= (reg_q1048 AND symb_decoder(16#72#));
reg_q2130_in <= (reg_q2128 AND symb_decoder(16#6d#)) OR
 					(reg_q2128 AND symb_decoder(16#4d#));
reg_q2166_in <= (reg_q2164 AND symb_decoder(16#5f#));
reg_q324_in <= (reg_q322 AND symb_decoder(16#72#)) OR
 					(reg_q322 AND symb_decoder(16#52#));
reg_q1882_in <= (reg_q1880 AND symb_decoder(16#23#));
reg_q2669_in <= (reg_q2667 AND symb_decoder(16#31#));
reg_q2102_in <= (reg_q2100 AND symb_decoder(16#6b#)) OR
 					(reg_q2100 AND symb_decoder(16#4b#));
reg_q908_in <= (reg_q906 AND symb_decoder(16#69#)) OR
 					(reg_q906 AND symb_decoder(16#49#));
reg_q1149_in <= (reg_q1147 AND symb_decoder(16#45#)) OR
 					(reg_q1147 AND symb_decoder(16#65#));
reg_q2104_in <= (reg_q2102 AND symb_decoder(16#5f#));
reg_q1838_in <= (reg_q1836 AND symb_decoder(16#62#)) OR
 					(reg_q1836 AND symb_decoder(16#42#));
reg_q1896_in <= (reg_q1894 AND symb_decoder(16#46#)) OR
 					(reg_q1894 AND symb_decoder(16#66#));
reg_q1772_in <= (reg_q1770 AND symb_decoder(16#52#)) OR
 					(reg_q1770 AND symb_decoder(16#72#));
reg_q1433_in <= (reg_q1431 AND symb_decoder(16#64#)) OR
 					(reg_q1431 AND symb_decoder(16#44#));
reg_q1554_in <= (reg_q1552 AND symb_decoder(16#52#)) OR
 					(reg_q1552 AND symb_decoder(16#72#));
reg_q940_in <= (reg_q938 AND symb_decoder(16#47#)) OR
 					(reg_q938 AND symb_decoder(16#67#));
reg_q1300_in <= (reg_q1298 AND symb_decoder(16#52#)) OR
 					(reg_q1298 AND symb_decoder(16#72#));
reg_q1836_in <= (reg_q1834 AND symb_decoder(16#6f#)) OR
 					(reg_q1834 AND symb_decoder(16#4f#));
reg_q2546_in <= (reg_q2544 AND symb_decoder(16#5c#));
reg_q902_in <= (reg_q900 AND symb_decoder(16#45#)) OR
 					(reg_q900 AND symb_decoder(16#65#));
reg_q1680_in <= (reg_q1678 AND symb_decoder(16#3d#));
reg_q1030_in <= (reg_q1028 AND symb_decoder(16#65#));
reg_q1032_in <= (reg_q1030 AND symb_decoder(16#66#));
reg_q1052_in <= (reg_q1050 AND symb_decoder(16#76#));
reg_q1898_in <= (reg_q1896 AND symb_decoder(16#23#));
reg_q1058_in <= (reg_q1056 AND symb_decoder(16#3a#));
reg_q427_in <= (reg_q425 AND symb_decoder(16#6f#)) OR
 					(reg_q425 AND symb_decoder(16#4f#));
reg_q2544_in <= (reg_q2542 AND symb_decoder(16#24#));
reg_fullgraph5_init <= "000000000";

reg_fullgraph5_sel <= "00000000000000000000" & reg_q2544_in & reg_q427_in & reg_q1058_in & reg_q1898_in & reg_q1052_in & reg_q1032_in & reg_q1030_in & reg_q1680_in & reg_q902_in & reg_q2546_in & reg_q1836_in & reg_q1300_in & reg_q940_in & reg_q1554_in & reg_q1433_in & reg_q1772_in & reg_q1896_in & reg_q1838_in & reg_q2104_in & reg_q1149_in & reg_q908_in & reg_q2102_in & reg_q2669_in & reg_q1882_in & reg_q324_in & reg_q2166_in & reg_q2130_in & reg_q1050_in & reg_q1048_in & reg_q2068_in & reg_q1038_in & reg_q1678_in & reg_q1441_in & reg_q1439_in & reg_q831_in & reg_q829_in & reg_q1920_in & reg_q409_in & reg_q2463_in & reg_q780_in & reg_q445_in & reg_q833_in & reg_q1437_in & reg_q1435_in & reg_q1876_in & reg_q1201_in & reg_q1199_in & reg_q1510_in & reg_q467_in & reg_q2574_in & reg_q1874_in & reg_q1268_in & reg_q1302_in & reg_q1826_in & reg_q1056_in & reg_q1054_in & reg_q2427_in & reg_q2425_in & reg_q1939_in & reg_q302_in & reg_q642_in & reg_q1228_in & reg_q1226_in & reg_q2461_in & reg_q2657_in & reg_q429_in & reg_q2675_in & reg_q896_in & reg_q1664_in & reg_q2100_in & reg_q304_in & reg_q2501_in & reg_q2399_in & reg_q2507_in & reg_q2136_in & reg_q421_in & reg_q2180_in & reg_q2086_in & reg_q2499_in & reg_q1880_in & reg_q1878_in & reg_q798_in & reg_q796_in & reg_q391_in & reg_q2517_in & reg_q1666_in & reg_q2128_in & reg_q1568_in & reg_q2481_in & reg_q2483_in & reg_q720_in & reg_q1774_in & reg_q1824_in & reg_q1840_in & reg_q449_in & reg_q447_in & reg_q2210_in & reg_q443_in & reg_q1862_in & reg_q1566_in & reg_q1564_in & reg_q2485_in & reg_q2138_in & reg_q2445_in & reg_q1894_in & reg_q886_in & reg_q658_in & reg_q1240_in & reg_q1294_in & reg_q1608_in & reg_q616_in & reg_q888_in & reg_q2144_in & reg_q1151_in & reg_q827_in & reg_q2098_in & reg_q2096_in & reg_q1040_in & reg_q2548_in & reg_q1415_in & reg_q1413_in & reg_q618_in & reg_q2443_in & reg_q1842_in & reg_q1544_in & reg_q1542_in & reg_q581_in & reg_q1953_in & reg_q744_in & reg_q650_in & reg_q2489_in & reg_q1383_in & reg_q1381_in & reg_q2515_in & reg_q1830_in & reg_q1828_in & reg_q1886_in & reg_q2142_in & reg_q2140_in & reg_q1403_in & reg_q1083_in & reg_q938_in & reg_q936_in & reg_q2196_in & reg_q1298_in & reg_q1292_in & reg_q1624_in & reg_q1532_in & reg_q1646_in & reg_q431_in & reg_q640_in & reg_q638_in & reg_q872_in & reg_q1419_in & reg_q1417_in & reg_q2134_in & reg_q2132_in & reg_q1556_in & reg_q451_in & reg_q914_in & reg_q2455_in & reg_q1586_in & reg_q1864_in & reg_q2182_in & reg_q2106_in & reg_q1224_in & reg_q1656_in & reg_q1654_in & reg_q920_in & reg_q1959_in & reg_q2580_in & reg_q2566_in & reg_q2663_in & reg_q2204_in & reg_q2202_in & reg_q1536_in & reg_q2491_in & reg_q453_in & reg_q1512_in & reg_q610_in & reg_q1264_in & reg_q765_in & reg_q573_in & reg_q300_in & reg_q338_in & reg_q336_in & reg_q1562_in & reg_q1560_in & reg_q459_in & reg_q457_in & reg_q1901_in & reg_q2475_in & reg_q322_in & reg_q320_in & reg_q465_in & reg_q463_in & reg_q2459_in & reg_q2457_in & reg_q922_in & reg_q1238_in & reg_q1957_in & reg_q1955_in & reg_q2084_in & reg_q1282_in & reg_q2174_in & reg_q306_in & reg_q1632_in & reg_q2477_in & reg_q2740_in & reg_q2564_in & reg_q407_in & reg_q405_in & reg_q413_in & reg_q577_in & reg_q1971_in & reg_q1969_in & reg_q1872_in & reg_q1870_in & reg_q2513_in & reg_q1306_in & reg_q1304_in & reg_q1868_in & reg_q1866_in & reg_q1967_in & reg_q1638_in & reg_q2667_in & reg_q2665_in & reg_q1367_in & reg_q1907_in & reg_q934_in & reg_q932_in & reg_q579_in & reg_q2423_in & reg_q2421_in & reg_q2742_in & reg_q1246_in & reg_q1471_in & reg_q326_in & reg_q2473_in & reg_q2471_in & reg_q1888_in & reg_q1401_in & reg_q1650_in & reg_q1648_in & reg_q2208_in & reg_q2206_in & reg_q825_in & reg_q614_in & reg_q612_in & reg_q1733_in & reg_q1731_in & reg_q1852_in & reg_q1850_in & reg_q1286_in & reg_q1284_in & reg_q2671_in & reg_q742_in & reg_q1552_in & reg_q1550_in & reg_q1540_in & reg_q1538_in & reg_q1036_in & reg_q1236_in & reg_q2120_in & reg_q1662_in & reg_q1822_in & reg_q433_in & reg_q2497_in & reg_q866_in & reg_q864_in & reg_q2186_in & reg_q2184_in & reg_q870_in & reg_q2066_in & reg_q2090_in & reg_q2088_in & reg_q924_in & reg_q2465_in & reg_q2158_in & reg_q2156_in & reg_q1244_in & reg_q1242_in & reg_q2072_in & reg_q2070_in & reg_q2178_in & reg_q2176_in & reg_q910_in & reg_q2542_in & reg_q2540_in & reg_q656_in & reg_q1280_in & reg_q1278_in & reg_q1138_in & reg_q1256_in & reg_q1254_in & reg_q1455_in & reg_q632_in & reg_q630_in & reg_q900_in & reg_q898_in & reg_q2188_in & reg_q403_in & reg_q549_in & reg_q1325_in & reg_q926_in & reg_q2148_in & reg_q2146_in & reg_q503_in & reg_q2200_in & reg_q2198_in & reg_q930_in & reg_q928_in & reg_q2532_in & reg_q2530_in & reg_q1614_in & reg_q1272_in & reg_q912_in & reg_q1421_in & reg_q839_in & reg_q1409_in & reg_q654_in & reg_q652_in & reg_q841_in & reg_q1582_in & reg_q1580_in & reg_q1572_in & reg_q1570_in & reg_q1670_in & reg_q1668_in & reg_q1558_in & reg_q1258_in & reg_q628_in & reg_q626_in & reg_q837_in & reg_q835_in & reg_q1451_in & reg_q1449_in & reg_q2558_in & reg_q2126_in & reg_q2124_in & reg_q334_in & reg_q585_in & reg_q181_in & reg_q1248_in & reg_q2078_in & reg_q2076_in & reg_q332_in & reg_q1590_in & reg_q1588_in & reg_q425_in & reg_q423_in & reg_q624_in & reg_q1622_in & reg_q340_in & reg_q1290_in & reg_q1288_in & reg_q2214_in & reg_q2212_in & reg_q1425_in & reg_q1423_in & reg_q1252_in & reg_q1250_in & reg_q1230_in & reg_q1477_in & reg_q1234_in & reg_q1232_in & reg_q1943_in & reg_q2469_in & reg_q2467_in & reg_q918_in & reg_q916_in & reg_q1407_in & reg_q1405_in & reg_q1375_in & reg_q2493_in & reg_q1276_in & reg_q1274_in & reg_q2661_in & reg_q2659_in & reg_q786_in & reg_q1373_in & reg_q1371_in & reg_q2110_in & reg_q2108_in & reg_q1266_in & reg_q417_in & reg_q415_in & reg_q419_in & reg_q1431_in & reg_q2568_in & reg_q583_in & reg_q2170_in & reg_q2168_in & reg_q2562_in & reg_q2560_in & reg_q1600_in & reg_q2190_in & reg_q330_in & reg_q328_in & reg_q437_in & reg_q1856_in & reg_q1854_in & reg_q1548_in & reg_q1546_in & reg_q767_in & reg_q1612_in & reg_q1610_in & reg_q1834_in & reg_q1832_in & reg_q862_in & reg_q906_in & reg_q904_in & reg_q1429_in & reg_q1427_in & reg_q575_in & reg_q1262_in & reg_q1260_in & reg_q1475_in & reg_q1473_in & reg_q2437_in & reg_q292_in & reg_q290_in & reg_q1860_in & reg_q1858_in & reg_q2511_in & reg_q2509_in & reg_q183_in & reg_q892_in & reg_q890_in & reg_q1844_in & reg_q1528_in & reg_q1526_in & reg_q2479_in & reg_q314_in & reg_q312_in & reg_q1606_in & reg_q794_in & reg_q792_in & reg_q1660_in & reg_q1658_in & reg_q608_in & reg_q2235_in & reg_q1044_in & reg_q1042_in & reg_q2578_in & reg_q2576_in & reg_q173_in & reg_q490_in & reg_q488_in & reg_q441_in & reg_q439_in & reg_q2094_in & reg_q2092_in & reg_q1524_in & reg_q2194_in & reg_q2192_in & reg_q2441_in & reg_q2439_in & reg_q2112_in & reg_q1616_in & reg_q622_in & reg_q620_in & reg_q318_in & reg_q316_in & reg_q2150_in & reg_q2627_in & reg_q2082_in & reg_q1892_in & reg_q1890_in & reg_q2534_in & reg_q1379_in & reg_q1377_in & reg_q819_in & reg_q2453_in & reg_q2451_in & reg_q2572_in & reg_q2570_in & reg_q636_in & reg_q634_in & reg_q179_in & reg_q646_in & reg_q644_in & reg_q1443_in & reg_q2651_in & reg_q308_in & reg_q1604_in & reg_q1602_in & reg_q2429_in & reg_q1672_in & reg_q1961_in & reg_q2233_in & reg_q2231_in;

	--coder fullgraph5
with reg_fullgraph5_sel select
reg_fullgraph5_in <=
	"000000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001",
	"000000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010",
	"000000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100",
	"000000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000",
	"000000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000",
	"000000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000",
	"000000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000",
	"000001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000",
	"000001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
	"000001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000",
	"000001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000",
	"000001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000",
	"000001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000",
	"000001110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000",
	"000001111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000",
	"000010000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000",
	"000010001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000",
	"000010010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000",
	"000010011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000",
	"000010100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000",
	"000010101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000",
	"000010110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000",
	"000010111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000",
	"000011000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000",
	"000011001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000",
	"000011010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000",
	"000011011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000",
	"000011100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000",
	"000011101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000",
	"000011110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000",
	"000011111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000",
	"000100000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000",
	"000100001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000",
	"000100010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000",
	"000100011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000",
	"000100100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000",
	"000100101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000",
	"000100110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000",
	"000100111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000",
	"000101000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000",
	"000101001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000",
	"000101010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000",
	"000101011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000",
	"000101100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000",
	"000101101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"000101110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000",
	"000101111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000",
	"000110000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000",
	"000110001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000",
	"000110010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000",
	"000110011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000",
	"000110100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000",
	"000110101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000",
	"000110110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000",
	"000110111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000",
	"000111000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000",
	"000111001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000",
	"000111010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000",
	"000111011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000",
	"000111100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000",
	"000111101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000",
	"000111110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000",
	"000111111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000",
	"001000000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000",
	"001000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000",
	"001000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000",
	"001000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000",
	"001000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000",
	"001000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000",
	"001000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000",
	"001000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000",
	"001001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000",
	"001001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000",
	"001001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000",
	"001001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000",
	"001001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001001110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001001111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101010000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101010001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101010010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101010011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101010100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101010101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101010110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101010111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101011000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101011001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101011010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101011011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101011100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101011101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101011110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101011111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101100000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101100001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101100010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101100011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101100100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101100101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101100110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101100111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101101000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101101001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101101010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101101011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101101100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101101101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101101110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101101111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101110000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101110001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101110010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101110011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101110100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101110101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101110110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101110111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101111000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101111001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101111010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101111011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101111100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101111101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101111110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101111111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110000000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110001110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110001111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110010000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110010001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110010010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110010011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110010100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110010101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110010110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110010111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110011000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110011001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110011010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110011011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110011100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110011101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110011110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110011111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110100000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110100001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110100010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110100011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110100100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110100101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110100110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110100111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110101000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110101001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110101010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110101011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110101100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110101101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110101110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110101111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110110000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110110001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110110010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110110011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110110100" when "00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110110101" when "00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110110110" when "00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110110111" when "00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110111000" when "00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110111001" when "00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110111010" when "00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110111011" when "00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110111100" when "00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110111101" when "00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110111110" when "00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"110111111" when "00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111000000" when "00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111000001" when "00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111000010" when "00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111000011" when "00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111000100" when "00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111000101" when "00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111000110" when "00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111000111" when "00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111001000" when "00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111001001" when "00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111001010" when "00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111001011" when "00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111001100" when "00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111001101" when "00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111001110" when "00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111001111" when "00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111010000" when "00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111010001" when "00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111010010" when "00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111010011" when "00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111010100" when "00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111010101" when "00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111010110" when "00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111010111" when "00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111011000" when "00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111011001" when "00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111011010" when "00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111011011" when "00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111011100" when "00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111011101" when "00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111011110" when "00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111011111" when "00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111100000" when "00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111100001" when "00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111100010" when "00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111100011" when "00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111100100" when "00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111100101" when "00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111100110" when "00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111100111" when "00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111101000" when "00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111101001" when "00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111101010" when "00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111101011" when "00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"111101100" when "00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"000000000" when others;
 --end coder

	p_reg_fullgraph5: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph5 <= reg_fullgraph5_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph5 <= reg_fullgraph5_init;
        else
          reg_fullgraph5 <= reg_fullgraph5_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph5

		reg_q2231 <= '1' when reg_fullgraph5 = "000000001" else '0'; 
		reg_q2233 <= '1' when reg_fullgraph5 = "000000010" else '0'; 
		reg_q1961 <= '1' when reg_fullgraph5 = "000000011" else '0'; 
		reg_q1672 <= '1' when reg_fullgraph5 = "000000100" else '0'; 
		reg_q2429 <= '1' when reg_fullgraph5 = "000000101" else '0'; 
		reg_q1602 <= '1' when reg_fullgraph5 = "000000110" else '0'; 
		reg_q1604 <= '1' when reg_fullgraph5 = "000000111" else '0'; 
		reg_q308 <= '1' when reg_fullgraph5 = "000001000" else '0'; 
		reg_q2651 <= '1' when reg_fullgraph5 = "000001001" else '0'; 
		reg_q1443 <= '1' when reg_fullgraph5 = "000001010" else '0'; 
		reg_q644 <= '1' when reg_fullgraph5 = "000001011" else '0'; 
		reg_q646 <= '1' when reg_fullgraph5 = "000001100" else '0'; 
		reg_q179 <= '1' when reg_fullgraph5 = "000001101" else '0'; 
		reg_q634 <= '1' when reg_fullgraph5 = "000001110" else '0'; 
		reg_q636 <= '1' when reg_fullgraph5 = "000001111" else '0'; 
		reg_q2570 <= '1' when reg_fullgraph5 = "000010000" else '0'; 
		reg_q2572 <= '1' when reg_fullgraph5 = "000010001" else '0'; 
		reg_q2451 <= '1' when reg_fullgraph5 = "000010010" else '0'; 
		reg_q2453 <= '1' when reg_fullgraph5 = "000010011" else '0'; 
		reg_q819 <= '1' when reg_fullgraph5 = "000010100" else '0'; 
		reg_q1377 <= '1' when reg_fullgraph5 = "000010101" else '0'; 
		reg_q1379 <= '1' when reg_fullgraph5 = "000010110" else '0'; 
		reg_q2534 <= '1' when reg_fullgraph5 = "000010111" else '0'; 
		reg_q1890 <= '1' when reg_fullgraph5 = "000011000" else '0'; 
		reg_q1892 <= '1' when reg_fullgraph5 = "000011001" else '0'; 
		reg_q2082 <= '1' when reg_fullgraph5 = "000011010" else '0'; 
		reg_q2627 <= '1' when reg_fullgraph5 = "000011011" else '0'; 
		reg_q2150 <= '1' when reg_fullgraph5 = "000011100" else '0'; 
		reg_q316 <= '1' when reg_fullgraph5 = "000011101" else '0'; 
		reg_q318 <= '1' when reg_fullgraph5 = "000011110" else '0'; 
		reg_q620 <= '1' when reg_fullgraph5 = "000011111" else '0'; 
		reg_q622 <= '1' when reg_fullgraph5 = "000100000" else '0'; 
		reg_q1616 <= '1' when reg_fullgraph5 = "000100001" else '0'; 
		reg_q2112 <= '1' when reg_fullgraph5 = "000100010" else '0'; 
		reg_q2439 <= '1' when reg_fullgraph5 = "000100011" else '0'; 
		reg_q2441 <= '1' when reg_fullgraph5 = "000100100" else '0'; 
		reg_q2192 <= '1' when reg_fullgraph5 = "000100101" else '0'; 
		reg_q2194 <= '1' when reg_fullgraph5 = "000100110" else '0'; 
		reg_q1524 <= '1' when reg_fullgraph5 = "000100111" else '0'; 
		reg_q2092 <= '1' when reg_fullgraph5 = "000101000" else '0'; 
		reg_q2094 <= '1' when reg_fullgraph5 = "000101001" else '0'; 
		reg_q439 <= '1' when reg_fullgraph5 = "000101010" else '0'; 
		reg_q441 <= '1' when reg_fullgraph5 = "000101011" else '0'; 
		reg_q488 <= '1' when reg_fullgraph5 = "000101100" else '0'; 
		reg_q490 <= '1' when reg_fullgraph5 = "000101101" else '0'; 
		reg_q173 <= '1' when reg_fullgraph5 = "000101110" else '0'; 
		reg_q2576 <= '1' when reg_fullgraph5 = "000101111" else '0'; 
		reg_q2578 <= '1' when reg_fullgraph5 = "000110000" else '0'; 
		reg_q1042 <= '1' when reg_fullgraph5 = "000110001" else '0'; 
		reg_q1044 <= '1' when reg_fullgraph5 = "000110010" else '0'; 
		reg_q2235 <= '1' when reg_fullgraph5 = "000110011" else '0'; 
		reg_q608 <= '1' when reg_fullgraph5 = "000110100" else '0'; 
		reg_q1658 <= '1' when reg_fullgraph5 = "000110101" else '0'; 
		reg_q1660 <= '1' when reg_fullgraph5 = "000110110" else '0'; 
		reg_q792 <= '1' when reg_fullgraph5 = "000110111" else '0'; 
		reg_q794 <= '1' when reg_fullgraph5 = "000111000" else '0'; 
		reg_q1606 <= '1' when reg_fullgraph5 = "000111001" else '0'; 
		reg_q312 <= '1' when reg_fullgraph5 = "000111010" else '0'; 
		reg_q314 <= '1' when reg_fullgraph5 = "000111011" else '0'; 
		reg_q2479 <= '1' when reg_fullgraph5 = "000111100" else '0'; 
		reg_q1526 <= '1' when reg_fullgraph5 = "000111101" else '0'; 
		reg_q1528 <= '1' when reg_fullgraph5 = "000111110" else '0'; 
		reg_q1844 <= '1' when reg_fullgraph5 = "000111111" else '0'; 
		reg_q890 <= '1' when reg_fullgraph5 = "001000000" else '0'; 
		reg_q892 <= '1' when reg_fullgraph5 = "001000001" else '0'; 
		reg_q183 <= '1' when reg_fullgraph5 = "001000010" else '0'; 
		reg_q2509 <= '1' when reg_fullgraph5 = "001000011" else '0'; 
		reg_q2511 <= '1' when reg_fullgraph5 = "001000100" else '0'; 
		reg_q1858 <= '1' when reg_fullgraph5 = "001000101" else '0'; 
		reg_q1860 <= '1' when reg_fullgraph5 = "001000110" else '0'; 
		reg_q290 <= '1' when reg_fullgraph5 = "001000111" else '0'; 
		reg_q292 <= '1' when reg_fullgraph5 = "001001000" else '0'; 
		reg_q2437 <= '1' when reg_fullgraph5 = "001001001" else '0'; 
		reg_q1473 <= '1' when reg_fullgraph5 = "001001010" else '0'; 
		reg_q1475 <= '1' when reg_fullgraph5 = "001001011" else '0'; 
		reg_q1260 <= '1' when reg_fullgraph5 = "001001100" else '0'; 
		reg_q1262 <= '1' when reg_fullgraph5 = "001001101" else '0'; 
		reg_q575 <= '1' when reg_fullgraph5 = "001001110" else '0'; 
		reg_q1427 <= '1' when reg_fullgraph5 = "001001111" else '0'; 
		reg_q1429 <= '1' when reg_fullgraph5 = "001010000" else '0'; 
		reg_q904 <= '1' when reg_fullgraph5 = "001010001" else '0'; 
		reg_q906 <= '1' when reg_fullgraph5 = "001010010" else '0'; 
		reg_q862 <= '1' when reg_fullgraph5 = "001010011" else '0'; 
		reg_q1832 <= '1' when reg_fullgraph5 = "001010100" else '0'; 
		reg_q1834 <= '1' when reg_fullgraph5 = "001010101" else '0'; 
		reg_q1610 <= '1' when reg_fullgraph5 = "001010110" else '0'; 
		reg_q1612 <= '1' when reg_fullgraph5 = "001010111" else '0'; 
		reg_q767 <= '1' when reg_fullgraph5 = "001011000" else '0'; 
		reg_q1546 <= '1' when reg_fullgraph5 = "001011001" else '0'; 
		reg_q1548 <= '1' when reg_fullgraph5 = "001011010" else '0'; 
		reg_q1854 <= '1' when reg_fullgraph5 = "001011011" else '0'; 
		reg_q1856 <= '1' when reg_fullgraph5 = "001011100" else '0'; 
		reg_q437 <= '1' when reg_fullgraph5 = "001011101" else '0'; 
		reg_q328 <= '1' when reg_fullgraph5 = "001011110" else '0'; 
		reg_q330 <= '1' when reg_fullgraph5 = "001011111" else '0'; 
		reg_q2190 <= '1' when reg_fullgraph5 = "001100000" else '0'; 
		reg_q1600 <= '1' when reg_fullgraph5 = "001100001" else '0'; 
		reg_q2560 <= '1' when reg_fullgraph5 = "001100010" else '0'; 
		reg_q2562 <= '1' when reg_fullgraph5 = "001100011" else '0'; 
		reg_q2168 <= '1' when reg_fullgraph5 = "001100100" else '0'; 
		reg_q2170 <= '1' when reg_fullgraph5 = "001100101" else '0'; 
		reg_q583 <= '1' when reg_fullgraph5 = "001100110" else '0'; 
		reg_q2568 <= '1' when reg_fullgraph5 = "001100111" else '0'; 
		reg_q1431 <= '1' when reg_fullgraph5 = "001101000" else '0'; 
		reg_q419 <= '1' when reg_fullgraph5 = "001101001" else '0'; 
		reg_q415 <= '1' when reg_fullgraph5 = "001101010" else '0'; 
		reg_q417 <= '1' when reg_fullgraph5 = "001101011" else '0'; 
		reg_q1266 <= '1' when reg_fullgraph5 = "001101100" else '0'; 
		reg_q2108 <= '1' when reg_fullgraph5 = "001101101" else '0'; 
		reg_q2110 <= '1' when reg_fullgraph5 = "001101110" else '0'; 
		reg_q1371 <= '1' when reg_fullgraph5 = "001101111" else '0'; 
		reg_q1373 <= '1' when reg_fullgraph5 = "001110000" else '0'; 
		reg_q786 <= '1' when reg_fullgraph5 = "001110001" else '0'; 
		reg_q2659 <= '1' when reg_fullgraph5 = "001110010" else '0'; 
		reg_q2661 <= '1' when reg_fullgraph5 = "001110011" else '0'; 
		reg_q1274 <= '1' when reg_fullgraph5 = "001110100" else '0'; 
		reg_q1276 <= '1' when reg_fullgraph5 = "001110101" else '0'; 
		reg_q2493 <= '1' when reg_fullgraph5 = "001110110" else '0'; 
		reg_q1375 <= '1' when reg_fullgraph5 = "001110111" else '0'; 
		reg_q1405 <= '1' when reg_fullgraph5 = "001111000" else '0'; 
		reg_q1407 <= '1' when reg_fullgraph5 = "001111001" else '0'; 
		reg_q916 <= '1' when reg_fullgraph5 = "001111010" else '0'; 
		reg_q918 <= '1' when reg_fullgraph5 = "001111011" else '0'; 
		reg_q2467 <= '1' when reg_fullgraph5 = "001111100" else '0'; 
		reg_q2469 <= '1' when reg_fullgraph5 = "001111101" else '0'; 
		reg_q1943 <= '1' when reg_fullgraph5 = "001111110" else '0'; 
		reg_q1232 <= '1' when reg_fullgraph5 = "001111111" else '0'; 
		reg_q1234 <= '1' when reg_fullgraph5 = "010000000" else '0'; 
		reg_q1477 <= '1' when reg_fullgraph5 = "010000001" else '0'; 
		reg_q1230 <= '1' when reg_fullgraph5 = "010000010" else '0'; 
		reg_q1250 <= '1' when reg_fullgraph5 = "010000011" else '0'; 
		reg_q1252 <= '1' when reg_fullgraph5 = "010000100" else '0'; 
		reg_q1423 <= '1' when reg_fullgraph5 = "010000101" else '0'; 
		reg_q1425 <= '1' when reg_fullgraph5 = "010000110" else '0'; 
		reg_q2212 <= '1' when reg_fullgraph5 = "010000111" else '0'; 
		reg_q2214 <= '1' when reg_fullgraph5 = "010001000" else '0'; 
		reg_q1288 <= '1' when reg_fullgraph5 = "010001001" else '0'; 
		reg_q1290 <= '1' when reg_fullgraph5 = "010001010" else '0'; 
		reg_q340 <= '1' when reg_fullgraph5 = "010001011" else '0'; 
		reg_q1622 <= '1' when reg_fullgraph5 = "010001100" else '0'; 
		reg_q624 <= '1' when reg_fullgraph5 = "010001101" else '0'; 
		reg_q423 <= '1' when reg_fullgraph5 = "010001110" else '0'; 
		reg_q425 <= '1' when reg_fullgraph5 = "010001111" else '0'; 
		reg_q1588 <= '1' when reg_fullgraph5 = "010010000" else '0'; 
		reg_q1590 <= '1' when reg_fullgraph5 = "010010001" else '0'; 
		reg_q332 <= '1' when reg_fullgraph5 = "010010010" else '0'; 
		reg_q2076 <= '1' when reg_fullgraph5 = "010010011" else '0'; 
		reg_q2078 <= '1' when reg_fullgraph5 = "010010100" else '0'; 
		reg_q1248 <= '1' when reg_fullgraph5 = "010010101" else '0'; 
		reg_q181 <= '1' when reg_fullgraph5 = "010010110" else '0'; 
		reg_q585 <= '1' when reg_fullgraph5 = "010010111" else '0'; 
		reg_q334 <= '1' when reg_fullgraph5 = "010011000" else '0'; 
		reg_q2124 <= '1' when reg_fullgraph5 = "010011001" else '0'; 
		reg_q2126 <= '1' when reg_fullgraph5 = "010011010" else '0'; 
		reg_q2558 <= '1' when reg_fullgraph5 = "010011011" else '0'; 
		reg_q1449 <= '1' when reg_fullgraph5 = "010011100" else '0'; 
		reg_q1451 <= '1' when reg_fullgraph5 = "010011101" else '0'; 
		reg_q835 <= '1' when reg_fullgraph5 = "010011110" else '0'; 
		reg_q837 <= '1' when reg_fullgraph5 = "010011111" else '0'; 
		reg_q626 <= '1' when reg_fullgraph5 = "010100000" else '0'; 
		reg_q628 <= '1' when reg_fullgraph5 = "010100001" else '0'; 
		reg_q1258 <= '1' when reg_fullgraph5 = "010100010" else '0'; 
		reg_q1558 <= '1' when reg_fullgraph5 = "010100011" else '0'; 
		reg_q1668 <= '1' when reg_fullgraph5 = "010100100" else '0'; 
		reg_q1670 <= '1' when reg_fullgraph5 = "010100101" else '0'; 
		reg_q1570 <= '1' when reg_fullgraph5 = "010100110" else '0'; 
		reg_q1572 <= '1' when reg_fullgraph5 = "010100111" else '0'; 
		reg_q1580 <= '1' when reg_fullgraph5 = "010101000" else '0'; 
		reg_q1582 <= '1' when reg_fullgraph5 = "010101001" else '0'; 
		reg_q841 <= '1' when reg_fullgraph5 = "010101010" else '0'; 
		reg_q652 <= '1' when reg_fullgraph5 = "010101011" else '0'; 
		reg_q654 <= '1' when reg_fullgraph5 = "010101100" else '0'; 
		reg_q1409 <= '1' when reg_fullgraph5 = "010101101" else '0'; 
		reg_q839 <= '1' when reg_fullgraph5 = "010101110" else '0'; 
		reg_q1421 <= '1' when reg_fullgraph5 = "010101111" else '0'; 
		reg_q912 <= '1' when reg_fullgraph5 = "010110000" else '0'; 
		reg_q1272 <= '1' when reg_fullgraph5 = "010110001" else '0'; 
		reg_q1614 <= '1' when reg_fullgraph5 = "010110010" else '0'; 
		reg_q2530 <= '1' when reg_fullgraph5 = "010110011" else '0'; 
		reg_q2532 <= '1' when reg_fullgraph5 = "010110100" else '0'; 
		reg_q928 <= '1' when reg_fullgraph5 = "010110101" else '0'; 
		reg_q930 <= '1' when reg_fullgraph5 = "010110110" else '0'; 
		reg_q2198 <= '1' when reg_fullgraph5 = "010110111" else '0'; 
		reg_q2200 <= '1' when reg_fullgraph5 = "010111000" else '0'; 
		reg_q503 <= '1' when reg_fullgraph5 = "010111001" else '0'; 
		reg_q2146 <= '1' when reg_fullgraph5 = "010111010" else '0'; 
		reg_q2148 <= '1' when reg_fullgraph5 = "010111011" else '0'; 
		reg_q926 <= '1' when reg_fullgraph5 = "010111100" else '0'; 
		reg_q1325 <= '1' when reg_fullgraph5 = "010111101" else '0'; 
		reg_q549 <= '1' when reg_fullgraph5 = "010111110" else '0'; 
		reg_q403 <= '1' when reg_fullgraph5 = "010111111" else '0'; 
		reg_q2188 <= '1' when reg_fullgraph5 = "011000000" else '0'; 
		reg_q898 <= '1' when reg_fullgraph5 = "011000001" else '0'; 
		reg_q900 <= '1' when reg_fullgraph5 = "011000010" else '0'; 
		reg_q630 <= '1' when reg_fullgraph5 = "011000011" else '0'; 
		reg_q632 <= '1' when reg_fullgraph5 = "011000100" else '0'; 
		reg_q1455 <= '1' when reg_fullgraph5 = "011000101" else '0'; 
		reg_q1254 <= '1' when reg_fullgraph5 = "011000110" else '0'; 
		reg_q1256 <= '1' when reg_fullgraph5 = "011000111" else '0'; 
		reg_q1138 <= '1' when reg_fullgraph5 = "011001000" else '0'; 
		reg_q1278 <= '1' when reg_fullgraph5 = "011001001" else '0'; 
		reg_q1280 <= '1' when reg_fullgraph5 = "011001010" else '0'; 
		reg_q656 <= '1' when reg_fullgraph5 = "011001011" else '0'; 
		reg_q2540 <= '1' when reg_fullgraph5 = "011001100" else '0'; 
		reg_q2542 <= '1' when reg_fullgraph5 = "011001101" else '0'; 
		reg_q910 <= '1' when reg_fullgraph5 = "011001110" else '0'; 
		reg_q2176 <= '1' when reg_fullgraph5 = "011001111" else '0'; 
		reg_q2178 <= '1' when reg_fullgraph5 = "011010000" else '0'; 
		reg_q2070 <= '1' when reg_fullgraph5 = "011010001" else '0'; 
		reg_q2072 <= '1' when reg_fullgraph5 = "011010010" else '0'; 
		reg_q1242 <= '1' when reg_fullgraph5 = "011010011" else '0'; 
		reg_q1244 <= '1' when reg_fullgraph5 = "011010100" else '0'; 
		reg_q2156 <= '1' when reg_fullgraph5 = "011010101" else '0'; 
		reg_q2158 <= '1' when reg_fullgraph5 = "011010110" else '0'; 
		reg_q2465 <= '1' when reg_fullgraph5 = "011010111" else '0'; 
		reg_q924 <= '1' when reg_fullgraph5 = "011011000" else '0'; 
		reg_q2088 <= '1' when reg_fullgraph5 = "011011001" else '0'; 
		reg_q2090 <= '1' when reg_fullgraph5 = "011011010" else '0'; 
		reg_q2066 <= '1' when reg_fullgraph5 = "011011011" else '0'; 
		reg_q870 <= '1' when reg_fullgraph5 = "011011100" else '0'; 
		reg_q2184 <= '1' when reg_fullgraph5 = "011011101" else '0'; 
		reg_q2186 <= '1' when reg_fullgraph5 = "011011110" else '0'; 
		reg_q864 <= '1' when reg_fullgraph5 = "011011111" else '0'; 
		reg_q866 <= '1' when reg_fullgraph5 = "011100000" else '0'; 
		reg_q2497 <= '1' when reg_fullgraph5 = "011100001" else '0'; 
		reg_q433 <= '1' when reg_fullgraph5 = "011100010" else '0'; 
		reg_q1822 <= '1' when reg_fullgraph5 = "011100011" else '0'; 
		reg_q1662 <= '1' when reg_fullgraph5 = "011100100" else '0'; 
		reg_q2120 <= '1' when reg_fullgraph5 = "011100101" else '0'; 
		reg_q1236 <= '1' when reg_fullgraph5 = "011100110" else '0'; 
		reg_q1036 <= '1' when reg_fullgraph5 = "011100111" else '0'; 
		reg_q1538 <= '1' when reg_fullgraph5 = "011101000" else '0'; 
		reg_q1540 <= '1' when reg_fullgraph5 = "011101001" else '0'; 
		reg_q1550 <= '1' when reg_fullgraph5 = "011101010" else '0'; 
		reg_q1552 <= '1' when reg_fullgraph5 = "011101011" else '0'; 
		reg_q742 <= '1' when reg_fullgraph5 = "011101100" else '0'; 
		reg_q2671 <= '1' when reg_fullgraph5 = "011101101" else '0'; 
		reg_q1284 <= '1' when reg_fullgraph5 = "011101110" else '0'; 
		reg_q1286 <= '1' when reg_fullgraph5 = "011101111" else '0'; 
		reg_q1850 <= '1' when reg_fullgraph5 = "011110000" else '0'; 
		reg_q1852 <= '1' when reg_fullgraph5 = "011110001" else '0'; 
		reg_q1731 <= '1' when reg_fullgraph5 = "011110010" else '0'; 
		reg_q1733 <= '1' when reg_fullgraph5 = "011110011" else '0'; 
		reg_q612 <= '1' when reg_fullgraph5 = "011110100" else '0'; 
		reg_q614 <= '1' when reg_fullgraph5 = "011110101" else '0'; 
		reg_q825 <= '1' when reg_fullgraph5 = "011110110" else '0'; 
		reg_q2206 <= '1' when reg_fullgraph5 = "011110111" else '0'; 
		reg_q2208 <= '1' when reg_fullgraph5 = "011111000" else '0'; 
		reg_q1648 <= '1' when reg_fullgraph5 = "011111001" else '0'; 
		reg_q1650 <= '1' when reg_fullgraph5 = "011111010" else '0'; 
		reg_q1401 <= '1' when reg_fullgraph5 = "011111011" else '0'; 
		reg_q1888 <= '1' when reg_fullgraph5 = "011111100" else '0'; 
		reg_q2471 <= '1' when reg_fullgraph5 = "011111101" else '0'; 
		reg_q2473 <= '1' when reg_fullgraph5 = "011111110" else '0'; 
		reg_q326 <= '1' when reg_fullgraph5 = "011111111" else '0'; 
		reg_q1471 <= '1' when reg_fullgraph5 = "100000000" else '0'; 
		reg_q1246 <= '1' when reg_fullgraph5 = "100000001" else '0'; 
		reg_q2742 <= '1' when reg_fullgraph5 = "100000010" else '0'; 
		reg_q2421 <= '1' when reg_fullgraph5 = "100000011" else '0'; 
		reg_q2423 <= '1' when reg_fullgraph5 = "100000100" else '0'; 
		reg_q579 <= '1' when reg_fullgraph5 = "100000101" else '0'; 
		reg_q932 <= '1' when reg_fullgraph5 = "100000110" else '0'; 
		reg_q934 <= '1' when reg_fullgraph5 = "100000111" else '0'; 
		reg_q1907 <= '1' when reg_fullgraph5 = "100001000" else '0'; 
		reg_q1367 <= '1' when reg_fullgraph5 = "100001001" else '0'; 
		reg_q2665 <= '1' when reg_fullgraph5 = "100001010" else '0'; 
		reg_q2667 <= '1' when reg_fullgraph5 = "100001011" else '0'; 
		reg_q1638 <= '1' when reg_fullgraph5 = "100001100" else '0'; 
		reg_q1967 <= '1' when reg_fullgraph5 = "100001101" else '0'; 
		reg_q1866 <= '1' when reg_fullgraph5 = "100001110" else '0'; 
		reg_q1868 <= '1' when reg_fullgraph5 = "100001111" else '0'; 
		reg_q1304 <= '1' when reg_fullgraph5 = "100010000" else '0'; 
		reg_q1306 <= '1' when reg_fullgraph5 = "100010001" else '0'; 
		reg_q2513 <= '1' when reg_fullgraph5 = "100010010" else '0'; 
		reg_q1870 <= '1' when reg_fullgraph5 = "100010011" else '0'; 
		reg_q1872 <= '1' when reg_fullgraph5 = "100010100" else '0'; 
		reg_q1969 <= '1' when reg_fullgraph5 = "100010101" else '0'; 
		reg_q1971 <= '1' when reg_fullgraph5 = "100010110" else '0'; 
		reg_q577 <= '1' when reg_fullgraph5 = "100010111" else '0'; 
		reg_q413 <= '1' when reg_fullgraph5 = "100011000" else '0'; 
		reg_q405 <= '1' when reg_fullgraph5 = "100011001" else '0'; 
		reg_q407 <= '1' when reg_fullgraph5 = "100011010" else '0'; 
		reg_q2564 <= '1' when reg_fullgraph5 = "100011011" else '0'; 
		reg_q2740 <= '1' when reg_fullgraph5 = "100011100" else '0'; 
		reg_q2477 <= '1' when reg_fullgraph5 = "100011101" else '0'; 
		reg_q1632 <= '1' when reg_fullgraph5 = "100011110" else '0'; 
		reg_q306 <= '1' when reg_fullgraph5 = "100011111" else '0'; 
		reg_q2174 <= '1' when reg_fullgraph5 = "100100000" else '0'; 
		reg_q1282 <= '1' when reg_fullgraph5 = "100100001" else '0'; 
		reg_q2084 <= '1' when reg_fullgraph5 = "100100010" else '0'; 
		reg_q1955 <= '1' when reg_fullgraph5 = "100100011" else '0'; 
		reg_q1957 <= '1' when reg_fullgraph5 = "100100100" else '0'; 
		reg_q1238 <= '1' when reg_fullgraph5 = "100100101" else '0'; 
		reg_q922 <= '1' when reg_fullgraph5 = "100100110" else '0'; 
		reg_q2457 <= '1' when reg_fullgraph5 = "100100111" else '0'; 
		reg_q2459 <= '1' when reg_fullgraph5 = "100101000" else '0'; 
		reg_q463 <= '1' when reg_fullgraph5 = "100101001" else '0'; 
		reg_q465 <= '1' when reg_fullgraph5 = "100101010" else '0'; 
		reg_q320 <= '1' when reg_fullgraph5 = "100101011" else '0'; 
		reg_q322 <= '1' when reg_fullgraph5 = "100101100" else '0'; 
		reg_q2475 <= '1' when reg_fullgraph5 = "100101101" else '0'; 
		reg_q1901 <= '1' when reg_fullgraph5 = "100101110" else '0'; 
		reg_q457 <= '1' when reg_fullgraph5 = "100101111" else '0'; 
		reg_q459 <= '1' when reg_fullgraph5 = "100110000" else '0'; 
		reg_q1560 <= '1' when reg_fullgraph5 = "100110001" else '0'; 
		reg_q1562 <= '1' when reg_fullgraph5 = "100110010" else '0'; 
		reg_q336 <= '1' when reg_fullgraph5 = "100110011" else '0'; 
		reg_q338 <= '1' when reg_fullgraph5 = "100110100" else '0'; 
		reg_q300 <= '1' when reg_fullgraph5 = "100110101" else '0'; 
		reg_q573 <= '1' when reg_fullgraph5 = "100110110" else '0'; 
		reg_q765 <= '1' when reg_fullgraph5 = "100110111" else '0'; 
		reg_q1264 <= '1' when reg_fullgraph5 = "100111000" else '0'; 
		reg_q610 <= '1' when reg_fullgraph5 = "100111001" else '0'; 
		reg_q1512 <= '1' when reg_fullgraph5 = "100111010" else '0'; 
		reg_q453 <= '1' when reg_fullgraph5 = "100111011" else '0'; 
		reg_q2491 <= '1' when reg_fullgraph5 = "100111100" else '0'; 
		reg_q1536 <= '1' when reg_fullgraph5 = "100111101" else '0'; 
		reg_q2202 <= '1' when reg_fullgraph5 = "100111110" else '0'; 
		reg_q2204 <= '1' when reg_fullgraph5 = "100111111" else '0'; 
		reg_q2663 <= '1' when reg_fullgraph5 = "101000000" else '0'; 
		reg_q2566 <= '1' when reg_fullgraph5 = "101000001" else '0'; 
		reg_q2580 <= '1' when reg_fullgraph5 = "101000010" else '0'; 
		reg_q1959 <= '1' when reg_fullgraph5 = "101000011" else '0'; 
		reg_q920 <= '1' when reg_fullgraph5 = "101000100" else '0'; 
		reg_q1654 <= '1' when reg_fullgraph5 = "101000101" else '0'; 
		reg_q1656 <= '1' when reg_fullgraph5 = "101000110" else '0'; 
		reg_q1224 <= '1' when reg_fullgraph5 = "101000111" else '0'; 
		reg_q2106 <= '1' when reg_fullgraph5 = "101001000" else '0'; 
		reg_q2182 <= '1' when reg_fullgraph5 = "101001001" else '0'; 
		reg_q1864 <= '1' when reg_fullgraph5 = "101001010" else '0'; 
		reg_q1586 <= '1' when reg_fullgraph5 = "101001011" else '0'; 
		reg_q2455 <= '1' when reg_fullgraph5 = "101001100" else '0'; 
		reg_q914 <= '1' when reg_fullgraph5 = "101001101" else '0'; 
		reg_q451 <= '1' when reg_fullgraph5 = "101001110" else '0'; 
		reg_q1556 <= '1' when reg_fullgraph5 = "101001111" else '0'; 
		reg_q2132 <= '1' when reg_fullgraph5 = "101010000" else '0'; 
		reg_q2134 <= '1' when reg_fullgraph5 = "101010001" else '0'; 
		reg_q1417 <= '1' when reg_fullgraph5 = "101010010" else '0'; 
		reg_q1419 <= '1' when reg_fullgraph5 = "101010011" else '0'; 
		reg_q872 <= '1' when reg_fullgraph5 = "101010100" else '0'; 
		reg_q638 <= '1' when reg_fullgraph5 = "101010101" else '0'; 
		reg_q640 <= '1' when reg_fullgraph5 = "101010110" else '0'; 
		reg_q431 <= '1' when reg_fullgraph5 = "101010111" else '0'; 
		reg_q1646 <= '1' when reg_fullgraph5 = "101011000" else '0'; 
		reg_q1532 <= '1' when reg_fullgraph5 = "101011001" else '0'; 
		reg_q1624 <= '1' when reg_fullgraph5 = "101011010" else '0'; 
		reg_q1292 <= '1' when reg_fullgraph5 = "101011011" else '0'; 
		reg_q1298 <= '1' when reg_fullgraph5 = "101011100" else '0'; 
		reg_q2196 <= '1' when reg_fullgraph5 = "101011101" else '0'; 
		reg_q936 <= '1' when reg_fullgraph5 = "101011110" else '0'; 
		reg_q938 <= '1' when reg_fullgraph5 = "101011111" else '0'; 
		reg_q1083 <= '1' when reg_fullgraph5 = "101100000" else '0'; 
		reg_q1403 <= '1' when reg_fullgraph5 = "101100001" else '0'; 
		reg_q2140 <= '1' when reg_fullgraph5 = "101100010" else '0'; 
		reg_q2142 <= '1' when reg_fullgraph5 = "101100011" else '0'; 
		reg_q1886 <= '1' when reg_fullgraph5 = "101100100" else '0'; 
		reg_q1828 <= '1' when reg_fullgraph5 = "101100101" else '0'; 
		reg_q1830 <= '1' when reg_fullgraph5 = "101100110" else '0'; 
		reg_q2515 <= '1' when reg_fullgraph5 = "101100111" else '0'; 
		reg_q1381 <= '1' when reg_fullgraph5 = "101101000" else '0'; 
		reg_q1383 <= '1' when reg_fullgraph5 = "101101001" else '0'; 
		reg_q2489 <= '1' when reg_fullgraph5 = "101101010" else '0'; 
		reg_q650 <= '1' when reg_fullgraph5 = "101101011" else '0'; 
		reg_q744 <= '1' when reg_fullgraph5 = "101101100" else '0'; 
		reg_q1953 <= '1' when reg_fullgraph5 = "101101101" else '0'; 
		reg_q581 <= '1' when reg_fullgraph5 = "101101110" else '0'; 
		reg_q1542 <= '1' when reg_fullgraph5 = "101101111" else '0'; 
		reg_q1544 <= '1' when reg_fullgraph5 = "101110000" else '0'; 
		reg_q1842 <= '1' when reg_fullgraph5 = "101110001" else '0'; 
		reg_q2443 <= '1' when reg_fullgraph5 = "101110010" else '0'; 
		reg_q618 <= '1' when reg_fullgraph5 = "101110011" else '0'; 
		reg_q1413 <= '1' when reg_fullgraph5 = "101110100" else '0'; 
		reg_q1415 <= '1' when reg_fullgraph5 = "101110101" else '0'; 
		reg_q2548 <= '1' when reg_fullgraph5 = "101110110" else '0'; 
		reg_q1040 <= '1' when reg_fullgraph5 = "101110111" else '0'; 
		reg_q2096 <= '1' when reg_fullgraph5 = "101111000" else '0'; 
		reg_q2098 <= '1' when reg_fullgraph5 = "101111001" else '0'; 
		reg_q827 <= '1' when reg_fullgraph5 = "101111010" else '0'; 
		reg_q1151 <= '1' when reg_fullgraph5 = "101111011" else '0'; 
		reg_q2144 <= '1' when reg_fullgraph5 = "101111100" else '0'; 
		reg_q888 <= '1' when reg_fullgraph5 = "101111101" else '0'; 
		reg_q616 <= '1' when reg_fullgraph5 = "101111110" else '0'; 
		reg_q1608 <= '1' when reg_fullgraph5 = "101111111" else '0'; 
		reg_q1294 <= '1' when reg_fullgraph5 = "110000000" else '0'; 
		reg_q1240 <= '1' when reg_fullgraph5 = "110000001" else '0'; 
		reg_q658 <= '1' when reg_fullgraph5 = "110000010" else '0'; 
		reg_q886 <= '1' when reg_fullgraph5 = "110000011" else '0'; 
		reg_q1894 <= '1' when reg_fullgraph5 = "110000100" else '0'; 
		reg_q2445 <= '1' when reg_fullgraph5 = "110000101" else '0'; 
		reg_q2138 <= '1' when reg_fullgraph5 = "110000110" else '0'; 
		reg_q2485 <= '1' when reg_fullgraph5 = "110000111" else '0'; 
		reg_q1564 <= '1' when reg_fullgraph5 = "110001000" else '0'; 
		reg_q1566 <= '1' when reg_fullgraph5 = "110001001" else '0'; 
		reg_q1862 <= '1' when reg_fullgraph5 = "110001010" else '0'; 
		reg_q443 <= '1' when reg_fullgraph5 = "110001011" else '0'; 
		reg_q2210 <= '1' when reg_fullgraph5 = "110001100" else '0'; 
		reg_q447 <= '1' when reg_fullgraph5 = "110001101" else '0'; 
		reg_q449 <= '1' when reg_fullgraph5 = "110001110" else '0'; 
		reg_q1840 <= '1' when reg_fullgraph5 = "110001111" else '0'; 
		reg_q1824 <= '1' when reg_fullgraph5 = "110010000" else '0'; 
		reg_q1774 <= '1' when reg_fullgraph5 = "110010001" else '0'; 
		reg_q720 <= '1' when reg_fullgraph5 = "110010010" else '0'; 
		reg_q2483 <= '1' when reg_fullgraph5 = "110010011" else '0'; 
		reg_q2481 <= '1' when reg_fullgraph5 = "110010100" else '0'; 
		reg_q1568 <= '1' when reg_fullgraph5 = "110010101" else '0'; 
		reg_q2128 <= '1' when reg_fullgraph5 = "110010110" else '0'; 
		reg_q1666 <= '1' when reg_fullgraph5 = "110010111" else '0'; 
		reg_q2517 <= '1' when reg_fullgraph5 = "110011000" else '0'; 
		reg_q391 <= '1' when reg_fullgraph5 = "110011001" else '0'; 
		reg_q796 <= '1' when reg_fullgraph5 = "110011010" else '0'; 
		reg_q798 <= '1' when reg_fullgraph5 = "110011011" else '0'; 
		reg_q1878 <= '1' when reg_fullgraph5 = "110011100" else '0'; 
		reg_q1880 <= '1' when reg_fullgraph5 = "110011101" else '0'; 
		reg_q2499 <= '1' when reg_fullgraph5 = "110011110" else '0'; 
		reg_q2086 <= '1' when reg_fullgraph5 = "110011111" else '0'; 
		reg_q2180 <= '1' when reg_fullgraph5 = "110100000" else '0'; 
		reg_q421 <= '1' when reg_fullgraph5 = "110100001" else '0'; 
		reg_q2136 <= '1' when reg_fullgraph5 = "110100010" else '0'; 
		reg_q2507 <= '1' when reg_fullgraph5 = "110100011" else '0'; 
		reg_q2399 <= '1' when reg_fullgraph5 = "110100100" else '0'; 
		reg_q2501 <= '1' when reg_fullgraph5 = "110100101" else '0'; 
		reg_q304 <= '1' when reg_fullgraph5 = "110100110" else '0'; 
		reg_q2100 <= '1' when reg_fullgraph5 = "110100111" else '0'; 
		reg_q1664 <= '1' when reg_fullgraph5 = "110101000" else '0'; 
		reg_q896 <= '1' when reg_fullgraph5 = "110101001" else '0'; 
		reg_q2675 <= '1' when reg_fullgraph5 = "110101010" else '0'; 
		reg_q429 <= '1' when reg_fullgraph5 = "110101011" else '0'; 
		reg_q2657 <= '1' when reg_fullgraph5 = "110101100" else '0'; 
		reg_q2461 <= '1' when reg_fullgraph5 = "110101101" else '0'; 
		reg_q1226 <= '1' when reg_fullgraph5 = "110101110" else '0'; 
		reg_q1228 <= '1' when reg_fullgraph5 = "110101111" else '0'; 
		reg_q642 <= '1' when reg_fullgraph5 = "110110000" else '0'; 
		reg_q302 <= '1' when reg_fullgraph5 = "110110001" else '0'; 
		reg_q1939 <= '1' when reg_fullgraph5 = "110110010" else '0'; 
		reg_q2425 <= '1' when reg_fullgraph5 = "110110011" else '0'; 
		reg_q2427 <= '1' when reg_fullgraph5 = "110110100" else '0'; 
		reg_q1054 <= '1' when reg_fullgraph5 = "110110101" else '0'; 
		reg_q1056 <= '1' when reg_fullgraph5 = "110110110" else '0'; 
		reg_q1826 <= '1' when reg_fullgraph5 = "110110111" else '0'; 
		reg_q1302 <= '1' when reg_fullgraph5 = "110111000" else '0'; 
		reg_q1268 <= '1' when reg_fullgraph5 = "110111001" else '0'; 
		reg_q1874 <= '1' when reg_fullgraph5 = "110111010" else '0'; 
		reg_q2574 <= '1' when reg_fullgraph5 = "110111011" else '0'; 
		reg_q467 <= '1' when reg_fullgraph5 = "110111100" else '0'; 
		reg_q1510 <= '1' when reg_fullgraph5 = "110111101" else '0'; 
		reg_q1199 <= '1' when reg_fullgraph5 = "110111110" else '0'; 
		reg_q1201 <= '1' when reg_fullgraph5 = "110111111" else '0'; 
		reg_q1876 <= '1' when reg_fullgraph5 = "111000000" else '0'; 
		reg_q1435 <= '1' when reg_fullgraph5 = "111000001" else '0'; 
		reg_q1437 <= '1' when reg_fullgraph5 = "111000010" else '0'; 
		reg_q833 <= '1' when reg_fullgraph5 = "111000011" else '0'; 
		reg_q445 <= '1' when reg_fullgraph5 = "111000100" else '0'; 
		reg_q780 <= '1' when reg_fullgraph5 = "111000101" else '0'; 
		reg_q2463 <= '1' when reg_fullgraph5 = "111000110" else '0'; 
		reg_q409 <= '1' when reg_fullgraph5 = "111000111" else '0'; 
		reg_q1920 <= '1' when reg_fullgraph5 = "111001000" else '0'; 
		reg_q829 <= '1' when reg_fullgraph5 = "111001001" else '0'; 
		reg_q831 <= '1' when reg_fullgraph5 = "111001010" else '0'; 
		reg_q1439 <= '1' when reg_fullgraph5 = "111001011" else '0'; 
		reg_q1441 <= '1' when reg_fullgraph5 = "111001100" else '0'; 
		reg_q1678 <= '1' when reg_fullgraph5 = "111001101" else '0'; 
		reg_q1038 <= '1' when reg_fullgraph5 = "111001110" else '0'; 
		reg_q2068 <= '1' when reg_fullgraph5 = "111001111" else '0'; 
		reg_q1048 <= '1' when reg_fullgraph5 = "111010000" else '0'; 
		reg_q1050 <= '1' when reg_fullgraph5 = "111010001" else '0'; 
		reg_q2130 <= '1' when reg_fullgraph5 = "111010010" else '0'; 
		reg_q2166 <= '1' when reg_fullgraph5 = "111010011" else '0'; 
		reg_q324 <= '1' when reg_fullgraph5 = "111010100" else '0'; 
		reg_q1882 <= '1' when reg_fullgraph5 = "111010101" else '0'; 
		reg_q2669 <= '1' when reg_fullgraph5 = "111010110" else '0'; 
		reg_q2102 <= '1' when reg_fullgraph5 = "111010111" else '0'; 
		reg_q908 <= '1' when reg_fullgraph5 = "111011000" else '0'; 
		reg_q1149 <= '1' when reg_fullgraph5 = "111011001" else '0'; 
		reg_q2104 <= '1' when reg_fullgraph5 = "111011010" else '0'; 
		reg_q1838 <= '1' when reg_fullgraph5 = "111011011" else '0'; 
		reg_q1896 <= '1' when reg_fullgraph5 = "111011100" else '0'; 
		reg_q1772 <= '1' when reg_fullgraph5 = "111011101" else '0'; 
		reg_q1433 <= '1' when reg_fullgraph5 = "111011110" else '0'; 
		reg_q1554 <= '1' when reg_fullgraph5 = "111011111" else '0'; 
		reg_q940 <= '1' when reg_fullgraph5 = "111100000" else '0'; 
		reg_q1300 <= '1' when reg_fullgraph5 = "111100001" else '0'; 
		reg_q1836 <= '1' when reg_fullgraph5 = "111100010" else '0'; 
		reg_q2546 <= '1' when reg_fullgraph5 = "111100011" else '0'; 
		reg_q902 <= '1' when reg_fullgraph5 = "111100100" else '0'; 
		reg_q1680 <= '1' when reg_fullgraph5 = "111100101" else '0'; 
		reg_q1030 <= '1' when reg_fullgraph5 = "111100110" else '0'; 
		reg_q1032 <= '1' when reg_fullgraph5 = "111100111" else '0'; 
		reg_q1052 <= '1' when reg_fullgraph5 = "111101000" else '0'; 
		reg_q1898 <= '1' when reg_fullgraph5 = "111101001" else '0'; 
		reg_q1058 <= '1' when reg_fullgraph5 = "111101010" else '0'; 
		reg_q427 <= '1' when reg_fullgraph5 = "111101011" else '0'; 
		reg_q2544 <= '1' when reg_fullgraph5 = "111101100" else '0'; 
--end decoder 

reg_q470_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q470 AND symb_decoder(16#57#)) OR
 					(reg_q470 AND symb_decoder(16#a6#)) OR
 					(reg_q470 AND symb_decoder(16#f7#)) OR
 					(reg_q470 AND symb_decoder(16#31#)) OR
 					(reg_q470 AND symb_decoder(16#e1#)) OR
 					(reg_q470 AND symb_decoder(16#32#)) OR
 					(reg_q470 AND symb_decoder(16#8c#)) OR
 					(reg_q470 AND symb_decoder(16#ee#)) OR
 					(reg_q470 AND symb_decoder(16#ed#)) OR
 					(reg_q470 AND symb_decoder(16#cf#)) OR
 					(reg_q470 AND symb_decoder(16#38#)) OR
 					(reg_q470 AND symb_decoder(16#a8#)) OR
 					(reg_q470 AND symb_decoder(16#86#)) OR
 					(reg_q470 AND symb_decoder(16#6e#)) OR
 					(reg_q470 AND symb_decoder(16#fa#)) OR
 					(reg_q470 AND symb_decoder(16#de#)) OR
 					(reg_q470 AND symb_decoder(16#a1#)) OR
 					(reg_q470 AND symb_decoder(16#00#)) OR
 					(reg_q470 AND symb_decoder(16#d2#)) OR
 					(reg_q470 AND symb_decoder(16#7e#)) OR
 					(reg_q470 AND symb_decoder(16#9b#)) OR
 					(reg_q470 AND symb_decoder(16#42#)) OR
 					(reg_q470 AND symb_decoder(16#cc#)) OR
 					(reg_q470 AND symb_decoder(16#b7#)) OR
 					(reg_q470 AND symb_decoder(16#92#)) OR
 					(reg_q470 AND symb_decoder(16#33#)) OR
 					(reg_q470 AND symb_decoder(16#6c#)) OR
 					(reg_q470 AND symb_decoder(16#f0#)) OR
 					(reg_q470 AND symb_decoder(16#55#)) OR
 					(reg_q470 AND symb_decoder(16#40#)) OR
 					(reg_q470 AND symb_decoder(16#30#)) OR
 					(reg_q470 AND symb_decoder(16#db#)) OR
 					(reg_q470 AND symb_decoder(16#0e#)) OR
 					(reg_q470 AND symb_decoder(16#4a#)) OR
 					(reg_q470 AND symb_decoder(16#a4#)) OR
 					(reg_q470 AND symb_decoder(16#9e#)) OR
 					(reg_q470 AND symb_decoder(16#b0#)) OR
 					(reg_q470 AND symb_decoder(16#63#)) OR
 					(reg_q470 AND symb_decoder(16#94#)) OR
 					(reg_q470 AND symb_decoder(16#ad#)) OR
 					(reg_q470 AND symb_decoder(16#73#)) OR
 					(reg_q470 AND symb_decoder(16#e6#)) OR
 					(reg_q470 AND symb_decoder(16#d3#)) OR
 					(reg_q470 AND symb_decoder(16#46#)) OR
 					(reg_q470 AND symb_decoder(16#f9#)) OR
 					(reg_q470 AND symb_decoder(16#56#)) OR
 					(reg_q470 AND symb_decoder(16#10#)) OR
 					(reg_q470 AND symb_decoder(16#71#)) OR
 					(reg_q470 AND symb_decoder(16#01#)) OR
 					(reg_q470 AND symb_decoder(16#b5#)) OR
 					(reg_q470 AND symb_decoder(16#77#)) OR
 					(reg_q470 AND symb_decoder(16#d4#)) OR
 					(reg_q470 AND symb_decoder(16#8b#)) OR
 					(reg_q470 AND symb_decoder(16#1c#)) OR
 					(reg_q470 AND symb_decoder(16#bf#)) OR
 					(reg_q470 AND symb_decoder(16#ef#)) OR
 					(reg_q470 AND symb_decoder(16#70#)) OR
 					(reg_q470 AND symb_decoder(16#50#)) OR
 					(reg_q470 AND symb_decoder(16#28#)) OR
 					(reg_q470 AND symb_decoder(16#60#)) OR
 					(reg_q470 AND symb_decoder(16#f5#)) OR
 					(reg_q470 AND symb_decoder(16#7c#)) OR
 					(reg_q470 AND symb_decoder(16#98#)) OR
 					(reg_q470 AND symb_decoder(16#09#)) OR
 					(reg_q470 AND symb_decoder(16#1a#)) OR
 					(reg_q470 AND symb_decoder(16#24#)) OR
 					(reg_q470 AND symb_decoder(16#dd#)) OR
 					(reg_q470 AND symb_decoder(16#02#)) OR
 					(reg_q470 AND symb_decoder(16#da#)) OR
 					(reg_q470 AND symb_decoder(16#1e#)) OR
 					(reg_q470 AND symb_decoder(16#15#)) OR
 					(reg_q470 AND symb_decoder(16#ce#)) OR
 					(reg_q470 AND symb_decoder(16#07#)) OR
 					(reg_q470 AND symb_decoder(16#0f#)) OR
 					(reg_q470 AND symb_decoder(16#b2#)) OR
 					(reg_q470 AND symb_decoder(16#b1#)) OR
 					(reg_q470 AND symb_decoder(16#2d#)) OR
 					(reg_q470 AND symb_decoder(16#34#)) OR
 					(reg_q470 AND symb_decoder(16#ea#)) OR
 					(reg_q470 AND symb_decoder(16#4c#)) OR
 					(reg_q470 AND symb_decoder(16#76#)) OR
 					(reg_q470 AND symb_decoder(16#3c#)) OR
 					(reg_q470 AND symb_decoder(16#27#)) OR
 					(reg_q470 AND symb_decoder(16#79#)) OR
 					(reg_q470 AND symb_decoder(16#4e#)) OR
 					(reg_q470 AND symb_decoder(16#b9#)) OR
 					(reg_q470 AND symb_decoder(16#19#)) OR
 					(reg_q470 AND symb_decoder(16#67#)) OR
 					(reg_q470 AND symb_decoder(16#d1#)) OR
 					(reg_q470 AND symb_decoder(16#5d#)) OR
 					(reg_q470 AND symb_decoder(16#c5#)) OR
 					(reg_q470 AND symb_decoder(16#4b#)) OR
 					(reg_q470 AND symb_decoder(16#2c#)) OR
 					(reg_q470 AND symb_decoder(16#ab#)) OR
 					(reg_q470 AND symb_decoder(16#43#)) OR
 					(reg_q470 AND symb_decoder(16#72#)) OR
 					(reg_q470 AND symb_decoder(16#8d#)) OR
 					(reg_q470 AND symb_decoder(16#06#)) OR
 					(reg_q470 AND symb_decoder(16#9f#)) OR
 					(reg_q470 AND symb_decoder(16#9c#)) OR
 					(reg_q470 AND symb_decoder(16#4d#)) OR
 					(reg_q470 AND symb_decoder(16#7a#)) OR
 					(reg_q470 AND symb_decoder(16#9a#)) OR
 					(reg_q470 AND symb_decoder(16#e4#)) OR
 					(reg_q470 AND symb_decoder(16#ca#)) OR
 					(reg_q470 AND symb_decoder(16#99#)) OR
 					(reg_q470 AND symb_decoder(16#74#)) OR
 					(reg_q470 AND symb_decoder(16#e9#)) OR
 					(reg_q470 AND symb_decoder(16#d8#)) OR
 					(reg_q470 AND symb_decoder(16#b3#)) OR
 					(reg_q470 AND symb_decoder(16#d7#)) OR
 					(reg_q470 AND symb_decoder(16#39#)) OR
 					(reg_q470 AND symb_decoder(16#a2#)) OR
 					(reg_q470 AND symb_decoder(16#05#)) OR
 					(reg_q470 AND symb_decoder(16#a5#)) OR
 					(reg_q470 AND symb_decoder(16#81#)) OR
 					(reg_q470 AND symb_decoder(16#bd#)) OR
 					(reg_q470 AND symb_decoder(16#c4#)) OR
 					(reg_q470 AND symb_decoder(16#0d#)) OR
 					(reg_q470 AND symb_decoder(16#58#)) OR
 					(reg_q470 AND symb_decoder(16#5c#)) OR
 					(reg_q470 AND symb_decoder(16#84#)) OR
 					(reg_q470 AND symb_decoder(16#c9#)) OR
 					(reg_q470 AND symb_decoder(16#8e#)) OR
 					(reg_q470 AND symb_decoder(16#c7#)) OR
 					(reg_q470 AND symb_decoder(16#be#)) OR
 					(reg_q470 AND symb_decoder(16#aa#)) OR
 					(reg_q470 AND symb_decoder(16#ae#)) OR
 					(reg_q470 AND symb_decoder(16#65#)) OR
 					(reg_q470 AND symb_decoder(16#f4#)) OR
 					(reg_q470 AND symb_decoder(16#6a#)) OR
 					(reg_q470 AND symb_decoder(16#3e#)) OR
 					(reg_q470 AND symb_decoder(16#47#)) OR
 					(reg_q470 AND symb_decoder(16#3f#)) OR
 					(reg_q470 AND symb_decoder(16#17#)) OR
 					(reg_q470 AND symb_decoder(16#f6#)) OR
 					(reg_q470 AND symb_decoder(16#25#)) OR
 					(reg_q470 AND symb_decoder(16#16#)) OR
 					(reg_q470 AND symb_decoder(16#54#)) OR
 					(reg_q470 AND symb_decoder(16#fe#)) OR
 					(reg_q470 AND symb_decoder(16#c6#)) OR
 					(reg_q470 AND symb_decoder(16#b6#)) OR
 					(reg_q470 AND symb_decoder(16#37#)) OR
 					(reg_q470 AND symb_decoder(16#d6#)) OR
 					(reg_q470 AND symb_decoder(16#0a#)) OR
 					(reg_q470 AND symb_decoder(16#7b#)) OR
 					(reg_q470 AND symb_decoder(16#e2#)) OR
 					(reg_q470 AND symb_decoder(16#0c#)) OR
 					(reg_q470 AND symb_decoder(16#36#)) OR
 					(reg_q470 AND symb_decoder(16#f3#)) OR
 					(reg_q470 AND symb_decoder(16#c3#)) OR
 					(reg_q470 AND symb_decoder(16#ba#)) OR
 					(reg_q470 AND symb_decoder(16#a7#)) OR
 					(reg_q470 AND symb_decoder(16#fc#)) OR
 					(reg_q470 AND symb_decoder(16#fb#)) OR
 					(reg_q470 AND symb_decoder(16#87#)) OR
 					(reg_q470 AND symb_decoder(16#13#)) OR
 					(reg_q470 AND symb_decoder(16#a3#)) OR
 					(reg_q470 AND symb_decoder(16#88#)) OR
 					(reg_q470 AND symb_decoder(16#2e#)) OR
 					(reg_q470 AND symb_decoder(16#22#)) OR
 					(reg_q470 AND symb_decoder(16#6d#)) OR
 					(reg_q470 AND symb_decoder(16#cb#)) OR
 					(reg_q470 AND symb_decoder(16#b8#)) OR
 					(reg_q470 AND symb_decoder(16#8f#)) OR
 					(reg_q470 AND symb_decoder(16#20#)) OR
 					(reg_q470 AND symb_decoder(16#96#)) OR
 					(reg_q470 AND symb_decoder(16#fd#)) OR
 					(reg_q470 AND symb_decoder(16#f1#)) OR
 					(reg_q470 AND symb_decoder(16#c0#)) OR
 					(reg_q470 AND symb_decoder(16#7f#)) OR
 					(reg_q470 AND symb_decoder(16#68#)) OR
 					(reg_q470 AND symb_decoder(16#11#)) OR
 					(reg_q470 AND symb_decoder(16#75#)) OR
 					(reg_q470 AND symb_decoder(16#97#)) OR
 					(reg_q470 AND symb_decoder(16#c1#)) OR
 					(reg_q470 AND symb_decoder(16#85#)) OR
 					(reg_q470 AND symb_decoder(16#bc#)) OR
 					(reg_q470 AND symb_decoder(16#59#)) OR
 					(reg_q470 AND symb_decoder(16#2b#)) OR
 					(reg_q470 AND symb_decoder(16#61#)) OR
 					(reg_q470 AND symb_decoder(16#23#)) OR
 					(reg_q470 AND symb_decoder(16#53#)) OR
 					(reg_q470 AND symb_decoder(16#29#)) OR
 					(reg_q470 AND symb_decoder(16#48#)) OR
 					(reg_q470 AND symb_decoder(16#26#)) OR
 					(reg_q470 AND symb_decoder(16#cd#)) OR
 					(reg_q470 AND symb_decoder(16#df#)) OR
 					(reg_q470 AND symb_decoder(16#64#)) OR
 					(reg_q470 AND symb_decoder(16#21#)) OR
 					(reg_q470 AND symb_decoder(16#1b#)) OR
 					(reg_q470 AND symb_decoder(16#3b#)) OR
 					(reg_q470 AND symb_decoder(16#5e#)) OR
 					(reg_q470 AND symb_decoder(16#80#)) OR
 					(reg_q470 AND symb_decoder(16#66#)) OR
 					(reg_q470 AND symb_decoder(16#b4#)) OR
 					(reg_q470 AND symb_decoder(16#51#)) OR
 					(reg_q470 AND symb_decoder(16#9d#)) OR
 					(reg_q470 AND symb_decoder(16#dc#)) OR
 					(reg_q470 AND symb_decoder(16#ec#)) OR
 					(reg_q470 AND symb_decoder(16#eb#)) OR
 					(reg_q470 AND symb_decoder(16#2a#)) OR
 					(reg_q470 AND symb_decoder(16#45#)) OR
 					(reg_q470 AND symb_decoder(16#90#)) OR
 					(reg_q470 AND symb_decoder(16#4f#)) OR
 					(reg_q470 AND symb_decoder(16#49#)) OR
 					(reg_q470 AND symb_decoder(16#7d#)) OR
 					(reg_q470 AND symb_decoder(16#d9#)) OR
 					(reg_q470 AND symb_decoder(16#44#)) OR
 					(reg_q470 AND symb_decoder(16#14#)) OR
 					(reg_q470 AND symb_decoder(16#41#)) OR
 					(reg_q470 AND symb_decoder(16#a9#)) OR
 					(reg_q470 AND symb_decoder(16#6b#)) OR
 					(reg_q470 AND symb_decoder(16#89#)) OR
 					(reg_q470 AND symb_decoder(16#04#)) OR
 					(reg_q470 AND symb_decoder(16#e3#)) OR
 					(reg_q470 AND symb_decoder(16#18#)) OR
 					(reg_q470 AND symb_decoder(16#e5#)) OR
 					(reg_q470 AND symb_decoder(16#e8#)) OR
 					(reg_q470 AND symb_decoder(16#3d#)) OR
 					(reg_q470 AND symb_decoder(16#69#)) OR
 					(reg_q470 AND symb_decoder(16#1f#)) OR
 					(reg_q470 AND symb_decoder(16#52#)) OR
 					(reg_q470 AND symb_decoder(16#0b#)) OR
 					(reg_q470 AND symb_decoder(16#91#)) OR
 					(reg_q470 AND symb_decoder(16#5f#)) OR
 					(reg_q470 AND symb_decoder(16#f2#)) OR
 					(reg_q470 AND symb_decoder(16#5a#)) OR
 					(reg_q470 AND symb_decoder(16#5b#)) OR
 					(reg_q470 AND symb_decoder(16#82#)) OR
 					(reg_q470 AND symb_decoder(16#8a#)) OR
 					(reg_q470 AND symb_decoder(16#a0#)) OR
 					(reg_q470 AND symb_decoder(16#2f#)) OR
 					(reg_q470 AND symb_decoder(16#3a#)) OR
 					(reg_q470 AND symb_decoder(16#35#)) OR
 					(reg_q470 AND symb_decoder(16#1d#)) OR
 					(reg_q470 AND symb_decoder(16#62#)) OR
 					(reg_q470 AND symb_decoder(16#95#)) OR
 					(reg_q470 AND symb_decoder(16#e7#)) OR
 					(reg_q470 AND symb_decoder(16#ac#)) OR
 					(reg_q470 AND symb_decoder(16#08#)) OR
 					(reg_q470 AND symb_decoder(16#e0#)) OR
 					(reg_q470 AND symb_decoder(16#d0#)) OR
 					(reg_q470 AND symb_decoder(16#12#)) OR
 					(reg_q470 AND symb_decoder(16#bb#)) OR
 					(reg_q470 AND symb_decoder(16#ff#)) OR
 					(reg_q470 AND symb_decoder(16#78#)) OR
 					(reg_q470 AND symb_decoder(16#d5#)) OR
 					(reg_q470 AND symb_decoder(16#93#)) OR
 					(reg_q470 AND symb_decoder(16#03#)) OR
 					(reg_q470 AND symb_decoder(16#83#)) OR
 					(reg_q470 AND symb_decoder(16#c8#)) OR
 					(reg_q470 AND symb_decoder(16#c2#)) OR
 					(reg_q470 AND symb_decoder(16#6f#)) OR
 					(reg_q470 AND symb_decoder(16#f8#)) OR
 					(reg_q470 AND symb_decoder(16#af#));
reg_q470_init <= '0' ;
	p_reg_q470: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q470 <= reg_q470_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q470 <= reg_q470_init;
        else
          reg_q470 <= reg_q470_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q694_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q694 AND symb_decoder(16#4e#)) OR
 					(reg_q694 AND symb_decoder(16#ab#)) OR
 					(reg_q694 AND symb_decoder(16#38#)) OR
 					(reg_q694 AND symb_decoder(16#d9#)) OR
 					(reg_q694 AND symb_decoder(16#35#)) OR
 					(reg_q694 AND symb_decoder(16#e1#)) OR
 					(reg_q694 AND symb_decoder(16#62#)) OR
 					(reg_q694 AND symb_decoder(16#a0#)) OR
 					(reg_q694 AND symb_decoder(16#29#)) OR
 					(reg_q694 AND symb_decoder(16#f0#)) OR
 					(reg_q694 AND symb_decoder(16#3d#)) OR
 					(reg_q694 AND symb_decoder(16#da#)) OR
 					(reg_q694 AND symb_decoder(16#c3#)) OR
 					(reg_q694 AND symb_decoder(16#7f#)) OR
 					(reg_q694 AND symb_decoder(16#8f#)) OR
 					(reg_q694 AND symb_decoder(16#de#)) OR
 					(reg_q694 AND symb_decoder(16#84#)) OR
 					(reg_q694 AND symb_decoder(16#70#)) OR
 					(reg_q694 AND symb_decoder(16#15#)) OR
 					(reg_q694 AND symb_decoder(16#b1#)) OR
 					(reg_q694 AND symb_decoder(16#9c#)) OR
 					(reg_q694 AND symb_decoder(16#6c#)) OR
 					(reg_q694 AND symb_decoder(16#42#)) OR
 					(reg_q694 AND symb_decoder(16#73#)) OR
 					(reg_q694 AND symb_decoder(16#b7#)) OR
 					(reg_q694 AND symb_decoder(16#d6#)) OR
 					(reg_q694 AND symb_decoder(16#4c#)) OR
 					(reg_q694 AND symb_decoder(16#fa#)) OR
 					(reg_q694 AND symb_decoder(16#07#)) OR
 					(reg_q694 AND symb_decoder(16#19#)) OR
 					(reg_q694 AND symb_decoder(16#2a#)) OR
 					(reg_q694 AND symb_decoder(16#01#)) OR
 					(reg_q694 AND symb_decoder(16#cf#)) OR
 					(reg_q694 AND symb_decoder(16#2c#)) OR
 					(reg_q694 AND symb_decoder(16#fe#)) OR
 					(reg_q694 AND symb_decoder(16#09#)) OR
 					(reg_q694 AND symb_decoder(16#80#)) OR
 					(reg_q694 AND symb_decoder(16#b3#)) OR
 					(reg_q694 AND symb_decoder(16#ce#)) OR
 					(reg_q694 AND symb_decoder(16#81#)) OR
 					(reg_q694 AND symb_decoder(16#a6#)) OR
 					(reg_q694 AND symb_decoder(16#4a#)) OR
 					(reg_q694 AND symb_decoder(16#4f#)) OR
 					(reg_q694 AND symb_decoder(16#ef#)) OR
 					(reg_q694 AND symb_decoder(16#1b#)) OR
 					(reg_q694 AND symb_decoder(16#ba#)) OR
 					(reg_q694 AND symb_decoder(16#79#)) OR
 					(reg_q694 AND symb_decoder(16#a4#)) OR
 					(reg_q694 AND symb_decoder(16#21#)) OR
 					(reg_q694 AND symb_decoder(16#30#)) OR
 					(reg_q694 AND symb_decoder(16#94#)) OR
 					(reg_q694 AND symb_decoder(16#e3#)) OR
 					(reg_q694 AND symb_decoder(16#b6#)) OR
 					(reg_q694 AND symb_decoder(16#ea#)) OR
 					(reg_q694 AND symb_decoder(16#91#)) OR
 					(reg_q694 AND symb_decoder(16#ec#)) OR
 					(reg_q694 AND symb_decoder(16#7d#)) OR
 					(reg_q694 AND symb_decoder(16#23#)) OR
 					(reg_q694 AND symb_decoder(16#1a#)) OR
 					(reg_q694 AND symb_decoder(16#e7#)) OR
 					(reg_q694 AND symb_decoder(16#1d#)) OR
 					(reg_q694 AND symb_decoder(16#3a#)) OR
 					(reg_q694 AND symb_decoder(16#66#)) OR
 					(reg_q694 AND symb_decoder(16#68#)) OR
 					(reg_q694 AND symb_decoder(16#39#)) OR
 					(reg_q694 AND symb_decoder(16#d0#)) OR
 					(reg_q694 AND symb_decoder(16#b4#)) OR
 					(reg_q694 AND symb_decoder(16#dd#)) OR
 					(reg_q694 AND symb_decoder(16#1c#)) OR
 					(reg_q694 AND symb_decoder(16#99#)) OR
 					(reg_q694 AND symb_decoder(16#1e#)) OR
 					(reg_q694 AND symb_decoder(16#6a#)) OR
 					(reg_q694 AND symb_decoder(16#fd#)) OR
 					(reg_q694 AND symb_decoder(16#69#)) OR
 					(reg_q694 AND symb_decoder(16#ae#)) OR
 					(reg_q694 AND symb_decoder(16#aa#)) OR
 					(reg_q694 AND symb_decoder(16#40#)) OR
 					(reg_q694 AND symb_decoder(16#b8#)) OR
 					(reg_q694 AND symb_decoder(16#89#)) OR
 					(reg_q694 AND symb_decoder(16#c6#)) OR
 					(reg_q694 AND symb_decoder(16#3f#)) OR
 					(reg_q694 AND symb_decoder(16#86#)) OR
 					(reg_q694 AND symb_decoder(16#bb#)) OR
 					(reg_q694 AND symb_decoder(16#6b#)) OR
 					(reg_q694 AND symb_decoder(16#e9#)) OR
 					(reg_q694 AND symb_decoder(16#67#)) OR
 					(reg_q694 AND symb_decoder(16#a2#)) OR
 					(reg_q694 AND symb_decoder(16#0b#)) OR
 					(reg_q694 AND symb_decoder(16#c8#)) OR
 					(reg_q694 AND symb_decoder(16#f6#)) OR
 					(reg_q694 AND symb_decoder(16#05#)) OR
 					(reg_q694 AND symb_decoder(16#bf#)) OR
 					(reg_q694 AND symb_decoder(16#f5#)) OR
 					(reg_q694 AND symb_decoder(16#5b#)) OR
 					(reg_q694 AND symb_decoder(16#96#)) OR
 					(reg_q694 AND symb_decoder(16#71#)) OR
 					(reg_q694 AND symb_decoder(16#d3#)) OR
 					(reg_q694 AND symb_decoder(16#46#)) OR
 					(reg_q694 AND symb_decoder(16#7a#)) OR
 					(reg_q694 AND symb_decoder(16#6e#)) OR
 					(reg_q694 AND symb_decoder(16#c0#)) OR
 					(reg_q694 AND symb_decoder(16#55#)) OR
 					(reg_q694 AND symb_decoder(16#5d#)) OR
 					(reg_q694 AND symb_decoder(16#3e#)) OR
 					(reg_q694 AND symb_decoder(16#7c#)) OR
 					(reg_q694 AND symb_decoder(16#e5#)) OR
 					(reg_q694 AND symb_decoder(16#48#)) OR
 					(reg_q694 AND symb_decoder(16#8d#)) OR
 					(reg_q694 AND symb_decoder(16#88#)) OR
 					(reg_q694 AND symb_decoder(16#9b#)) OR
 					(reg_q694 AND symb_decoder(16#db#)) OR
 					(reg_q694 AND symb_decoder(16#0a#)) OR
 					(reg_q694 AND symb_decoder(16#18#)) OR
 					(reg_q694 AND symb_decoder(16#52#)) OR
 					(reg_q694 AND symb_decoder(16#16#)) OR
 					(reg_q694 AND symb_decoder(16#14#)) OR
 					(reg_q694 AND symb_decoder(16#a9#)) OR
 					(reg_q694 AND symb_decoder(16#8a#)) OR
 					(reg_q694 AND symb_decoder(16#b2#)) OR
 					(reg_q694 AND symb_decoder(16#44#)) OR
 					(reg_q694 AND symb_decoder(16#58#)) OR
 					(reg_q694 AND symb_decoder(16#32#)) OR
 					(reg_q694 AND symb_decoder(16#0e#)) OR
 					(reg_q694 AND symb_decoder(16#36#)) OR
 					(reg_q694 AND symb_decoder(16#a8#)) OR
 					(reg_q694 AND symb_decoder(16#74#)) OR
 					(reg_q694 AND symb_decoder(16#2b#)) OR
 					(reg_q694 AND symb_decoder(16#72#)) OR
 					(reg_q694 AND symb_decoder(16#f4#)) OR
 					(reg_q694 AND symb_decoder(16#fc#)) OR
 					(reg_q694 AND symb_decoder(16#ac#)) OR
 					(reg_q694 AND symb_decoder(16#e6#)) OR
 					(reg_q694 AND symb_decoder(16#27#)) OR
 					(reg_q694 AND symb_decoder(16#c9#)) OR
 					(reg_q694 AND symb_decoder(16#e0#)) OR
 					(reg_q694 AND symb_decoder(16#ad#)) OR
 					(reg_q694 AND symb_decoder(16#28#)) OR
 					(reg_q694 AND symb_decoder(16#e2#)) OR
 					(reg_q694 AND symb_decoder(16#df#)) OR
 					(reg_q694 AND symb_decoder(16#5a#)) OR
 					(reg_q694 AND symb_decoder(16#f1#)) OR
 					(reg_q694 AND symb_decoder(16#c4#)) OR
 					(reg_q694 AND symb_decoder(16#85#)) OR
 					(reg_q694 AND symb_decoder(16#cc#)) OR
 					(reg_q694 AND symb_decoder(16#3b#)) OR
 					(reg_q694 AND symb_decoder(16#f2#)) OR
 					(reg_q694 AND symb_decoder(16#c1#)) OR
 					(reg_q694 AND symb_decoder(16#f9#)) OR
 					(reg_q694 AND symb_decoder(16#b9#)) OR
 					(reg_q694 AND symb_decoder(16#8c#)) OR
 					(reg_q694 AND symb_decoder(16#af#)) OR
 					(reg_q694 AND symb_decoder(16#9d#)) OR
 					(reg_q694 AND symb_decoder(16#78#)) OR
 					(reg_q694 AND symb_decoder(16#17#)) OR
 					(reg_q694 AND symb_decoder(16#2d#)) OR
 					(reg_q694 AND symb_decoder(16#82#)) OR
 					(reg_q694 AND symb_decoder(16#59#)) OR
 					(reg_q694 AND symb_decoder(16#8e#)) OR
 					(reg_q694 AND symb_decoder(16#95#)) OR
 					(reg_q694 AND symb_decoder(16#22#)) OR
 					(reg_q694 AND symb_decoder(16#c5#)) OR
 					(reg_q694 AND symb_decoder(16#9f#)) OR
 					(reg_q694 AND symb_decoder(16#02#)) OR
 					(reg_q694 AND symb_decoder(16#08#)) OR
 					(reg_q694 AND symb_decoder(16#c7#)) OR
 					(reg_q694 AND symb_decoder(16#54#)) OR
 					(reg_q694 AND symb_decoder(16#6f#)) OR
 					(reg_q694 AND symb_decoder(16#90#)) OR
 					(reg_q694 AND symb_decoder(16#d1#)) OR
 					(reg_q694 AND symb_decoder(16#4b#)) OR
 					(reg_q694 AND symb_decoder(16#47#)) OR
 					(reg_q694 AND symb_decoder(16#04#)) OR
 					(reg_q694 AND symb_decoder(16#75#)) OR
 					(reg_q694 AND symb_decoder(16#98#)) OR
 					(reg_q694 AND symb_decoder(16#37#)) OR
 					(reg_q694 AND symb_decoder(16#87#)) OR
 					(reg_q694 AND symb_decoder(16#e8#)) OR
 					(reg_q694 AND symb_decoder(16#9e#)) OR
 					(reg_q694 AND symb_decoder(16#76#)) OR
 					(reg_q694 AND symb_decoder(16#d4#)) OR
 					(reg_q694 AND symb_decoder(16#57#)) OR
 					(reg_q694 AND symb_decoder(16#97#)) OR
 					(reg_q694 AND symb_decoder(16#53#)) OR
 					(reg_q694 AND symb_decoder(16#0d#)) OR
 					(reg_q694 AND symb_decoder(16#f3#)) OR
 					(reg_q694 AND symb_decoder(16#92#)) OR
 					(reg_q694 AND symb_decoder(16#e4#)) OR
 					(reg_q694 AND symb_decoder(16#65#)) OR
 					(reg_q694 AND symb_decoder(16#8b#)) OR
 					(reg_q694 AND symb_decoder(16#c2#)) OR
 					(reg_q694 AND symb_decoder(16#7e#)) OR
 					(reg_q694 AND symb_decoder(16#12#)) OR
 					(reg_q694 AND symb_decoder(16#dc#)) OR
 					(reg_q694 AND symb_decoder(16#6d#)) OR
 					(reg_q694 AND symb_decoder(16#41#)) OR
 					(reg_q694 AND symb_decoder(16#10#)) OR
 					(reg_q694 AND symb_decoder(16#cd#)) OR
 					(reg_q694 AND symb_decoder(16#56#)) OR
 					(reg_q694 AND symb_decoder(16#d5#)) OR
 					(reg_q694 AND symb_decoder(16#d7#)) OR
 					(reg_q694 AND symb_decoder(16#ff#)) OR
 					(reg_q694 AND symb_decoder(16#b5#)) OR
 					(reg_q694 AND symb_decoder(16#64#)) OR
 					(reg_q694 AND symb_decoder(16#b0#)) OR
 					(reg_q694 AND symb_decoder(16#13#)) OR
 					(reg_q694 AND symb_decoder(16#5e#)) OR
 					(reg_q694 AND symb_decoder(16#25#)) OR
 					(reg_q694 AND symb_decoder(16#ca#)) OR
 					(reg_q694 AND symb_decoder(16#ed#)) OR
 					(reg_q694 AND symb_decoder(16#1f#)) OR
 					(reg_q694 AND symb_decoder(16#83#)) OR
 					(reg_q694 AND symb_decoder(16#51#)) OR
 					(reg_q694 AND symb_decoder(16#49#)) OR
 					(reg_q694 AND symb_decoder(16#20#)) OR
 					(reg_q694 AND symb_decoder(16#2f#)) OR
 					(reg_q694 AND symb_decoder(16#31#)) OR
 					(reg_q694 AND symb_decoder(16#a5#)) OR
 					(reg_q694 AND symb_decoder(16#43#)) OR
 					(reg_q694 AND symb_decoder(16#a7#)) OR
 					(reg_q694 AND symb_decoder(16#f8#)) OR
 					(reg_q694 AND symb_decoder(16#26#)) OR
 					(reg_q694 AND symb_decoder(16#be#)) OR
 					(reg_q694 AND symb_decoder(16#45#)) OR
 					(reg_q694 AND symb_decoder(16#bd#)) OR
 					(reg_q694 AND symb_decoder(16#06#)) OR
 					(reg_q694 AND symb_decoder(16#5f#)) OR
 					(reg_q694 AND symb_decoder(16#d2#)) OR
 					(reg_q694 AND symb_decoder(16#7b#)) OR
 					(reg_q694 AND symb_decoder(16#d8#)) OR
 					(reg_q694 AND symb_decoder(16#33#)) OR
 					(reg_q694 AND symb_decoder(16#4d#)) OR
 					(reg_q694 AND symb_decoder(16#9a#)) OR
 					(reg_q694 AND symb_decoder(16#bc#)) OR
 					(reg_q694 AND symb_decoder(16#eb#)) OR
 					(reg_q694 AND symb_decoder(16#34#)) OR
 					(reg_q694 AND symb_decoder(16#50#)) OR
 					(reg_q694 AND symb_decoder(16#11#)) OR
 					(reg_q694 AND symb_decoder(16#0f#)) OR
 					(reg_q694 AND symb_decoder(16#cb#)) OR
 					(reg_q694 AND symb_decoder(16#a3#)) OR
 					(reg_q694 AND symb_decoder(16#03#)) OR
 					(reg_q694 AND symb_decoder(16#00#)) OR
 					(reg_q694 AND symb_decoder(16#fb#)) OR
 					(reg_q694 AND symb_decoder(16#0c#)) OR
 					(reg_q694 AND symb_decoder(16#3c#)) OR
 					(reg_q694 AND symb_decoder(16#63#)) OR
 					(reg_q694 AND symb_decoder(16#5c#)) OR
 					(reg_q694 AND symb_decoder(16#24#)) OR
 					(reg_q694 AND symb_decoder(16#77#)) OR
 					(reg_q694 AND symb_decoder(16#a1#)) OR
 					(reg_q694 AND symb_decoder(16#61#)) OR
 					(reg_q694 AND symb_decoder(16#f7#)) OR
 					(reg_q694 AND symb_decoder(16#60#)) OR
 					(reg_q694 AND symb_decoder(16#93#)) OR
 					(reg_q694 AND symb_decoder(16#ee#)) OR
 					(reg_q694 AND symb_decoder(16#2e#));
reg_q694_init <= '0' ;
	p_reg_q694: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q694 <= reg_q694_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q694 <= reg_q694_init;
        else
          reg_q694 <= reg_q694_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2229_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q2229 AND symb_decoder(16#dd#)) OR
 					(reg_q2229 AND symb_decoder(16#de#)) OR
 					(reg_q2229 AND symb_decoder(16#55#)) OR
 					(reg_q2229 AND symb_decoder(16#d0#)) OR
 					(reg_q2229 AND symb_decoder(16#24#)) OR
 					(reg_q2229 AND symb_decoder(16#5d#)) OR
 					(reg_q2229 AND symb_decoder(16#04#)) OR
 					(reg_q2229 AND symb_decoder(16#45#)) OR
 					(reg_q2229 AND symb_decoder(16#a2#)) OR
 					(reg_q2229 AND symb_decoder(16#20#)) OR
 					(reg_q2229 AND symb_decoder(16#98#)) OR
 					(reg_q2229 AND symb_decoder(16#9b#)) OR
 					(reg_q2229 AND symb_decoder(16#92#)) OR
 					(reg_q2229 AND symb_decoder(16#db#)) OR
 					(reg_q2229 AND symb_decoder(16#cc#)) OR
 					(reg_q2229 AND symb_decoder(16#13#)) OR
 					(reg_q2229 AND symb_decoder(16#f3#)) OR
 					(reg_q2229 AND symb_decoder(16#79#)) OR
 					(reg_q2229 AND symb_decoder(16#9a#)) OR
 					(reg_q2229 AND symb_decoder(16#ca#)) OR
 					(reg_q2229 AND symb_decoder(16#bd#)) OR
 					(reg_q2229 AND symb_decoder(16#46#)) OR
 					(reg_q2229 AND symb_decoder(16#b9#)) OR
 					(reg_q2229 AND symb_decoder(16#87#)) OR
 					(reg_q2229 AND symb_decoder(16#81#)) OR
 					(reg_q2229 AND symb_decoder(16#c8#)) OR
 					(reg_q2229 AND symb_decoder(16#ef#)) OR
 					(reg_q2229 AND symb_decoder(16#cf#)) OR
 					(reg_q2229 AND symb_decoder(16#32#)) OR
 					(reg_q2229 AND symb_decoder(16#4d#)) OR
 					(reg_q2229 AND symb_decoder(16#38#)) OR
 					(reg_q2229 AND symb_decoder(16#6b#)) OR
 					(reg_q2229 AND symb_decoder(16#12#)) OR
 					(reg_q2229 AND symb_decoder(16#a7#)) OR
 					(reg_q2229 AND symb_decoder(16#36#)) OR
 					(reg_q2229 AND symb_decoder(16#7b#)) OR
 					(reg_q2229 AND symb_decoder(16#97#)) OR
 					(reg_q2229 AND symb_decoder(16#71#)) OR
 					(reg_q2229 AND symb_decoder(16#6e#)) OR
 					(reg_q2229 AND symb_decoder(16#52#)) OR
 					(reg_q2229 AND symb_decoder(16#c9#)) OR
 					(reg_q2229 AND symb_decoder(16#0a#)) OR
 					(reg_q2229 AND symb_decoder(16#23#)) OR
 					(reg_q2229 AND symb_decoder(16#90#)) OR
 					(reg_q2229 AND symb_decoder(16#ae#)) OR
 					(reg_q2229 AND symb_decoder(16#f1#)) OR
 					(reg_q2229 AND symb_decoder(16#84#)) OR
 					(reg_q2229 AND symb_decoder(16#d5#)) OR
 					(reg_q2229 AND symb_decoder(16#c7#)) OR
 					(reg_q2229 AND symb_decoder(16#29#)) OR
 					(reg_q2229 AND symb_decoder(16#7f#)) OR
 					(reg_q2229 AND symb_decoder(16#e0#)) OR
 					(reg_q2229 AND symb_decoder(16#c6#)) OR
 					(reg_q2229 AND symb_decoder(16#2f#)) OR
 					(reg_q2229 AND symb_decoder(16#1a#)) OR
 					(reg_q2229 AND symb_decoder(16#48#)) OR
 					(reg_q2229 AND symb_decoder(16#58#)) OR
 					(reg_q2229 AND symb_decoder(16#07#)) OR
 					(reg_q2229 AND symb_decoder(16#91#)) OR
 					(reg_q2229 AND symb_decoder(16#9d#)) OR
 					(reg_q2229 AND symb_decoder(16#67#)) OR
 					(reg_q2229 AND symb_decoder(16#3e#)) OR
 					(reg_q2229 AND symb_decoder(16#33#)) OR
 					(reg_q2229 AND symb_decoder(16#b2#)) OR
 					(reg_q2229 AND symb_decoder(16#50#)) OR
 					(reg_q2229 AND symb_decoder(16#2a#)) OR
 					(reg_q2229 AND symb_decoder(16#fc#)) OR
 					(reg_q2229 AND symb_decoder(16#d4#)) OR
 					(reg_q2229 AND symb_decoder(16#f9#)) OR
 					(reg_q2229 AND symb_decoder(16#be#)) OR
 					(reg_q2229 AND symb_decoder(16#43#)) OR
 					(reg_q2229 AND symb_decoder(16#75#)) OR
 					(reg_q2229 AND symb_decoder(16#ee#)) OR
 					(reg_q2229 AND symb_decoder(16#99#)) OR
 					(reg_q2229 AND symb_decoder(16#63#)) OR
 					(reg_q2229 AND symb_decoder(16#f4#)) OR
 					(reg_q2229 AND symb_decoder(16#0b#)) OR
 					(reg_q2229 AND symb_decoder(16#e7#)) OR
 					(reg_q2229 AND symb_decoder(16#8d#)) OR
 					(reg_q2229 AND symb_decoder(16#ea#)) OR
 					(reg_q2229 AND symb_decoder(16#80#)) OR
 					(reg_q2229 AND symb_decoder(16#c2#)) OR
 					(reg_q2229 AND symb_decoder(16#aa#)) OR
 					(reg_q2229 AND symb_decoder(16#ad#)) OR
 					(reg_q2229 AND symb_decoder(16#d1#)) OR
 					(reg_q2229 AND symb_decoder(16#8e#)) OR
 					(reg_q2229 AND symb_decoder(16#b4#)) OR
 					(reg_q2229 AND symb_decoder(16#61#)) OR
 					(reg_q2229 AND symb_decoder(16#c1#)) OR
 					(reg_q2229 AND symb_decoder(16#a1#)) OR
 					(reg_q2229 AND symb_decoder(16#ab#)) OR
 					(reg_q2229 AND symb_decoder(16#2e#)) OR
 					(reg_q2229 AND symb_decoder(16#89#)) OR
 					(reg_q2229 AND symb_decoder(16#3d#)) OR
 					(reg_q2229 AND symb_decoder(16#05#)) OR
 					(reg_q2229 AND symb_decoder(16#f0#)) OR
 					(reg_q2229 AND symb_decoder(16#4f#)) OR
 					(reg_q2229 AND symb_decoder(16#d7#)) OR
 					(reg_q2229 AND symb_decoder(16#00#)) OR
 					(reg_q2229 AND symb_decoder(16#34#)) OR
 					(reg_q2229 AND symb_decoder(16#4b#)) OR
 					(reg_q2229 AND symb_decoder(16#6a#)) OR
 					(reg_q2229 AND symb_decoder(16#1f#)) OR
 					(reg_q2229 AND symb_decoder(16#42#)) OR
 					(reg_q2229 AND symb_decoder(16#26#)) OR
 					(reg_q2229 AND symb_decoder(16#b5#)) OR
 					(reg_q2229 AND symb_decoder(16#44#)) OR
 					(reg_q2229 AND symb_decoder(16#d3#)) OR
 					(reg_q2229 AND symb_decoder(16#5b#)) OR
 					(reg_q2229 AND symb_decoder(16#d2#)) OR
 					(reg_q2229 AND symb_decoder(16#b7#)) OR
 					(reg_q2229 AND symb_decoder(16#1e#)) OR
 					(reg_q2229 AND symb_decoder(16#14#)) OR
 					(reg_q2229 AND symb_decoder(16#30#)) OR
 					(reg_q2229 AND symb_decoder(16#17#)) OR
 					(reg_q2229 AND symb_decoder(16#1d#)) OR
 					(reg_q2229 AND symb_decoder(16#a4#)) OR
 					(reg_q2229 AND symb_decoder(16#57#)) OR
 					(reg_q2229 AND symb_decoder(16#51#)) OR
 					(reg_q2229 AND symb_decoder(16#8c#)) OR
 					(reg_q2229 AND symb_decoder(16#c3#)) OR
 					(reg_q2229 AND symb_decoder(16#2b#)) OR
 					(reg_q2229 AND symb_decoder(16#4c#)) OR
 					(reg_q2229 AND symb_decoder(16#06#)) OR
 					(reg_q2229 AND symb_decoder(16#76#)) OR
 					(reg_q2229 AND symb_decoder(16#86#)) OR
 					(reg_q2229 AND symb_decoder(16#ce#)) OR
 					(reg_q2229 AND symb_decoder(16#ba#)) OR
 					(reg_q2229 AND symb_decoder(16#d9#)) OR
 					(reg_q2229 AND symb_decoder(16#f5#)) OR
 					(reg_q2229 AND symb_decoder(16#0e#)) OR
 					(reg_q2229 AND symb_decoder(16#f8#)) OR
 					(reg_q2229 AND symb_decoder(16#8b#)) OR
 					(reg_q2229 AND symb_decoder(16#95#)) OR
 					(reg_q2229 AND symb_decoder(16#a0#)) OR
 					(reg_q2229 AND symb_decoder(16#ac#)) OR
 					(reg_q2229 AND symb_decoder(16#6c#)) OR
 					(reg_q2229 AND symb_decoder(16#e4#)) OR
 					(reg_q2229 AND symb_decoder(16#70#)) OR
 					(reg_q2229 AND symb_decoder(16#a5#)) OR
 					(reg_q2229 AND symb_decoder(16#0f#)) OR
 					(reg_q2229 AND symb_decoder(16#72#)) OR
 					(reg_q2229 AND symb_decoder(16#e9#)) OR
 					(reg_q2229 AND symb_decoder(16#7c#)) OR
 					(reg_q2229 AND symb_decoder(16#d8#)) OR
 					(reg_q2229 AND symb_decoder(16#e2#)) OR
 					(reg_q2229 AND symb_decoder(16#31#)) OR
 					(reg_q2229 AND symb_decoder(16#03#)) OR
 					(reg_q2229 AND symb_decoder(16#b8#)) OR
 					(reg_q2229 AND symb_decoder(16#c5#)) OR
 					(reg_q2229 AND symb_decoder(16#3a#)) OR
 					(reg_q2229 AND symb_decoder(16#df#)) OR
 					(reg_q2229 AND symb_decoder(16#22#)) OR
 					(reg_q2229 AND symb_decoder(16#1c#)) OR
 					(reg_q2229 AND symb_decoder(16#25#)) OR
 					(reg_q2229 AND symb_decoder(16#cd#)) OR
 					(reg_q2229 AND symb_decoder(16#bc#)) OR
 					(reg_q2229 AND symb_decoder(16#fd#)) OR
 					(reg_q2229 AND symb_decoder(16#16#)) OR
 					(reg_q2229 AND symb_decoder(16#3b#)) OR
 					(reg_q2229 AND symb_decoder(16#35#)) OR
 					(reg_q2229 AND symb_decoder(16#64#)) OR
 					(reg_q2229 AND symb_decoder(16#65#)) OR
 					(reg_q2229 AND symb_decoder(16#c0#)) OR
 					(reg_q2229 AND symb_decoder(16#2d#)) OR
 					(reg_q2229 AND symb_decoder(16#8a#)) OR
 					(reg_q2229 AND symb_decoder(16#5c#)) OR
 					(reg_q2229 AND symb_decoder(16#77#)) OR
 					(reg_q2229 AND symb_decoder(16#3f#)) OR
 					(reg_q2229 AND symb_decoder(16#60#)) OR
 					(reg_q2229 AND symb_decoder(16#fe#)) OR
 					(reg_q2229 AND symb_decoder(16#47#)) OR
 					(reg_q2229 AND symb_decoder(16#62#)) OR
 					(reg_q2229 AND symb_decoder(16#f2#)) OR
 					(reg_q2229 AND symb_decoder(16#bb#)) OR
 					(reg_q2229 AND symb_decoder(16#e3#)) OR
 					(reg_q2229 AND symb_decoder(16#09#)) OR
 					(reg_q2229 AND symb_decoder(16#cb#)) OR
 					(reg_q2229 AND symb_decoder(16#96#)) OR
 					(reg_q2229 AND symb_decoder(16#dc#)) OR
 					(reg_q2229 AND symb_decoder(16#6f#)) OR
 					(reg_q2229 AND symb_decoder(16#b1#)) OR
 					(reg_q2229 AND symb_decoder(16#68#)) OR
 					(reg_q2229 AND symb_decoder(16#a6#)) OR
 					(reg_q2229 AND symb_decoder(16#9c#)) OR
 					(reg_q2229 AND symb_decoder(16#fa#)) OR
 					(reg_q2229 AND symb_decoder(16#78#)) OR
 					(reg_q2229 AND symb_decoder(16#5a#)) OR
 					(reg_q2229 AND symb_decoder(16#fb#)) OR
 					(reg_q2229 AND symb_decoder(16#08#)) OR
 					(reg_q2229 AND symb_decoder(16#d6#)) OR
 					(reg_q2229 AND symb_decoder(16#4e#)) OR
 					(reg_q2229 AND symb_decoder(16#37#)) OR
 					(reg_q2229 AND symb_decoder(16#a9#)) OR
 					(reg_q2229 AND symb_decoder(16#59#)) OR
 					(reg_q2229 AND symb_decoder(16#a3#)) OR
 					(reg_q2229 AND symb_decoder(16#e1#)) OR
 					(reg_q2229 AND symb_decoder(16#02#)) OR
 					(reg_q2229 AND symb_decoder(16#7d#)) OR
 					(reg_q2229 AND symb_decoder(16#88#)) OR
 					(reg_q2229 AND symb_decoder(16#b3#)) OR
 					(reg_q2229 AND symb_decoder(16#3c#)) OR
 					(reg_q2229 AND symb_decoder(16#41#)) OR
 					(reg_q2229 AND symb_decoder(16#ec#)) OR
 					(reg_q2229 AND symb_decoder(16#85#)) OR
 					(reg_q2229 AND symb_decoder(16#11#)) OR
 					(reg_q2229 AND symb_decoder(16#2c#)) OR
 					(reg_q2229 AND symb_decoder(16#a8#)) OR
 					(reg_q2229 AND symb_decoder(16#af#)) OR
 					(reg_q2229 AND symb_decoder(16#b6#)) OR
 					(reg_q2229 AND symb_decoder(16#5f#)) OR
 					(reg_q2229 AND symb_decoder(16#9f#)) OR
 					(reg_q2229 AND symb_decoder(16#83#)) OR
 					(reg_q2229 AND symb_decoder(16#69#)) OR
 					(reg_q2229 AND symb_decoder(16#ed#)) OR
 					(reg_q2229 AND symb_decoder(16#93#)) OR
 					(reg_q2229 AND symb_decoder(16#74#)) OR
 					(reg_q2229 AND symb_decoder(16#53#)) OR
 					(reg_q2229 AND symb_decoder(16#7a#)) OR
 					(reg_q2229 AND symb_decoder(16#0c#)) OR
 					(reg_q2229 AND symb_decoder(16#7e#)) OR
 					(reg_q2229 AND symb_decoder(16#da#)) OR
 					(reg_q2229 AND symb_decoder(16#56#)) OR
 					(reg_q2229 AND symb_decoder(16#8f#)) OR
 					(reg_q2229 AND symb_decoder(16#01#)) OR
 					(reg_q2229 AND symb_decoder(16#eb#)) OR
 					(reg_q2229 AND symb_decoder(16#54#)) OR
 					(reg_q2229 AND symb_decoder(16#73#)) OR
 					(reg_q2229 AND symb_decoder(16#5e#)) OR
 					(reg_q2229 AND symb_decoder(16#27#)) OR
 					(reg_q2229 AND symb_decoder(16#bf#)) OR
 					(reg_q2229 AND symb_decoder(16#f6#)) OR
 					(reg_q2229 AND symb_decoder(16#10#)) OR
 					(reg_q2229 AND symb_decoder(16#b0#)) OR
 					(reg_q2229 AND symb_decoder(16#1b#)) OR
 					(reg_q2229 AND symb_decoder(16#f7#)) OR
 					(reg_q2229 AND symb_decoder(16#49#)) OR
 					(reg_q2229 AND symb_decoder(16#ff#)) OR
 					(reg_q2229 AND symb_decoder(16#15#)) OR
 					(reg_q2229 AND symb_decoder(16#0d#)) OR
 					(reg_q2229 AND symb_decoder(16#18#)) OR
 					(reg_q2229 AND symb_decoder(16#66#)) OR
 					(reg_q2229 AND symb_decoder(16#19#)) OR
 					(reg_q2229 AND symb_decoder(16#c4#)) OR
 					(reg_q2229 AND symb_decoder(16#28#)) OR
 					(reg_q2229 AND symb_decoder(16#e6#)) OR
 					(reg_q2229 AND symb_decoder(16#e5#)) OR
 					(reg_q2229 AND symb_decoder(16#6d#)) OR
 					(reg_q2229 AND symb_decoder(16#82#)) OR
 					(reg_q2229 AND symb_decoder(16#4a#)) OR
 					(reg_q2229 AND symb_decoder(16#e8#)) OR
 					(reg_q2229 AND symb_decoder(16#40#)) OR
 					(reg_q2229 AND symb_decoder(16#39#)) OR
 					(reg_q2229 AND symb_decoder(16#9e#)) OR
 					(reg_q2229 AND symb_decoder(16#21#)) OR
 					(reg_q2229 AND symb_decoder(16#94#));
reg_q2229_init <= '0' ;
	p_reg_q2229: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2229 <= reg_q2229_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2229 <= reg_q2229_init;
        else
          reg_q2229 <= reg_q2229_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1756_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1756 AND symb_decoder(16#73#)) OR
 					(reg_q1756 AND symb_decoder(16#56#)) OR
 					(reg_q1756 AND symb_decoder(16#a8#)) OR
 					(reg_q1756 AND symb_decoder(16#03#)) OR
 					(reg_q1756 AND symb_decoder(16#28#)) OR
 					(reg_q1756 AND symb_decoder(16#67#)) OR
 					(reg_q1756 AND symb_decoder(16#4c#)) OR
 					(reg_q1756 AND symb_decoder(16#0b#)) OR
 					(reg_q1756 AND symb_decoder(16#91#)) OR
 					(reg_q1756 AND symb_decoder(16#c7#)) OR
 					(reg_q1756 AND symb_decoder(16#ea#)) OR
 					(reg_q1756 AND symb_decoder(16#93#)) OR
 					(reg_q1756 AND symb_decoder(16#0d#)) OR
 					(reg_q1756 AND symb_decoder(16#d2#)) OR
 					(reg_q1756 AND symb_decoder(16#b8#)) OR
 					(reg_q1756 AND symb_decoder(16#79#)) OR
 					(reg_q1756 AND symb_decoder(16#3b#)) OR
 					(reg_q1756 AND symb_decoder(16#14#)) OR
 					(reg_q1756 AND symb_decoder(16#01#)) OR
 					(reg_q1756 AND symb_decoder(16#ee#)) OR
 					(reg_q1756 AND symb_decoder(16#dc#)) OR
 					(reg_q1756 AND symb_decoder(16#be#)) OR
 					(reg_q1756 AND symb_decoder(16#1f#)) OR
 					(reg_q1756 AND symb_decoder(16#f7#)) OR
 					(reg_q1756 AND symb_decoder(16#20#)) OR
 					(reg_q1756 AND symb_decoder(16#0e#)) OR
 					(reg_q1756 AND symb_decoder(16#4d#)) OR
 					(reg_q1756 AND symb_decoder(16#da#)) OR
 					(reg_q1756 AND symb_decoder(16#1b#)) OR
 					(reg_q1756 AND symb_decoder(16#8e#)) OR
 					(reg_q1756 AND symb_decoder(16#45#)) OR
 					(reg_q1756 AND symb_decoder(16#d4#)) OR
 					(reg_q1756 AND symb_decoder(16#21#)) OR
 					(reg_q1756 AND symb_decoder(16#84#)) OR
 					(reg_q1756 AND symb_decoder(16#74#)) OR
 					(reg_q1756 AND symb_decoder(16#d9#)) OR
 					(reg_q1756 AND symb_decoder(16#d5#)) OR
 					(reg_q1756 AND symb_decoder(16#3a#)) OR
 					(reg_q1756 AND symb_decoder(16#f0#)) OR
 					(reg_q1756 AND symb_decoder(16#ba#)) OR
 					(reg_q1756 AND symb_decoder(16#1c#)) OR
 					(reg_q1756 AND symb_decoder(16#c4#)) OR
 					(reg_q1756 AND symb_decoder(16#00#)) OR
 					(reg_q1756 AND symb_decoder(16#49#)) OR
 					(reg_q1756 AND symb_decoder(16#3c#)) OR
 					(reg_q1756 AND symb_decoder(16#c8#)) OR
 					(reg_q1756 AND symb_decoder(16#8a#)) OR
 					(reg_q1756 AND symb_decoder(16#57#)) OR
 					(reg_q1756 AND symb_decoder(16#77#)) OR
 					(reg_q1756 AND symb_decoder(16#9a#)) OR
 					(reg_q1756 AND symb_decoder(16#92#)) OR
 					(reg_q1756 AND symb_decoder(16#9c#)) OR
 					(reg_q1756 AND symb_decoder(16#04#)) OR
 					(reg_q1756 AND symb_decoder(16#e8#)) OR
 					(reg_q1756 AND symb_decoder(16#b9#)) OR
 					(reg_q1756 AND symb_decoder(16#29#)) OR
 					(reg_q1756 AND symb_decoder(16#8b#)) OR
 					(reg_q1756 AND symb_decoder(16#75#)) OR
 					(reg_q1756 AND symb_decoder(16#6a#)) OR
 					(reg_q1756 AND symb_decoder(16#47#)) OR
 					(reg_q1756 AND symb_decoder(16#09#)) OR
 					(reg_q1756 AND symb_decoder(16#a9#)) OR
 					(reg_q1756 AND symb_decoder(16#3f#)) OR
 					(reg_q1756 AND symb_decoder(16#f6#)) OR
 					(reg_q1756 AND symb_decoder(16#a0#)) OR
 					(reg_q1756 AND symb_decoder(16#6b#)) OR
 					(reg_q1756 AND symb_decoder(16#78#)) OR
 					(reg_q1756 AND symb_decoder(16#fb#)) OR
 					(reg_q1756 AND symb_decoder(16#42#)) OR
 					(reg_q1756 AND symb_decoder(16#30#)) OR
 					(reg_q1756 AND symb_decoder(16#d3#)) OR
 					(reg_q1756 AND symb_decoder(16#f3#)) OR
 					(reg_q1756 AND symb_decoder(16#64#)) OR
 					(reg_q1756 AND symb_decoder(16#88#)) OR
 					(reg_q1756 AND symb_decoder(16#2b#)) OR
 					(reg_q1756 AND symb_decoder(16#38#)) OR
 					(reg_q1756 AND symb_decoder(16#dd#)) OR
 					(reg_q1756 AND symb_decoder(16#c5#)) OR
 					(reg_q1756 AND symb_decoder(16#99#)) OR
 					(reg_q1756 AND symb_decoder(16#eb#)) OR
 					(reg_q1756 AND symb_decoder(16#b6#)) OR
 					(reg_q1756 AND symb_decoder(16#05#)) OR
 					(reg_q1756 AND symb_decoder(16#af#)) OR
 					(reg_q1756 AND symb_decoder(16#3e#)) OR
 					(reg_q1756 AND symb_decoder(16#39#)) OR
 					(reg_q1756 AND symb_decoder(16#e6#)) OR
 					(reg_q1756 AND symb_decoder(16#22#)) OR
 					(reg_q1756 AND symb_decoder(16#32#)) OR
 					(reg_q1756 AND symb_decoder(16#15#)) OR
 					(reg_q1756 AND symb_decoder(16#a3#)) OR
 					(reg_q1756 AND symb_decoder(16#c1#)) OR
 					(reg_q1756 AND symb_decoder(16#ca#)) OR
 					(reg_q1756 AND symb_decoder(16#58#)) OR
 					(reg_q1756 AND symb_decoder(16#8f#)) OR
 					(reg_q1756 AND symb_decoder(16#27#)) OR
 					(reg_q1756 AND symb_decoder(16#86#)) OR
 					(reg_q1756 AND symb_decoder(16#36#)) OR
 					(reg_q1756 AND symb_decoder(16#5e#)) OR
 					(reg_q1756 AND symb_decoder(16#95#)) OR
 					(reg_q1756 AND symb_decoder(16#7c#)) OR
 					(reg_q1756 AND symb_decoder(16#23#)) OR
 					(reg_q1756 AND symb_decoder(16#98#)) OR
 					(reg_q1756 AND symb_decoder(16#bc#)) OR
 					(reg_q1756 AND symb_decoder(16#82#)) OR
 					(reg_q1756 AND symb_decoder(16#9d#)) OR
 					(reg_q1756 AND symb_decoder(16#8d#)) OR
 					(reg_q1756 AND symb_decoder(16#37#)) OR
 					(reg_q1756 AND symb_decoder(16#19#)) OR
 					(reg_q1756 AND symb_decoder(16#cb#)) OR
 					(reg_q1756 AND symb_decoder(16#b5#)) OR
 					(reg_q1756 AND symb_decoder(16#71#)) OR
 					(reg_q1756 AND symb_decoder(16#bd#)) OR
 					(reg_q1756 AND symb_decoder(16#44#)) OR
 					(reg_q1756 AND symb_decoder(16#a5#)) OR
 					(reg_q1756 AND symb_decoder(16#5a#)) OR
 					(reg_q1756 AND symb_decoder(16#b3#)) OR
 					(reg_q1756 AND symb_decoder(16#69#)) OR
 					(reg_q1756 AND symb_decoder(16#2c#)) OR
 					(reg_q1756 AND symb_decoder(16#bf#)) OR
 					(reg_q1756 AND symb_decoder(16#b0#)) OR
 					(reg_q1756 AND symb_decoder(16#a2#)) OR
 					(reg_q1756 AND symb_decoder(16#76#)) OR
 					(reg_q1756 AND symb_decoder(16#89#)) OR
 					(reg_q1756 AND symb_decoder(16#f1#)) OR
 					(reg_q1756 AND symb_decoder(16#52#)) OR
 					(reg_q1756 AND symb_decoder(16#5f#)) OR
 					(reg_q1756 AND symb_decoder(16#25#)) OR
 					(reg_q1756 AND symb_decoder(16#24#)) OR
 					(reg_q1756 AND symb_decoder(16#c6#)) OR
 					(reg_q1756 AND symb_decoder(16#ae#)) OR
 					(reg_q1756 AND symb_decoder(16#cd#)) OR
 					(reg_q1756 AND symb_decoder(16#18#)) OR
 					(reg_q1756 AND symb_decoder(16#f8#)) OR
 					(reg_q1756 AND symb_decoder(16#ff#)) OR
 					(reg_q1756 AND symb_decoder(16#4a#)) OR
 					(reg_q1756 AND symb_decoder(16#48#)) OR
 					(reg_q1756 AND symb_decoder(16#9b#)) OR
 					(reg_q1756 AND symb_decoder(16#43#)) OR
 					(reg_q1756 AND symb_decoder(16#70#)) OR
 					(reg_q1756 AND symb_decoder(16#90#)) OR
 					(reg_q1756 AND symb_decoder(16#a6#)) OR
 					(reg_q1756 AND symb_decoder(16#9f#)) OR
 					(reg_q1756 AND symb_decoder(16#54#)) OR
 					(reg_q1756 AND symb_decoder(16#6d#)) OR
 					(reg_q1756 AND symb_decoder(16#7f#)) OR
 					(reg_q1756 AND symb_decoder(16#f5#)) OR
 					(reg_q1756 AND symb_decoder(16#4b#)) OR
 					(reg_q1756 AND symb_decoder(16#5c#)) OR
 					(reg_q1756 AND symb_decoder(16#d6#)) OR
 					(reg_q1756 AND symb_decoder(16#07#)) OR
 					(reg_q1756 AND symb_decoder(16#50#)) OR
 					(reg_q1756 AND symb_decoder(16#ab#)) OR
 					(reg_q1756 AND symb_decoder(16#4f#)) OR
 					(reg_q1756 AND symb_decoder(16#b4#)) OR
 					(reg_q1756 AND symb_decoder(16#7e#)) OR
 					(reg_q1756 AND symb_decoder(16#34#)) OR
 					(reg_q1756 AND symb_decoder(16#fe#)) OR
 					(reg_q1756 AND symb_decoder(16#1d#)) OR
 					(reg_q1756 AND symb_decoder(16#3d#)) OR
 					(reg_q1756 AND symb_decoder(16#8c#)) OR
 					(reg_q1756 AND symb_decoder(16#c0#)) OR
 					(reg_q1756 AND symb_decoder(16#ec#)) OR
 					(reg_q1756 AND symb_decoder(16#5b#)) OR
 					(reg_q1756 AND symb_decoder(16#aa#)) OR
 					(reg_q1756 AND symb_decoder(16#94#)) OR
 					(reg_q1756 AND symb_decoder(16#a4#)) OR
 					(reg_q1756 AND symb_decoder(16#4e#)) OR
 					(reg_q1756 AND symb_decoder(16#55#)) OR
 					(reg_q1756 AND symb_decoder(16#f2#)) OR
 					(reg_q1756 AND symb_decoder(16#83#)) OR
 					(reg_q1756 AND symb_decoder(16#60#)) OR
 					(reg_q1756 AND symb_decoder(16#5d#)) OR
 					(reg_q1756 AND symb_decoder(16#17#)) OR
 					(reg_q1756 AND symb_decoder(16#96#)) OR
 					(reg_q1756 AND symb_decoder(16#9e#)) OR
 					(reg_q1756 AND symb_decoder(16#51#)) OR
 					(reg_q1756 AND symb_decoder(16#c2#)) OR
 					(reg_q1756 AND symb_decoder(16#40#)) OR
 					(reg_q1756 AND symb_decoder(16#fd#)) OR
 					(reg_q1756 AND symb_decoder(16#ef#)) OR
 					(reg_q1756 AND symb_decoder(16#61#)) OR
 					(reg_q1756 AND symb_decoder(16#e2#)) OR
 					(reg_q1756 AND symb_decoder(16#81#)) OR
 					(reg_q1756 AND symb_decoder(16#97#)) OR
 					(reg_q1756 AND symb_decoder(16#7a#)) OR
 					(reg_q1756 AND symb_decoder(16#33#)) OR
 					(reg_q1756 AND symb_decoder(16#12#)) OR
 					(reg_q1756 AND symb_decoder(16#bb#)) OR
 					(reg_q1756 AND symb_decoder(16#ad#)) OR
 					(reg_q1756 AND symb_decoder(16#63#)) OR
 					(reg_q1756 AND symb_decoder(16#7b#)) OR
 					(reg_q1756 AND symb_decoder(16#a1#)) OR
 					(reg_q1756 AND symb_decoder(16#16#)) OR
 					(reg_q1756 AND symb_decoder(16#c9#)) OR
 					(reg_q1756 AND symb_decoder(16#6c#)) OR
 					(reg_q1756 AND symb_decoder(16#fc#)) OR
 					(reg_q1756 AND symb_decoder(16#46#)) OR
 					(reg_q1756 AND symb_decoder(16#e5#)) OR
 					(reg_q1756 AND symb_decoder(16#de#)) OR
 					(reg_q1756 AND symb_decoder(16#1a#)) OR
 					(reg_q1756 AND symb_decoder(16#41#)) OR
 					(reg_q1756 AND symb_decoder(16#0f#)) OR
 					(reg_q1756 AND symb_decoder(16#ce#)) OR
 					(reg_q1756 AND symb_decoder(16#02#)) OR
 					(reg_q1756 AND symb_decoder(16#31#)) OR
 					(reg_q1756 AND symb_decoder(16#1e#)) OR
 					(reg_q1756 AND symb_decoder(16#fa#)) OR
 					(reg_q1756 AND symb_decoder(16#6e#)) OR
 					(reg_q1756 AND symb_decoder(16#e0#)) OR
 					(reg_q1756 AND symb_decoder(16#0a#)) OR
 					(reg_q1756 AND symb_decoder(16#d0#)) OR
 					(reg_q1756 AND symb_decoder(16#b2#)) OR
 					(reg_q1756 AND symb_decoder(16#a7#)) OR
 					(reg_q1756 AND symb_decoder(16#b7#)) OR
 					(reg_q1756 AND symb_decoder(16#11#)) OR
 					(reg_q1756 AND symb_decoder(16#cc#)) OR
 					(reg_q1756 AND symb_decoder(16#85#)) OR
 					(reg_q1756 AND symb_decoder(16#e3#)) OR
 					(reg_q1756 AND symb_decoder(16#80#)) OR
 					(reg_q1756 AND symb_decoder(16#df#)) OR
 					(reg_q1756 AND symb_decoder(16#ed#)) OR
 					(reg_q1756 AND symb_decoder(16#cf#)) OR
 					(reg_q1756 AND symb_decoder(16#f4#)) OR
 					(reg_q1756 AND symb_decoder(16#2a#)) OR
 					(reg_q1756 AND symb_decoder(16#59#)) OR
 					(reg_q1756 AND symb_decoder(16#68#)) OR
 					(reg_q1756 AND symb_decoder(16#e9#)) OR
 					(reg_q1756 AND symb_decoder(16#66#)) OR
 					(reg_q1756 AND symb_decoder(16#d7#)) OR
 					(reg_q1756 AND symb_decoder(16#7d#)) OR
 					(reg_q1756 AND symb_decoder(16#d8#)) OR
 					(reg_q1756 AND symb_decoder(16#e4#)) OR
 					(reg_q1756 AND symb_decoder(16#ac#)) OR
 					(reg_q1756 AND symb_decoder(16#f9#)) OR
 					(reg_q1756 AND symb_decoder(16#2e#)) OR
 					(reg_q1756 AND symb_decoder(16#13#)) OR
 					(reg_q1756 AND symb_decoder(16#c3#)) OR
 					(reg_q1756 AND symb_decoder(16#db#)) OR
 					(reg_q1756 AND symb_decoder(16#10#)) OR
 					(reg_q1756 AND symb_decoder(16#2d#)) OR
 					(reg_q1756 AND symb_decoder(16#e7#)) OR
 					(reg_q1756 AND symb_decoder(16#53#)) OR
 					(reg_q1756 AND symb_decoder(16#62#)) OR
 					(reg_q1756 AND symb_decoder(16#d1#)) OR
 					(reg_q1756 AND symb_decoder(16#08#)) OR
 					(reg_q1756 AND symb_decoder(16#e1#)) OR
 					(reg_q1756 AND symb_decoder(16#72#)) OR
 					(reg_q1756 AND symb_decoder(16#26#)) OR
 					(reg_q1756 AND symb_decoder(16#35#)) OR
 					(reg_q1756 AND symb_decoder(16#65#)) OR
 					(reg_q1756 AND symb_decoder(16#2f#)) OR
 					(reg_q1756 AND symb_decoder(16#87#)) OR
 					(reg_q1756 AND symb_decoder(16#06#)) OR
 					(reg_q1756 AND symb_decoder(16#6f#)) OR
 					(reg_q1756 AND symb_decoder(16#0c#)) OR
 					(reg_q1756 AND symb_decoder(16#b1#));
reg_q1756_init <= '0' ;
	p_reg_q1756: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1756 <= reg_q1756_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1756 <= reg_q1756_init;
        else
          reg_q1756 <= reg_q1756_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q860_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q860 AND symb_decoder(16#30#)) OR
 					(reg_q860 AND symb_decoder(16#42#)) OR
 					(reg_q860 AND symb_decoder(16#8b#)) OR
 					(reg_q860 AND symb_decoder(16#72#)) OR
 					(reg_q860 AND symb_decoder(16#53#)) OR
 					(reg_q860 AND symb_decoder(16#ef#)) OR
 					(reg_q860 AND symb_decoder(16#cf#)) OR
 					(reg_q860 AND symb_decoder(16#3f#)) OR
 					(reg_q860 AND symb_decoder(16#12#)) OR
 					(reg_q860 AND symb_decoder(16#88#)) OR
 					(reg_q860 AND symb_decoder(16#23#)) OR
 					(reg_q860 AND symb_decoder(16#c3#)) OR
 					(reg_q860 AND symb_decoder(16#ed#)) OR
 					(reg_q860 AND symb_decoder(16#ba#)) OR
 					(reg_q860 AND symb_decoder(16#55#)) OR
 					(reg_q860 AND symb_decoder(16#35#)) OR
 					(reg_q860 AND symb_decoder(16#39#)) OR
 					(reg_q860 AND symb_decoder(16#4e#)) OR
 					(reg_q860 AND symb_decoder(16#3a#)) OR
 					(reg_q860 AND symb_decoder(16#1c#)) OR
 					(reg_q860 AND symb_decoder(16#8e#)) OR
 					(reg_q860 AND symb_decoder(16#14#)) OR
 					(reg_q860 AND symb_decoder(16#9c#)) OR
 					(reg_q860 AND symb_decoder(16#b0#)) OR
 					(reg_q860 AND symb_decoder(16#3d#)) OR
 					(reg_q860 AND symb_decoder(16#43#)) OR
 					(reg_q860 AND symb_decoder(16#5a#)) OR
 					(reg_q860 AND symb_decoder(16#cc#)) OR
 					(reg_q860 AND symb_decoder(16#a7#)) OR
 					(reg_q860 AND symb_decoder(16#e6#)) OR
 					(reg_q860 AND symb_decoder(16#b9#)) OR
 					(reg_q860 AND symb_decoder(16#4d#)) OR
 					(reg_q860 AND symb_decoder(16#24#)) OR
 					(reg_q860 AND symb_decoder(16#0b#)) OR
 					(reg_q860 AND symb_decoder(16#97#)) OR
 					(reg_q860 AND symb_decoder(16#de#)) OR
 					(reg_q860 AND symb_decoder(16#11#)) OR
 					(reg_q860 AND symb_decoder(16#78#)) OR
 					(reg_q860 AND symb_decoder(16#46#)) OR
 					(reg_q860 AND symb_decoder(16#ae#)) OR
 					(reg_q860 AND symb_decoder(16#da#)) OR
 					(reg_q860 AND symb_decoder(16#c1#)) OR
 					(reg_q860 AND symb_decoder(16#27#)) OR
 					(reg_q860 AND symb_decoder(16#9a#)) OR
 					(reg_q860 AND symb_decoder(16#64#)) OR
 					(reg_q860 AND symb_decoder(16#f6#)) OR
 					(reg_q860 AND symb_decoder(16#1b#)) OR
 					(reg_q860 AND symb_decoder(16#63#)) OR
 					(reg_q860 AND symb_decoder(16#f3#)) OR
 					(reg_q860 AND symb_decoder(16#03#)) OR
 					(reg_q860 AND symb_decoder(16#58#)) OR
 					(reg_q860 AND symb_decoder(16#93#)) OR
 					(reg_q860 AND symb_decoder(16#82#)) OR
 					(reg_q860 AND symb_decoder(16#b8#)) OR
 					(reg_q860 AND symb_decoder(16#ff#)) OR
 					(reg_q860 AND symb_decoder(16#b1#)) OR
 					(reg_q860 AND symb_decoder(16#49#)) OR
 					(reg_q860 AND symb_decoder(16#4f#)) OR
 					(reg_q860 AND symb_decoder(16#9f#)) OR
 					(reg_q860 AND symb_decoder(16#44#)) OR
 					(reg_q860 AND symb_decoder(16#b2#)) OR
 					(reg_q860 AND symb_decoder(16#aa#)) OR
 					(reg_q860 AND symb_decoder(16#4c#)) OR
 					(reg_q860 AND symb_decoder(16#33#)) OR
 					(reg_q860 AND symb_decoder(16#48#)) OR
 					(reg_q860 AND symb_decoder(16#86#)) OR
 					(reg_q860 AND symb_decoder(16#62#)) OR
 					(reg_q860 AND symb_decoder(16#00#)) OR
 					(reg_q860 AND symb_decoder(16#75#)) OR
 					(reg_q860 AND symb_decoder(16#f0#)) OR
 					(reg_q860 AND symb_decoder(16#a1#)) OR
 					(reg_q860 AND symb_decoder(16#09#)) OR
 					(reg_q860 AND symb_decoder(16#a4#)) OR
 					(reg_q860 AND symb_decoder(16#c2#)) OR
 					(reg_q860 AND symb_decoder(16#22#)) OR
 					(reg_q860 AND symb_decoder(16#66#)) OR
 					(reg_q860 AND symb_decoder(16#e7#)) OR
 					(reg_q860 AND symb_decoder(16#ac#)) OR
 					(reg_q860 AND symb_decoder(16#8c#)) OR
 					(reg_q860 AND symb_decoder(16#c4#)) OR
 					(reg_q860 AND symb_decoder(16#32#)) OR
 					(reg_q860 AND symb_decoder(16#13#)) OR
 					(reg_q860 AND symb_decoder(16#0d#)) OR
 					(reg_q860 AND symb_decoder(16#80#)) OR
 					(reg_q860 AND symb_decoder(16#85#)) OR
 					(reg_q860 AND symb_decoder(16#59#)) OR
 					(reg_q860 AND symb_decoder(16#f7#)) OR
 					(reg_q860 AND symb_decoder(16#ee#)) OR
 					(reg_q860 AND symb_decoder(16#73#)) OR
 					(reg_q860 AND symb_decoder(16#6e#)) OR
 					(reg_q860 AND symb_decoder(16#b3#)) OR
 					(reg_q860 AND symb_decoder(16#08#)) OR
 					(reg_q860 AND symb_decoder(16#d5#)) OR
 					(reg_q860 AND symb_decoder(16#18#)) OR
 					(reg_q860 AND symb_decoder(16#74#)) OR
 					(reg_q860 AND symb_decoder(16#b5#)) OR
 					(reg_q860 AND symb_decoder(16#dd#)) OR
 					(reg_q860 AND symb_decoder(16#a3#)) OR
 					(reg_q860 AND symb_decoder(16#df#)) OR
 					(reg_q860 AND symb_decoder(16#ec#)) OR
 					(reg_q860 AND symb_decoder(16#40#)) OR
 					(reg_q860 AND symb_decoder(16#60#)) OR
 					(reg_q860 AND symb_decoder(16#fa#)) OR
 					(reg_q860 AND symb_decoder(16#e3#)) OR
 					(reg_q860 AND symb_decoder(16#eb#)) OR
 					(reg_q860 AND symb_decoder(16#be#)) OR
 					(reg_q860 AND symb_decoder(16#b6#)) OR
 					(reg_q860 AND symb_decoder(16#2b#)) OR
 					(reg_q860 AND symb_decoder(16#bf#)) OR
 					(reg_q860 AND symb_decoder(16#7c#)) OR
 					(reg_q860 AND symb_decoder(16#06#)) OR
 					(reg_q860 AND symb_decoder(16#5c#)) OR
 					(reg_q860 AND symb_decoder(16#db#)) OR
 					(reg_q860 AND symb_decoder(16#7f#)) OR
 					(reg_q860 AND symb_decoder(16#5f#)) OR
 					(reg_q860 AND symb_decoder(16#6b#)) OR
 					(reg_q860 AND symb_decoder(16#6f#)) OR
 					(reg_q860 AND symb_decoder(16#ab#)) OR
 					(reg_q860 AND symb_decoder(16#7e#)) OR
 					(reg_q860 AND symb_decoder(16#cd#)) OR
 					(reg_q860 AND symb_decoder(16#fc#)) OR
 					(reg_q860 AND symb_decoder(16#9b#)) OR
 					(reg_q860 AND symb_decoder(16#6d#)) OR
 					(reg_q860 AND symb_decoder(16#d2#)) OR
 					(reg_q860 AND symb_decoder(16#8f#)) OR
 					(reg_q860 AND symb_decoder(16#9e#)) OR
 					(reg_q860 AND symb_decoder(16#b4#)) OR
 					(reg_q860 AND symb_decoder(16#a9#)) OR
 					(reg_q860 AND symb_decoder(16#2c#)) OR
 					(reg_q860 AND symb_decoder(16#c0#)) OR
 					(reg_q860 AND symb_decoder(16#20#)) OR
 					(reg_q860 AND symb_decoder(16#47#)) OR
 					(reg_q860 AND symb_decoder(16#28#)) OR
 					(reg_q860 AND symb_decoder(16#f1#)) OR
 					(reg_q860 AND symb_decoder(16#2d#)) OR
 					(reg_q860 AND symb_decoder(16#3c#)) OR
 					(reg_q860 AND symb_decoder(16#99#)) OR
 					(reg_q860 AND symb_decoder(16#61#)) OR
 					(reg_q860 AND symb_decoder(16#c5#)) OR
 					(reg_q860 AND symb_decoder(16#57#)) OR
 					(reg_q860 AND symb_decoder(16#38#)) OR
 					(reg_q860 AND symb_decoder(16#a8#)) OR
 					(reg_q860 AND symb_decoder(16#8a#)) OR
 					(reg_q860 AND symb_decoder(16#31#)) OR
 					(reg_q860 AND symb_decoder(16#87#)) OR
 					(reg_q860 AND symb_decoder(16#15#)) OR
 					(reg_q860 AND symb_decoder(16#25#)) OR
 					(reg_q860 AND symb_decoder(16#34#)) OR
 					(reg_q860 AND symb_decoder(16#54#)) OR
 					(reg_q860 AND symb_decoder(16#ea#)) OR
 					(reg_q860 AND symb_decoder(16#79#)) OR
 					(reg_q860 AND symb_decoder(16#01#)) OR
 					(reg_q860 AND symb_decoder(16#36#)) OR
 					(reg_q860 AND symb_decoder(16#70#)) OR
 					(reg_q860 AND symb_decoder(16#19#)) OR
 					(reg_q860 AND symb_decoder(16#4b#)) OR
 					(reg_q860 AND symb_decoder(16#71#)) OR
 					(reg_q860 AND symb_decoder(16#a0#)) OR
 					(reg_q860 AND symb_decoder(16#c9#)) OR
 					(reg_q860 AND symb_decoder(16#a2#)) OR
 					(reg_q860 AND symb_decoder(16#37#)) OR
 					(reg_q860 AND symb_decoder(16#fe#)) OR
 					(reg_q860 AND symb_decoder(16#98#)) OR
 					(reg_q860 AND symb_decoder(16#fd#)) OR
 					(reg_q860 AND symb_decoder(16#d7#)) OR
 					(reg_q860 AND symb_decoder(16#e8#)) OR
 					(reg_q860 AND symb_decoder(16#cb#)) OR
 					(reg_q860 AND symb_decoder(16#02#)) OR
 					(reg_q860 AND symb_decoder(16#83#)) OR
 					(reg_q860 AND symb_decoder(16#af#)) OR
 					(reg_q860 AND symb_decoder(16#91#)) OR
 					(reg_q860 AND symb_decoder(16#26#)) OR
 					(reg_q860 AND symb_decoder(16#1a#)) OR
 					(reg_q860 AND symb_decoder(16#5b#)) OR
 					(reg_q860 AND symb_decoder(16#e5#)) OR
 					(reg_q860 AND symb_decoder(16#e1#)) OR
 					(reg_q860 AND symb_decoder(16#68#)) OR
 					(reg_q860 AND symb_decoder(16#bb#)) OR
 					(reg_q860 AND symb_decoder(16#5d#)) OR
 					(reg_q860 AND symb_decoder(16#90#)) OR
 					(reg_q860 AND symb_decoder(16#f5#)) OR
 					(reg_q860 AND symb_decoder(16#84#)) OR
 					(reg_q860 AND symb_decoder(16#16#)) OR
 					(reg_q860 AND symb_decoder(16#c7#)) OR
 					(reg_q860 AND symb_decoder(16#45#)) OR
 					(reg_q860 AND symb_decoder(16#f4#)) OR
 					(reg_q860 AND symb_decoder(16#0f#)) OR
 					(reg_q860 AND symb_decoder(16#07#)) OR
 					(reg_q860 AND symb_decoder(16#92#)) OR
 					(reg_q860 AND symb_decoder(16#67#)) OR
 					(reg_q860 AND symb_decoder(16#51#)) OR
 					(reg_q860 AND symb_decoder(16#50#)) OR
 					(reg_q860 AND symb_decoder(16#0a#)) OR
 					(reg_q860 AND symb_decoder(16#9d#)) OR
 					(reg_q860 AND symb_decoder(16#bd#)) OR
 					(reg_q860 AND symb_decoder(16#d1#)) OR
 					(reg_q860 AND symb_decoder(16#4a#)) OR
 					(reg_q860 AND symb_decoder(16#1d#)) OR
 					(reg_q860 AND symb_decoder(16#41#)) OR
 					(reg_q860 AND symb_decoder(16#1e#)) OR
 					(reg_q860 AND symb_decoder(16#69#)) OR
 					(reg_q860 AND symb_decoder(16#21#)) OR
 					(reg_q860 AND symb_decoder(16#7a#)) OR
 					(reg_q860 AND symb_decoder(16#81#)) OR
 					(reg_q860 AND symb_decoder(16#c8#)) OR
 					(reg_q860 AND symb_decoder(16#ca#)) OR
 					(reg_q860 AND symb_decoder(16#d3#)) OR
 					(reg_q860 AND symb_decoder(16#d6#)) OR
 					(reg_q860 AND symb_decoder(16#6a#)) OR
 					(reg_q860 AND symb_decoder(16#8d#)) OR
 					(reg_q860 AND symb_decoder(16#d8#)) OR
 					(reg_q860 AND symb_decoder(16#d4#)) OR
 					(reg_q860 AND symb_decoder(16#5e#)) OR
 					(reg_q860 AND symb_decoder(16#29#)) OR
 					(reg_q860 AND symb_decoder(16#3b#)) OR
 					(reg_q860 AND symb_decoder(16#f2#)) OR
 					(reg_q860 AND symb_decoder(16#2e#)) OR
 					(reg_q860 AND symb_decoder(16#6c#)) OR
 					(reg_q860 AND symb_decoder(16#a5#)) OR
 					(reg_q860 AND symb_decoder(16#0c#)) OR
 					(reg_q860 AND symb_decoder(16#ce#)) OR
 					(reg_q860 AND symb_decoder(16#ad#)) OR
 					(reg_q860 AND symb_decoder(16#a6#)) OR
 					(reg_q860 AND symb_decoder(16#0e#)) OR
 					(reg_q860 AND symb_decoder(16#c6#)) OR
 					(reg_q860 AND symb_decoder(16#65#)) OR
 					(reg_q860 AND symb_decoder(16#52#)) OR
 					(reg_q860 AND symb_decoder(16#17#)) OR
 					(reg_q860 AND symb_decoder(16#e9#)) OR
 					(reg_q860 AND symb_decoder(16#e4#)) OR
 					(reg_q860 AND symb_decoder(16#89#)) OR
 					(reg_q860 AND symb_decoder(16#f9#)) OR
 					(reg_q860 AND symb_decoder(16#04#)) OR
 					(reg_q860 AND symb_decoder(16#e2#)) OR
 					(reg_q860 AND symb_decoder(16#dc#)) OR
 					(reg_q860 AND symb_decoder(16#e0#)) OR
 					(reg_q860 AND symb_decoder(16#fb#)) OR
 					(reg_q860 AND symb_decoder(16#96#)) OR
 					(reg_q860 AND symb_decoder(16#d9#)) OR
 					(reg_q860 AND symb_decoder(16#f8#)) OR
 					(reg_q860 AND symb_decoder(16#7d#)) OR
 					(reg_q860 AND symb_decoder(16#05#)) OR
 					(reg_q860 AND symb_decoder(16#7b#)) OR
 					(reg_q860 AND symb_decoder(16#95#)) OR
 					(reg_q860 AND symb_decoder(16#2a#)) OR
 					(reg_q860 AND symb_decoder(16#76#)) OR
 					(reg_q860 AND symb_decoder(16#bc#)) OR
 					(reg_q860 AND symb_decoder(16#1f#)) OR
 					(reg_q860 AND symb_decoder(16#2f#)) OR
 					(reg_q860 AND symb_decoder(16#d0#)) OR
 					(reg_q860 AND symb_decoder(16#77#)) OR
 					(reg_q860 AND symb_decoder(16#94#)) OR
 					(reg_q860 AND symb_decoder(16#56#)) OR
 					(reg_q860 AND symb_decoder(16#b7#)) OR
 					(reg_q860 AND symb_decoder(16#10#)) OR
 					(reg_q860 AND symb_decoder(16#3e#));
reg_q860_init <= '0' ;
	p_reg_q860: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q860 <= reg_q860_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q860 <= reg_q860_init;
        else
          reg_q860 <= reg_q860_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph11

reg_q1975_in <= (reg_q1961 AND symb_decoder(16#a9#)) OR
 					(reg_q1961 AND symb_decoder(16#4f#)) OR
 					(reg_q1961 AND symb_decoder(16#d7#)) OR
 					(reg_q1961 AND symb_decoder(16#40#)) OR
 					(reg_q1961 AND symb_decoder(16#1a#)) OR
 					(reg_q1961 AND symb_decoder(16#f3#)) OR
 					(reg_q1961 AND symb_decoder(16#8c#)) OR
 					(reg_q1961 AND symb_decoder(16#a5#)) OR
 					(reg_q1961 AND symb_decoder(16#1e#)) OR
 					(reg_q1961 AND symb_decoder(16#b3#)) OR
 					(reg_q1961 AND symb_decoder(16#b5#)) OR
 					(reg_q1961 AND symb_decoder(16#ba#)) OR
 					(reg_q1961 AND symb_decoder(16#fb#)) OR
 					(reg_q1961 AND symb_decoder(16#9f#)) OR
 					(reg_q1961 AND symb_decoder(16#2c#)) OR
 					(reg_q1961 AND symb_decoder(16#0f#)) OR
 					(reg_q1961 AND symb_decoder(16#21#)) OR
 					(reg_q1961 AND symb_decoder(16#62#)) OR
 					(reg_q1961 AND symb_decoder(16#6d#)) OR
 					(reg_q1961 AND symb_decoder(16#e7#)) OR
 					(reg_q1961 AND symb_decoder(16#e6#)) OR
 					(reg_q1961 AND symb_decoder(16#93#)) OR
 					(reg_q1961 AND symb_decoder(16#5b#)) OR
 					(reg_q1961 AND symb_decoder(16#74#)) OR
 					(reg_q1961 AND symb_decoder(16#ce#)) OR
 					(reg_q1961 AND symb_decoder(16#65#)) OR
 					(reg_q1961 AND symb_decoder(16#07#)) OR
 					(reg_q1961 AND symb_decoder(16#d4#)) OR
 					(reg_q1961 AND symb_decoder(16#29#)) OR
 					(reg_q1961 AND symb_decoder(16#70#)) OR
 					(reg_q1961 AND symb_decoder(16#cb#)) OR
 					(reg_q1961 AND symb_decoder(16#44#)) OR
 					(reg_q1961 AND symb_decoder(16#f2#)) OR
 					(reg_q1961 AND symb_decoder(16#4e#)) OR
 					(reg_q1961 AND symb_decoder(16#c2#)) OR
 					(reg_q1961 AND symb_decoder(16#eb#)) OR
 					(reg_q1961 AND symb_decoder(16#8b#)) OR
 					(reg_q1961 AND symb_decoder(16#56#)) OR
 					(reg_q1961 AND symb_decoder(16#6b#)) OR
 					(reg_q1961 AND symb_decoder(16#a8#)) OR
 					(reg_q1961 AND symb_decoder(16#69#)) OR
 					(reg_q1961 AND symb_decoder(16#72#)) OR
 					(reg_q1961 AND symb_decoder(16#2a#)) OR
 					(reg_q1961 AND symb_decoder(16#33#)) OR
 					(reg_q1961 AND symb_decoder(16#5e#)) OR
 					(reg_q1961 AND symb_decoder(16#58#)) OR
 					(reg_q1961 AND symb_decoder(16#32#)) OR
 					(reg_q1961 AND symb_decoder(16#f6#)) OR
 					(reg_q1961 AND symb_decoder(16#48#)) OR
 					(reg_q1961 AND symb_decoder(16#c1#)) OR
 					(reg_q1961 AND symb_decoder(16#66#)) OR
 					(reg_q1961 AND symb_decoder(16#08#)) OR
 					(reg_q1961 AND symb_decoder(16#9a#)) OR
 					(reg_q1961 AND symb_decoder(16#63#)) OR
 					(reg_q1961 AND symb_decoder(16#dd#)) OR
 					(reg_q1961 AND symb_decoder(16#af#)) OR
 					(reg_q1961 AND symb_decoder(16#bd#)) OR
 					(reg_q1961 AND symb_decoder(16#20#)) OR
 					(reg_q1961 AND symb_decoder(16#64#)) OR
 					(reg_q1961 AND symb_decoder(16#79#)) OR
 					(reg_q1961 AND symb_decoder(16#7b#)) OR
 					(reg_q1961 AND symb_decoder(16#d2#)) OR
 					(reg_q1961 AND symb_decoder(16#26#)) OR
 					(reg_q1961 AND symb_decoder(16#c6#)) OR
 					(reg_q1961 AND symb_decoder(16#e5#)) OR
 					(reg_q1961 AND symb_decoder(16#90#)) OR
 					(reg_q1961 AND symb_decoder(16#95#)) OR
 					(reg_q1961 AND symb_decoder(16#6f#)) OR
 					(reg_q1961 AND symb_decoder(16#6e#)) OR
 					(reg_q1961 AND symb_decoder(16#99#)) OR
 					(reg_q1961 AND symb_decoder(16#1c#)) OR
 					(reg_q1961 AND symb_decoder(16#87#)) OR
 					(reg_q1961 AND symb_decoder(16#24#)) OR
 					(reg_q1961 AND symb_decoder(16#cd#)) OR
 					(reg_q1961 AND symb_decoder(16#25#)) OR
 					(reg_q1961 AND symb_decoder(16#6a#)) OR
 					(reg_q1961 AND symb_decoder(16#9b#)) OR
 					(reg_q1961 AND symb_decoder(16#68#)) OR
 					(reg_q1961 AND symb_decoder(16#ad#)) OR
 					(reg_q1961 AND symb_decoder(16#55#)) OR
 					(reg_q1961 AND symb_decoder(16#39#)) OR
 					(reg_q1961 AND symb_decoder(16#cf#)) OR
 					(reg_q1961 AND symb_decoder(16#3f#)) OR
 					(reg_q1961 AND symb_decoder(16#fd#)) OR
 					(reg_q1961 AND symb_decoder(16#27#)) OR
 					(reg_q1961 AND symb_decoder(16#d8#)) OR
 					(reg_q1961 AND symb_decoder(16#5c#)) OR
 					(reg_q1961 AND symb_decoder(16#30#)) OR
 					(reg_q1961 AND symb_decoder(16#aa#)) OR
 					(reg_q1961 AND symb_decoder(16#81#)) OR
 					(reg_q1961 AND symb_decoder(16#df#)) OR
 					(reg_q1961 AND symb_decoder(16#98#)) OR
 					(reg_q1961 AND symb_decoder(16#14#)) OR
 					(reg_q1961 AND symb_decoder(16#06#)) OR
 					(reg_q1961 AND symb_decoder(16#13#)) OR
 					(reg_q1961 AND symb_decoder(16#ef#)) OR
 					(reg_q1961 AND symb_decoder(16#2d#)) OR
 					(reg_q1961 AND symb_decoder(16#57#)) OR
 					(reg_q1961 AND symb_decoder(16#e4#)) OR
 					(reg_q1961 AND symb_decoder(16#73#)) OR
 					(reg_q1961 AND symb_decoder(16#a0#)) OR
 					(reg_q1961 AND symb_decoder(16#75#)) OR
 					(reg_q1961 AND symb_decoder(16#7c#)) OR
 					(reg_q1961 AND symb_decoder(16#67#)) OR
 					(reg_q1961 AND symb_decoder(16#6c#)) OR
 					(reg_q1961 AND symb_decoder(16#91#)) OR
 					(reg_q1961 AND symb_decoder(16#85#)) OR
 					(reg_q1961 AND symb_decoder(16#89#)) OR
 					(reg_q1961 AND symb_decoder(16#50#)) OR
 					(reg_q1961 AND symb_decoder(16#2e#)) OR
 					(reg_q1961 AND symb_decoder(16#ac#)) OR
 					(reg_q1961 AND symb_decoder(16#96#)) OR
 					(reg_q1961 AND symb_decoder(16#ff#)) OR
 					(reg_q1961 AND symb_decoder(16#ee#)) OR
 					(reg_q1961 AND symb_decoder(16#bf#)) OR
 					(reg_q1961 AND symb_decoder(16#23#)) OR
 					(reg_q1961 AND symb_decoder(16#d5#)) OR
 					(reg_q1961 AND symb_decoder(16#e1#)) OR
 					(reg_q1961 AND symb_decoder(16#35#)) OR
 					(reg_q1961 AND symb_decoder(16#d9#)) OR
 					(reg_q1961 AND symb_decoder(16#00#)) OR
 					(reg_q1961 AND symb_decoder(16#47#)) OR
 					(reg_q1961 AND symb_decoder(16#db#)) OR
 					(reg_q1961 AND symb_decoder(16#92#)) OR
 					(reg_q1961 AND symb_decoder(16#03#)) OR
 					(reg_q1961 AND symb_decoder(16#3d#)) OR
 					(reg_q1961 AND symb_decoder(16#60#)) OR
 					(reg_q1961 AND symb_decoder(16#cc#)) OR
 					(reg_q1961 AND symb_decoder(16#d1#)) OR
 					(reg_q1961 AND symb_decoder(16#c8#)) OR
 					(reg_q1961 AND symb_decoder(16#88#)) OR
 					(reg_q1961 AND symb_decoder(16#c9#)) OR
 					(reg_q1961 AND symb_decoder(16#c4#)) OR
 					(reg_q1961 AND symb_decoder(16#a4#)) OR
 					(reg_q1961 AND symb_decoder(16#dc#)) OR
 					(reg_q1961 AND symb_decoder(16#a3#)) OR
 					(reg_q1961 AND symb_decoder(16#46#)) OR
 					(reg_q1961 AND symb_decoder(16#e9#)) OR
 					(reg_q1961 AND symb_decoder(16#a6#)) OR
 					(reg_q1961 AND symb_decoder(16#15#)) OR
 					(reg_q1961 AND symb_decoder(16#12#)) OR
 					(reg_q1961 AND symb_decoder(16#0c#)) OR
 					(reg_q1961 AND symb_decoder(16#bc#)) OR
 					(reg_q1961 AND symb_decoder(16#da#)) OR
 					(reg_q1961 AND symb_decoder(16#fa#)) OR
 					(reg_q1961 AND symb_decoder(16#be#)) OR
 					(reg_q1961 AND symb_decoder(16#f4#)) OR
 					(reg_q1961 AND symb_decoder(16#9c#)) OR
 					(reg_q1961 AND symb_decoder(16#49#)) OR
 					(reg_q1961 AND symb_decoder(16#b0#)) OR
 					(reg_q1961 AND symb_decoder(16#ed#)) OR
 					(reg_q1961 AND symb_decoder(16#86#)) OR
 					(reg_q1961 AND symb_decoder(16#fe#)) OR
 					(reg_q1961 AND symb_decoder(16#31#)) OR
 					(reg_q1961 AND symb_decoder(16#10#)) OR
 					(reg_q1961 AND symb_decoder(16#7e#)) OR
 					(reg_q1961 AND symb_decoder(16#ab#)) OR
 					(reg_q1961 AND symb_decoder(16#7f#)) OR
 					(reg_q1961 AND symb_decoder(16#3b#)) OR
 					(reg_q1961 AND symb_decoder(16#16#)) OR
 					(reg_q1961 AND symb_decoder(16#e0#)) OR
 					(reg_q1961 AND symb_decoder(16#f0#)) OR
 					(reg_q1961 AND symb_decoder(16#1f#)) OR
 					(reg_q1961 AND symb_decoder(16#77#)) OR
 					(reg_q1961 AND symb_decoder(16#ec#)) OR
 					(reg_q1961 AND symb_decoder(16#83#)) OR
 					(reg_q1961 AND symb_decoder(16#0e#)) OR
 					(reg_q1961 AND symb_decoder(16#e2#)) OR
 					(reg_q1961 AND symb_decoder(16#c0#)) OR
 					(reg_q1961 AND symb_decoder(16#8e#)) OR
 					(reg_q1961 AND symb_decoder(16#22#)) OR
 					(reg_q1961 AND symb_decoder(16#5d#)) OR
 					(reg_q1961 AND symb_decoder(16#59#)) OR
 					(reg_q1961 AND symb_decoder(16#5f#)) OR
 					(reg_q1961 AND symb_decoder(16#3a#)) OR
 					(reg_q1961 AND symb_decoder(16#2f#)) OR
 					(reg_q1961 AND symb_decoder(16#11#)) OR
 					(reg_q1961 AND symb_decoder(16#4d#)) OR
 					(reg_q1961 AND symb_decoder(16#b4#)) OR
 					(reg_q1961 AND symb_decoder(16#04#)) OR
 					(reg_q1961 AND symb_decoder(16#43#)) OR
 					(reg_q1961 AND symb_decoder(16#de#)) OR
 					(reg_q1961 AND symb_decoder(16#45#)) OR
 					(reg_q1961 AND symb_decoder(16#9d#)) OR
 					(reg_q1961 AND symb_decoder(16#0b#)) OR
 					(reg_q1961 AND symb_decoder(16#c7#)) OR
 					(reg_q1961 AND symb_decoder(16#8a#)) OR
 					(reg_q1961 AND symb_decoder(16#f5#)) OR
 					(reg_q1961 AND symb_decoder(16#52#)) OR
 					(reg_q1961 AND symb_decoder(16#a1#)) OR
 					(reg_q1961 AND symb_decoder(16#7a#)) OR
 					(reg_q1961 AND symb_decoder(16#bb#)) OR
 					(reg_q1961 AND symb_decoder(16#53#)) OR
 					(reg_q1961 AND symb_decoder(16#97#)) OR
 					(reg_q1961 AND symb_decoder(16#17#)) OR
 					(reg_q1961 AND symb_decoder(16#e8#)) OR
 					(reg_q1961 AND symb_decoder(16#d6#)) OR
 					(reg_q1961 AND symb_decoder(16#8f#)) OR
 					(reg_q1961 AND symb_decoder(16#2b#)) OR
 					(reg_q1961 AND symb_decoder(16#f7#)) OR
 					(reg_q1961 AND symb_decoder(16#b1#)) OR
 					(reg_q1961 AND symb_decoder(16#ea#)) OR
 					(reg_q1961 AND symb_decoder(16#94#)) OR
 					(reg_q1961 AND symb_decoder(16#28#)) OR
 					(reg_q1961 AND symb_decoder(16#1d#)) OR
 					(reg_q1961 AND symb_decoder(16#f9#)) OR
 					(reg_q1961 AND symb_decoder(16#b7#)) OR
 					(reg_q1961 AND symb_decoder(16#8d#)) OR
 					(reg_q1961 AND symb_decoder(16#34#)) OR
 					(reg_q1961 AND symb_decoder(16#4b#)) OR
 					(reg_q1961 AND symb_decoder(16#fc#)) OR
 					(reg_q1961 AND symb_decoder(16#02#)) OR
 					(reg_q1961 AND symb_decoder(16#61#)) OR
 					(reg_q1961 AND symb_decoder(16#d3#)) OR
 					(reg_q1961 AND symb_decoder(16#f8#)) OR
 					(reg_q1961 AND symb_decoder(16#3c#)) OR
 					(reg_q1961 AND symb_decoder(16#5a#)) OR
 					(reg_q1961 AND symb_decoder(16#51#)) OR
 					(reg_q1961 AND symb_decoder(16#b8#)) OR
 					(reg_q1961 AND symb_decoder(16#76#)) OR
 					(reg_q1961 AND symb_decoder(16#84#)) OR
 					(reg_q1961 AND symb_decoder(16#38#)) OR
 					(reg_q1961 AND symb_decoder(16#41#)) OR
 					(reg_q1961 AND symb_decoder(16#18#)) OR
 					(reg_q1961 AND symb_decoder(16#54#)) OR
 					(reg_q1961 AND symb_decoder(16#ca#)) OR
 					(reg_q1961 AND symb_decoder(16#09#)) OR
 					(reg_q1961 AND symb_decoder(16#71#)) OR
 					(reg_q1961 AND symb_decoder(16#36#)) OR
 					(reg_q1961 AND symb_decoder(16#c3#)) OR
 					(reg_q1961 AND symb_decoder(16#9e#)) OR
 					(reg_q1961 AND symb_decoder(16#82#)) OR
 					(reg_q1961 AND symb_decoder(16#4c#)) OR
 					(reg_q1961 AND symb_decoder(16#b9#)) OR
 					(reg_q1961 AND symb_decoder(16#19#)) OR
 					(reg_q1961 AND symb_decoder(16#a7#)) OR
 					(reg_q1961 AND symb_decoder(16#3e#)) OR
 					(reg_q1961 AND symb_decoder(16#f1#)) OR
 					(reg_q1961 AND symb_decoder(16#01#)) OR
 					(reg_q1961 AND symb_decoder(16#a2#)) OR
 					(reg_q1961 AND symb_decoder(16#c5#)) OR
 					(reg_q1961 AND symb_decoder(16#d0#)) OR
 					(reg_q1961 AND symb_decoder(16#1b#)) OR
 					(reg_q1961 AND symb_decoder(16#e3#)) OR
 					(reg_q1961 AND symb_decoder(16#80#)) OR
 					(reg_q1961 AND symb_decoder(16#7d#)) OR
 					(reg_q1961 AND symb_decoder(16#05#)) OR
 					(reg_q1961 AND symb_decoder(16#b6#)) OR
 					(reg_q1961 AND symb_decoder(16#b2#)) OR
 					(reg_q1961 AND symb_decoder(16#ae#)) OR
 					(reg_q1961 AND symb_decoder(16#42#)) OR
 					(reg_q1961 AND symb_decoder(16#37#)) OR
 					(reg_q1961 AND symb_decoder(16#4a#)) OR
 					(reg_q1961 AND symb_decoder(16#78#)) OR
 					(reg_q1975 AND symb_decoder(16#46#)) OR
 					(reg_q1975 AND symb_decoder(16#55#)) OR
 					(reg_q1975 AND symb_decoder(16#db#)) OR
 					(reg_q1975 AND symb_decoder(16#d7#)) OR
 					(reg_q1975 AND symb_decoder(16#66#)) OR
 					(reg_q1975 AND symb_decoder(16#56#)) OR
 					(reg_q1975 AND symb_decoder(16#84#)) OR
 					(reg_q1975 AND symb_decoder(16#27#)) OR
 					(reg_q1975 AND symb_decoder(16#0c#)) OR
 					(reg_q1975 AND symb_decoder(16#04#)) OR
 					(reg_q1975 AND symb_decoder(16#24#)) OR
 					(reg_q1975 AND symb_decoder(16#bd#)) OR
 					(reg_q1975 AND symb_decoder(16#61#)) OR
 					(reg_q1975 AND symb_decoder(16#3a#)) OR
 					(reg_q1975 AND symb_decoder(16#b1#)) OR
 					(reg_q1975 AND symb_decoder(16#bb#)) OR
 					(reg_q1975 AND symb_decoder(16#ad#)) OR
 					(reg_q1975 AND symb_decoder(16#10#)) OR
 					(reg_q1975 AND symb_decoder(16#fc#)) OR
 					(reg_q1975 AND symb_decoder(16#6a#)) OR
 					(reg_q1975 AND symb_decoder(16#2c#)) OR
 					(reg_q1975 AND symb_decoder(16#65#)) OR
 					(reg_q1975 AND symb_decoder(16#4f#)) OR
 					(reg_q1975 AND symb_decoder(16#35#)) OR
 					(reg_q1975 AND symb_decoder(16#f4#)) OR
 					(reg_q1975 AND symb_decoder(16#ac#)) OR
 					(reg_q1975 AND symb_decoder(16#18#)) OR
 					(reg_q1975 AND symb_decoder(16#c7#)) OR
 					(reg_q1975 AND symb_decoder(16#05#)) OR
 					(reg_q1975 AND symb_decoder(16#cd#)) OR
 					(reg_q1975 AND symb_decoder(16#2b#)) OR
 					(reg_q1975 AND symb_decoder(16#4c#)) OR
 					(reg_q1975 AND symb_decoder(16#64#)) OR
 					(reg_q1975 AND symb_decoder(16#f6#)) OR
 					(reg_q1975 AND symb_decoder(16#63#)) OR
 					(reg_q1975 AND symb_decoder(16#02#)) OR
 					(reg_q1975 AND symb_decoder(16#ee#)) OR
 					(reg_q1975 AND symb_decoder(16#c6#)) OR
 					(reg_q1975 AND symb_decoder(16#bc#)) OR
 					(reg_q1975 AND symb_decoder(16#77#)) OR
 					(reg_q1975 AND symb_decoder(16#51#)) OR
 					(reg_q1975 AND symb_decoder(16#07#)) OR
 					(reg_q1975 AND symb_decoder(16#4a#)) OR
 					(reg_q1975 AND symb_decoder(16#33#)) OR
 					(reg_q1975 AND symb_decoder(16#70#)) OR
 					(reg_q1975 AND symb_decoder(16#fb#)) OR
 					(reg_q1975 AND symb_decoder(16#94#)) OR
 					(reg_q1975 AND symb_decoder(16#9f#)) OR
 					(reg_q1975 AND symb_decoder(16#e9#)) OR
 					(reg_q1975 AND symb_decoder(16#c1#)) OR
 					(reg_q1975 AND symb_decoder(16#08#)) OR
 					(reg_q1975 AND symb_decoder(16#3e#)) OR
 					(reg_q1975 AND symb_decoder(16#6d#)) OR
 					(reg_q1975 AND symb_decoder(16#30#)) OR
 					(reg_q1975 AND symb_decoder(16#41#)) OR
 					(reg_q1975 AND symb_decoder(16#d6#)) OR
 					(reg_q1975 AND symb_decoder(16#38#)) OR
 					(reg_q1975 AND symb_decoder(16#c0#)) OR
 					(reg_q1975 AND symb_decoder(16#9b#)) OR
 					(reg_q1975 AND symb_decoder(16#c8#)) OR
 					(reg_q1975 AND symb_decoder(16#39#)) OR
 					(reg_q1975 AND symb_decoder(16#4d#)) OR
 					(reg_q1975 AND symb_decoder(16#03#)) OR
 					(reg_q1975 AND symb_decoder(16#97#)) OR
 					(reg_q1975 AND symb_decoder(16#85#)) OR
 					(reg_q1975 AND symb_decoder(16#0f#)) OR
 					(reg_q1975 AND symb_decoder(16#a7#)) OR
 					(reg_q1975 AND symb_decoder(16#e1#)) OR
 					(reg_q1975 AND symb_decoder(16#c5#)) OR
 					(reg_q1975 AND symb_decoder(16#00#)) OR
 					(reg_q1975 AND symb_decoder(16#be#)) OR
 					(reg_q1975 AND symb_decoder(16#60#)) OR
 					(reg_q1975 AND symb_decoder(16#36#)) OR
 					(reg_q1975 AND symb_decoder(16#23#)) OR
 					(reg_q1975 AND symb_decoder(16#1d#)) OR
 					(reg_q1975 AND symb_decoder(16#3b#)) OR
 					(reg_q1975 AND symb_decoder(16#26#)) OR
 					(reg_q1975 AND symb_decoder(16#25#)) OR
 					(reg_q1975 AND symb_decoder(16#d0#)) OR
 					(reg_q1975 AND symb_decoder(16#de#)) OR
 					(reg_q1975 AND symb_decoder(16#01#)) OR
 					(reg_q1975 AND symb_decoder(16#19#)) OR
 					(reg_q1975 AND symb_decoder(16#e7#)) OR
 					(reg_q1975 AND symb_decoder(16#9e#)) OR
 					(reg_q1975 AND symb_decoder(16#20#)) OR
 					(reg_q1975 AND symb_decoder(16#5b#)) OR
 					(reg_q1975 AND symb_decoder(16#b3#)) OR
 					(reg_q1975 AND symb_decoder(16#b5#)) OR
 					(reg_q1975 AND symb_decoder(16#74#)) OR
 					(reg_q1975 AND symb_decoder(16#d2#)) OR
 					(reg_q1975 AND symb_decoder(16#29#)) OR
 					(reg_q1975 AND symb_decoder(16#48#)) OR
 					(reg_q1975 AND symb_decoder(16#ae#)) OR
 					(reg_q1975 AND symb_decoder(16#eb#)) OR
 					(reg_q1975 AND symb_decoder(16#90#)) OR
 					(reg_q1975 AND symb_decoder(16#9c#)) OR
 					(reg_q1975 AND symb_decoder(16#c4#)) OR
 					(reg_q1975 AND symb_decoder(16#82#)) OR
 					(reg_q1975 AND symb_decoder(16#f1#)) OR
 					(reg_q1975 AND symb_decoder(16#df#)) OR
 					(reg_q1975 AND symb_decoder(16#75#)) OR
 					(reg_q1975 AND symb_decoder(16#b4#)) OR
 					(reg_q1975 AND symb_decoder(16#b9#)) OR
 					(reg_q1975 AND symb_decoder(16#fa#)) OR
 					(reg_q1975 AND symb_decoder(16#59#)) OR
 					(reg_q1975 AND symb_decoder(16#5c#)) OR
 					(reg_q1975 AND symb_decoder(16#d8#)) OR
 					(reg_q1975 AND symb_decoder(16#81#)) OR
 					(reg_q1975 AND symb_decoder(16#93#)) OR
 					(reg_q1975 AND symb_decoder(16#88#)) OR
 					(reg_q1975 AND symb_decoder(16#12#)) OR
 					(reg_q1975 AND symb_decoder(16#ec#)) OR
 					(reg_q1975 AND symb_decoder(16#b0#)) OR
 					(reg_q1975 AND symb_decoder(16#0e#)) OR
 					(reg_q1975 AND symb_decoder(16#a2#)) OR
 					(reg_q1975 AND symb_decoder(16#e5#)) OR
 					(reg_q1975 AND symb_decoder(16#7c#)) OR
 					(reg_q1975 AND symb_decoder(16#68#)) OR
 					(reg_q1975 AND symb_decoder(16#5f#)) OR
 					(reg_q1975 AND symb_decoder(16#45#)) OR
 					(reg_q1975 AND symb_decoder(16#98#)) OR
 					(reg_q1975 AND symb_decoder(16#58#)) OR
 					(reg_q1975 AND symb_decoder(16#72#)) OR
 					(reg_q1975 AND symb_decoder(16#f3#)) OR
 					(reg_q1975 AND symb_decoder(16#1c#)) OR
 					(reg_q1975 AND symb_decoder(16#5d#)) OR
 					(reg_q1975 AND symb_decoder(16#aa#)) OR
 					(reg_q1975 AND symb_decoder(16#cc#)) OR
 					(reg_q1975 AND symb_decoder(16#67#)) OR
 					(reg_q1975 AND symb_decoder(16#e6#)) OR
 					(reg_q1975 AND symb_decoder(16#6b#)) OR
 					(reg_q1975 AND symb_decoder(16#9d#)) OR
 					(reg_q1975 AND symb_decoder(16#89#)) OR
 					(reg_q1975 AND symb_decoder(16#50#)) OR
 					(reg_q1975 AND symb_decoder(16#cf#)) OR
 					(reg_q1975 AND symb_decoder(16#dd#)) OR
 					(reg_q1975 AND symb_decoder(16#2a#)) OR
 					(reg_q1975 AND symb_decoder(16#8f#)) OR
 					(reg_q1975 AND symb_decoder(16#4b#)) OR
 					(reg_q1975 AND symb_decoder(16#f2#)) OR
 					(reg_q1975 AND symb_decoder(16#5a#)) OR
 					(reg_q1975 AND symb_decoder(16#11#)) OR
 					(reg_q1975 AND symb_decoder(16#e4#)) OR
 					(reg_q1975 AND symb_decoder(16#a9#)) OR
 					(reg_q1975 AND symb_decoder(16#d9#)) OR
 					(reg_q1975 AND symb_decoder(16#6c#)) OR
 					(reg_q1975 AND symb_decoder(16#f9#)) OR
 					(reg_q1975 AND symb_decoder(16#37#)) OR
 					(reg_q1975 AND symb_decoder(16#d3#)) OR
 					(reg_q1975 AND symb_decoder(16#87#)) OR
 					(reg_q1975 AND symb_decoder(16#8d#)) OR
 					(reg_q1975 AND symb_decoder(16#da#)) OR
 					(reg_q1975 AND symb_decoder(16#a3#)) OR
 					(reg_q1975 AND symb_decoder(16#5e#)) OR
 					(reg_q1975 AND symb_decoder(16#f0#)) OR
 					(reg_q1975 AND symb_decoder(16#1e#)) OR
 					(reg_q1975 AND symb_decoder(16#43#)) OR
 					(reg_q1975 AND symb_decoder(16#bf#)) OR
 					(reg_q1975 AND symb_decoder(16#80#)) OR
 					(reg_q1975 AND symb_decoder(16#f8#)) OR
 					(reg_q1975 AND symb_decoder(16#fe#)) OR
 					(reg_q1975 AND symb_decoder(16#96#)) OR
 					(reg_q1975 AND symb_decoder(16#44#)) OR
 					(reg_q1975 AND symb_decoder(16#6e#)) OR
 					(reg_q1975 AND symb_decoder(16#1a#)) OR
 					(reg_q1975 AND symb_decoder(16#32#)) OR
 					(reg_q1975 AND symb_decoder(16#b8#)) OR
 					(reg_q1975 AND symb_decoder(16#2e#)) OR
 					(reg_q1975 AND symb_decoder(16#fd#)) OR
 					(reg_q1975 AND symb_decoder(16#ef#)) OR
 					(reg_q1975 AND symb_decoder(16#71#)) OR
 					(reg_q1975 AND symb_decoder(16#6f#)) OR
 					(reg_q1975 AND symb_decoder(16#b7#)) OR
 					(reg_q1975 AND symb_decoder(16#ff#)) OR
 					(reg_q1975 AND symb_decoder(16#1b#)) OR
 					(reg_q1975 AND symb_decoder(16#ed#)) OR
 					(reg_q1975 AND symb_decoder(16#83#)) OR
 					(reg_q1975 AND symb_decoder(16#ca#)) OR
 					(reg_q1975 AND symb_decoder(16#c9#)) OR
 					(reg_q1975 AND symb_decoder(16#69#)) OR
 					(reg_q1975 AND symb_decoder(16#e8#)) OR
 					(reg_q1975 AND symb_decoder(16#f7#)) OR
 					(reg_q1975 AND symb_decoder(16#8a#)) OR
 					(reg_q1975 AND symb_decoder(16#16#)) OR
 					(reg_q1975 AND symb_decoder(16#7f#)) OR
 					(reg_q1975 AND symb_decoder(16#a4#)) OR
 					(reg_q1975 AND symb_decoder(16#c2#)) OR
 					(reg_q1975 AND symb_decoder(16#28#)) OR
 					(reg_q1975 AND symb_decoder(16#a5#)) OR
 					(reg_q1975 AND symb_decoder(16#79#)) OR
 					(reg_q1975 AND symb_decoder(16#d1#)) OR
 					(reg_q1975 AND symb_decoder(16#17#)) OR
 					(reg_q1975 AND symb_decoder(16#73#)) OR
 					(reg_q1975 AND symb_decoder(16#d4#)) OR
 					(reg_q1975 AND symb_decoder(16#49#)) OR
 					(reg_q1975 AND symb_decoder(16#14#)) OR
 					(reg_q1975 AND symb_decoder(16#b2#)) OR
 					(reg_q1975 AND symb_decoder(16#ea#)) OR
 					(reg_q1975 AND symb_decoder(16#ce#)) OR
 					(reg_q1975 AND symb_decoder(16#86#)) OR
 					(reg_q1975 AND symb_decoder(16#15#)) OR
 					(reg_q1975 AND symb_decoder(16#21#)) OR
 					(reg_q1975 AND symb_decoder(16#3f#)) OR
 					(reg_q1975 AND symb_decoder(16#e2#)) OR
 					(reg_q1975 AND symb_decoder(16#c3#)) OR
 					(reg_q1975 AND symb_decoder(16#af#)) OR
 					(reg_q1975 AND symb_decoder(16#22#)) OR
 					(reg_q1975 AND symb_decoder(16#ba#)) OR
 					(reg_q1975 AND symb_decoder(16#f5#)) OR
 					(reg_q1975 AND symb_decoder(16#7d#)) OR
 					(reg_q1975 AND symb_decoder(16#e0#)) OR
 					(reg_q1975 AND symb_decoder(16#7b#)) OR
 					(reg_q1975 AND symb_decoder(16#95#)) OR
 					(reg_q1975 AND symb_decoder(16#cb#)) OR
 					(reg_q1975 AND symb_decoder(16#a0#)) OR
 					(reg_q1975 AND symb_decoder(16#a8#)) OR
 					(reg_q1975 AND symb_decoder(16#8e#)) OR
 					(reg_q1975 AND symb_decoder(16#99#)) OR
 					(reg_q1975 AND symb_decoder(16#76#)) OR
 					(reg_q1975 AND symb_decoder(16#a1#)) OR
 					(reg_q1975 AND symb_decoder(16#57#)) OR
 					(reg_q1975 AND symb_decoder(16#8c#)) OR
 					(reg_q1975 AND symb_decoder(16#78#)) OR
 					(reg_q1975 AND symb_decoder(16#09#)) OR
 					(reg_q1975 AND symb_decoder(16#7a#)) OR
 					(reg_q1975 AND symb_decoder(16#a6#)) OR
 					(reg_q1975 AND symb_decoder(16#1f#)) OR
 					(reg_q1975 AND symb_decoder(16#0b#)) OR
 					(reg_q1975 AND symb_decoder(16#62#)) OR
 					(reg_q1975 AND symb_decoder(16#b6#)) OR
 					(reg_q1975 AND symb_decoder(16#9a#)) OR
 					(reg_q1975 AND symb_decoder(16#52#)) OR
 					(reg_q1975 AND symb_decoder(16#e3#)) OR
 					(reg_q1975 AND symb_decoder(16#42#)) OR
 					(reg_q1975 AND symb_decoder(16#dc#)) OR
 					(reg_q1975 AND symb_decoder(16#34#)) OR
 					(reg_q1975 AND symb_decoder(16#40#)) OR
 					(reg_q1975 AND symb_decoder(16#d5#)) OR
 					(reg_q1975 AND symb_decoder(16#31#)) OR
 					(reg_q1975 AND symb_decoder(16#54#)) OR
 					(reg_q1975 AND symb_decoder(16#06#)) OR
 					(reg_q1975 AND symb_decoder(16#4e#)) OR
 					(reg_q1975 AND symb_decoder(16#7e#)) OR
 					(reg_q1975 AND symb_decoder(16#91#)) OR
 					(reg_q1975 AND symb_decoder(16#47#)) OR
 					(reg_q1975 AND symb_decoder(16#53#)) OR
 					(reg_q1975 AND symb_decoder(16#3c#)) OR
 					(reg_q1975 AND symb_decoder(16#8b#)) OR
 					(reg_q1975 AND symb_decoder(16#ab#)) OR
 					(reg_q1975 AND symb_decoder(16#2f#)) OR
 					(reg_q1975 AND symb_decoder(16#2d#)) OR
 					(reg_q1975 AND symb_decoder(16#13#)) OR
 					(reg_q1975 AND symb_decoder(16#92#)) OR
 					(reg_q1975 AND symb_decoder(16#3d#));
reg_q1686_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q1685 AND symb_decoder(16#0d#)) OR
 					(reg_q1685 AND symb_decoder(16#0a#));
reg_q788_in <= (reg_q786 AND symb_decoder(16#3a#));
reg_q2631_in <= (reg_q2629 AND symb_decoder(16#36#)) OR
 					(reg_q2629 AND symb_decoder(16#33#)) OR
 					(reg_q2629 AND symb_decoder(16#39#)) OR
 					(reg_q2629 AND symb_decoder(16#31#)) OR
 					(reg_q2629 AND symb_decoder(16#38#)) OR
 					(reg_q2629 AND symb_decoder(16#37#)) OR
 					(reg_q2629 AND symb_decoder(16#32#)) OR
 					(reg_q2629 AND symb_decoder(16#35#)) OR
 					(reg_q2629 AND symb_decoder(16#30#)) OR
 					(reg_q2629 AND symb_decoder(16#34#)) OR
 					(reg_q2631 AND symb_decoder(16#33#)) OR
 					(reg_q2631 AND symb_decoder(16#37#)) OR
 					(reg_q2631 AND symb_decoder(16#38#)) OR
 					(reg_q2631 AND symb_decoder(16#34#)) OR
 					(reg_q2631 AND symb_decoder(16#31#)) OR
 					(reg_q2631 AND symb_decoder(16#35#)) OR
 					(reg_q2631 AND symb_decoder(16#32#)) OR
 					(reg_q2631 AND symb_decoder(16#30#)) OR
 					(reg_q2631 AND symb_decoder(16#39#)) OR
 					(reg_q2631 AND symb_decoder(16#36#));
reg_q518_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q517 AND symb_decoder(16#53#)) OR
 					(reg_q517 AND symb_decoder(16#73#));
reg_q474_in <= (reg_q472 AND symb_decoder(16#69#)) OR
 					(reg_q472 AND symb_decoder(16#49#));
reg_q1311_in <= (reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q1310 AND symb_decoder(16#57#)) OR
 					(reg_q1310 AND symb_decoder(16#77#));
reg_q3_in <= (reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2 AND symb_decoder(16#50#)) OR
 					(reg_q2 AND symb_decoder(16#70#));
reg_q118_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q117 AND symb_decoder(16#72#)) OR
 					(reg_q117 AND symb_decoder(16#52#));
reg_q2246_in <= (reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2245 AND symb_decoder(16#2f#));
reg_q476_in <= (reg_q474 AND symb_decoder(16#6e#)) OR
 					(reg_q474 AND symb_decoder(16#4e#));
reg_q763_in <= (reg_q761 AND symb_decoder(16#41#)) OR
 					(reg_q761 AND symb_decoder(16#61#));
reg_q761_in <= (reg_q759 AND symb_decoder(16#74#)) OR
 					(reg_q759 AND symb_decoder(16#54#));
reg_q952_in <= (reg_q950 AND symb_decoder(16#4e#));
reg_q1098_in <= (reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q1097 AND symb_decoder(16#74#)) OR
 					(reg_q1097 AND symb_decoder(16#54#));
reg_q349_in <= (reg_q347 AND symb_decoder(16#65#)) OR
 					(reg_q347 AND symb_decoder(16#45#));
reg_q1909_in <= (reg_q1907 AND symb_decoder(16#54#));
reg_q1147_in <= (reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q1146 AND symb_decoder(16#76#)) OR
 					(reg_q1146 AND symb_decoder(16#56#));
reg_q874_in <= (reg_q872 AND symb_decoder(16#54#)) OR
 					(reg_q872 AND symb_decoder(16#74#));
reg_q1486_in <= (reg_q1484 AND symb_decoder(16#49#)) OR
 					(reg_q1484 AND symb_decoder(16#69#));
reg_q1935_in <= (reg_q2757 AND symb_decoder(16#2a#));
reg_q813_in <= (reg_q811 AND symb_decoder(16#65#)) OR
 					(reg_q811 AND symb_decoder(16#45#));
reg_q815_in <= (reg_q813 AND symb_decoder(16#43#)) OR
 					(reg_q813 AND symb_decoder(16#63#));
reg_q1941_in <= (reg_q1939 AND symb_decoder(16#52#));
reg_q353_in <= (reg_q351 AND symb_decoder(16#76#)) OR
 					(reg_q351 AND symb_decoder(16#56#));
reg_q351_in <= (reg_q349 AND symb_decoder(16#72#)) OR
 					(reg_q349 AND symb_decoder(16#52#));
reg_q1065_in <= (reg_q1063 AND symb_decoder(16#68#)) OR
 					(reg_q1063 AND symb_decoder(16#48#));
reg_q811_in <= (reg_q809 AND symb_decoder(16#6a#)) OR
 					(reg_q809 AND symb_decoder(16#4a#));
reg_q1903_in <= (reg_q1901 AND symb_decoder(16#50#));
reg_q807_in <= (reg_q805 AND symb_decoder(16#55#)) OR
 					(reg_q805 AND symb_decoder(16#75#));
reg_q809_in <= (reg_q807 AND symb_decoder(16#62#)) OR
 					(reg_q807 AND symb_decoder(16#42#));
reg_q1922_in <= (reg_q1920 AND symb_decoder(16#4f#));
reg_fullgraph11_init <= "000000";

reg_fullgraph11_sel <= "00000000000000000000000000000000" & reg_q1922_in & reg_q809_in & reg_q807_in & reg_q1903_in & reg_q811_in & reg_q1065_in & reg_q351_in & reg_q353_in & reg_q1941_in & reg_q815_in & reg_q813_in & reg_q1935_in & reg_q1486_in & reg_q874_in & reg_q1147_in & reg_q1909_in & reg_q349_in & reg_q1098_in & reg_q952_in & reg_q761_in & reg_q763_in & reg_q476_in & reg_q2246_in & reg_q118_in & reg_q3_in & reg_q1311_in & reg_q474_in & reg_q518_in & reg_q2631_in & reg_q788_in & reg_q1686_in & reg_q1975_in;

	--coder fullgraph11
with reg_fullgraph11_sel select
reg_fullgraph11_in <=
	"000001" when "0000000000000000000000000000000000000000000000000000000000000001",
	"000010" when "0000000000000000000000000000000000000000000000000000000000000010",
	"000011" when "0000000000000000000000000000000000000000000000000000000000000100",
	"000100" when "0000000000000000000000000000000000000000000000000000000000001000",
	"000101" when "0000000000000000000000000000000000000000000000000000000000010000",
	"000110" when "0000000000000000000000000000000000000000000000000000000000100000",
	"000111" when "0000000000000000000000000000000000000000000000000000000001000000",
	"001000" when "0000000000000000000000000000000000000000000000000000000010000000",
	"001001" when "0000000000000000000000000000000000000000000000000000000100000000",
	"001010" when "0000000000000000000000000000000000000000000000000000001000000000",
	"001011" when "0000000000000000000000000000000000000000000000000000010000000000",
	"001100" when "0000000000000000000000000000000000000000000000000000100000000000",
	"001101" when "0000000000000000000000000000000000000000000000000001000000000000",
	"001110" when "0000000000000000000000000000000000000000000000000010000000000000",
	"001111" when "0000000000000000000000000000000000000000000000000100000000000000",
	"010000" when "0000000000000000000000000000000000000000000000001000000000000000",
	"010001" when "0000000000000000000000000000000000000000000000010000000000000000",
	"010010" when "0000000000000000000000000000000000000000000000100000000000000000",
	"010011" when "0000000000000000000000000000000000000000000001000000000000000000",
	"010100" when "0000000000000000000000000000000000000000000010000000000000000000",
	"010101" when "0000000000000000000000000000000000000000000100000000000000000000",
	"010110" when "0000000000000000000000000000000000000000001000000000000000000000",
	"010111" when "0000000000000000000000000000000000000000010000000000000000000000",
	"011000" when "0000000000000000000000000000000000000000100000000000000000000000",
	"011001" when "0000000000000000000000000000000000000001000000000000000000000000",
	"011010" when "0000000000000000000000000000000000000010000000000000000000000000",
	"011011" when "0000000000000000000000000000000000000100000000000000000000000000",
	"011100" when "0000000000000000000000000000000000001000000000000000000000000000",
	"011101" when "0000000000000000000000000000000000010000000000000000000000000000",
	"011110" when "0000000000000000000000000000000000100000000000000000000000000000",
	"011111" when "0000000000000000000000000000000001000000000000000000000000000000",
	"100000" when "0000000000000000000000000000000010000000000000000000000000000000",
	"000000" when others;
 --end coder

	p_reg_fullgraph11: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph11 <= reg_fullgraph11_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph11 <= reg_fullgraph11_init;
        else
          reg_fullgraph11 <= reg_fullgraph11_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph11

		reg_q1975 <= '1' when reg_fullgraph11 = "000001" else '0'; 
		reg_q1686 <= '1' when reg_fullgraph11 = "000010" else '0'; 
		reg_q788 <= '1' when reg_fullgraph11 = "000011" else '0'; 
		reg_q2631 <= '1' when reg_fullgraph11 = "000100" else '0'; 
		reg_q518 <= '1' when reg_fullgraph11 = "000101" else '0'; 
		reg_q474 <= '1' when reg_fullgraph11 = "000110" else '0'; 
		reg_q1311 <= '1' when reg_fullgraph11 = "000111" else '0'; 
		reg_q3 <= '1' when reg_fullgraph11 = "001000" else '0'; 
		reg_q118 <= '1' when reg_fullgraph11 = "001001" else '0'; 
		reg_q2246 <= '1' when reg_fullgraph11 = "001010" else '0'; 
		reg_q476 <= '1' when reg_fullgraph11 = "001011" else '0'; 
		reg_q763 <= '1' when reg_fullgraph11 = "001100" else '0'; 
		reg_q761 <= '1' when reg_fullgraph11 = "001101" else '0'; 
		reg_q952 <= '1' when reg_fullgraph11 = "001110" else '0'; 
		reg_q1098 <= '1' when reg_fullgraph11 = "001111" else '0'; 
		reg_q349 <= '1' when reg_fullgraph11 = "010000" else '0'; 
		reg_q1909 <= '1' when reg_fullgraph11 = "010001" else '0'; 
		reg_q1147 <= '1' when reg_fullgraph11 = "010010" else '0'; 
		reg_q874 <= '1' when reg_fullgraph11 = "010011" else '0'; 
		reg_q1486 <= '1' when reg_fullgraph11 = "010100" else '0'; 
		reg_q1935 <= '1' when reg_fullgraph11 = "010101" else '0'; 
		reg_q813 <= '1' when reg_fullgraph11 = "010110" else '0'; 
		reg_q815 <= '1' when reg_fullgraph11 = "010111" else '0'; 
		reg_q1941 <= '1' when reg_fullgraph11 = "011000" else '0'; 
		reg_q353 <= '1' when reg_fullgraph11 = "011001" else '0'; 
		reg_q351 <= '1' when reg_fullgraph11 = "011010" else '0'; 
		reg_q1065 <= '1' when reg_fullgraph11 = "011011" else '0'; 
		reg_q811 <= '1' when reg_fullgraph11 = "011100" else '0'; 
		reg_q1903 <= '1' when reg_fullgraph11 = "011101" else '0'; 
		reg_q807 <= '1' when reg_fullgraph11 = "011110" else '0'; 
		reg_q809 <= '1' when reg_fullgraph11 = "011111" else '0'; 
		reg_q1922 <= '1' when reg_fullgraph11 = "100000" else '0'; 
--end decoder 

reg_q286_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q286 AND symb_decoder(16#ec#)) OR
 					(reg_q286 AND symb_decoder(16#c5#)) OR
 					(reg_q286 AND symb_decoder(16#bf#)) OR
 					(reg_q286 AND symb_decoder(16#38#)) OR
 					(reg_q286 AND symb_decoder(16#b9#)) OR
 					(reg_q286 AND symb_decoder(16#4d#)) OR
 					(reg_q286 AND symb_decoder(16#7f#)) OR
 					(reg_q286 AND symb_decoder(16#ba#)) OR
 					(reg_q286 AND symb_decoder(16#19#)) OR
 					(reg_q286 AND symb_decoder(16#0d#)) OR
 					(reg_q286 AND symb_decoder(16#9e#)) OR
 					(reg_q286 AND symb_decoder(16#f4#)) OR
 					(reg_q286 AND symb_decoder(16#c0#)) OR
 					(reg_q286 AND symb_decoder(16#28#)) OR
 					(reg_q286 AND symb_decoder(16#db#)) OR
 					(reg_q286 AND symb_decoder(16#03#)) OR
 					(reg_q286 AND symb_decoder(16#4c#)) OR
 					(reg_q286 AND symb_decoder(16#bc#)) OR
 					(reg_q286 AND symb_decoder(16#fa#)) OR
 					(reg_q286 AND symb_decoder(16#60#)) OR
 					(reg_q286 AND symb_decoder(16#0b#)) OR
 					(reg_q286 AND symb_decoder(16#82#)) OR
 					(reg_q286 AND symb_decoder(16#b0#)) OR
 					(reg_q286 AND symb_decoder(16#e0#)) OR
 					(reg_q286 AND symb_decoder(16#ac#)) OR
 					(reg_q286 AND symb_decoder(16#4e#)) OR
 					(reg_q286 AND symb_decoder(16#98#)) OR
 					(reg_q286 AND symb_decoder(16#9f#)) OR
 					(reg_q286 AND symb_decoder(16#55#)) OR
 					(reg_q286 AND symb_decoder(16#63#)) OR
 					(reg_q286 AND symb_decoder(16#be#)) OR
 					(reg_q286 AND symb_decoder(16#66#)) OR
 					(reg_q286 AND symb_decoder(16#36#)) OR
 					(reg_q286 AND symb_decoder(16#88#)) OR
 					(reg_q286 AND symb_decoder(16#13#)) OR
 					(reg_q286 AND symb_decoder(16#04#)) OR
 					(reg_q286 AND symb_decoder(16#b3#)) OR
 					(reg_q286 AND symb_decoder(16#a4#)) OR
 					(reg_q286 AND symb_decoder(16#fe#)) OR
 					(reg_q286 AND symb_decoder(16#e8#)) OR
 					(reg_q286 AND symb_decoder(16#9b#)) OR
 					(reg_q286 AND symb_decoder(16#25#)) OR
 					(reg_q286 AND symb_decoder(16#39#)) OR
 					(reg_q286 AND symb_decoder(16#0a#)) OR
 					(reg_q286 AND symb_decoder(16#a6#)) OR
 					(reg_q286 AND symb_decoder(16#1e#)) OR
 					(reg_q286 AND symb_decoder(16#29#)) OR
 					(reg_q286 AND symb_decoder(16#35#)) OR
 					(reg_q286 AND symb_decoder(16#f3#)) OR
 					(reg_q286 AND symb_decoder(16#d6#)) OR
 					(reg_q286 AND symb_decoder(16#08#)) OR
 					(reg_q286 AND symb_decoder(16#a1#)) OR
 					(reg_q286 AND symb_decoder(16#d4#)) OR
 					(reg_q286 AND symb_decoder(16#57#)) OR
 					(reg_q286 AND symb_decoder(16#59#)) OR
 					(reg_q286 AND symb_decoder(16#c3#)) OR
 					(reg_q286 AND symb_decoder(16#b2#)) OR
 					(reg_q286 AND symb_decoder(16#ca#)) OR
 					(reg_q286 AND symb_decoder(16#8b#)) OR
 					(reg_q286 AND symb_decoder(16#dc#)) OR
 					(reg_q286 AND symb_decoder(16#6a#)) OR
 					(reg_q286 AND symb_decoder(16#ee#)) OR
 					(reg_q286 AND symb_decoder(16#90#)) OR
 					(reg_q286 AND symb_decoder(16#1b#)) OR
 					(reg_q286 AND symb_decoder(16#53#)) OR
 					(reg_q286 AND symb_decoder(16#67#)) OR
 					(reg_q286 AND symb_decoder(16#b4#)) OR
 					(reg_q286 AND symb_decoder(16#d1#)) OR
 					(reg_q286 AND symb_decoder(16#c7#)) OR
 					(reg_q286 AND symb_decoder(16#9a#)) OR
 					(reg_q286 AND symb_decoder(16#c2#)) OR
 					(reg_q286 AND symb_decoder(16#74#)) OR
 					(reg_q286 AND symb_decoder(16#f9#)) OR
 					(reg_q286 AND symb_decoder(16#75#)) OR
 					(reg_q286 AND symb_decoder(16#d9#)) OR
 					(reg_q286 AND symb_decoder(16#73#)) OR
 					(reg_q286 AND symb_decoder(16#84#)) OR
 					(reg_q286 AND symb_decoder(16#49#)) OR
 					(reg_q286 AND symb_decoder(16#11#)) OR
 					(reg_q286 AND symb_decoder(16#61#)) OR
 					(reg_q286 AND symb_decoder(16#42#)) OR
 					(reg_q286 AND symb_decoder(16#ef#)) OR
 					(reg_q286 AND symb_decoder(16#94#)) OR
 					(reg_q286 AND symb_decoder(16#77#)) OR
 					(reg_q286 AND symb_decoder(16#3c#)) OR
 					(reg_q286 AND symb_decoder(16#d2#)) OR
 					(reg_q286 AND symb_decoder(16#d5#)) OR
 					(reg_q286 AND symb_decoder(16#16#)) OR
 					(reg_q286 AND symb_decoder(16#f0#)) OR
 					(reg_q286 AND symb_decoder(16#96#)) OR
 					(reg_q286 AND symb_decoder(16#7c#)) OR
 					(reg_q286 AND symb_decoder(16#40#)) OR
 					(reg_q286 AND symb_decoder(16#97#)) OR
 					(reg_q286 AND symb_decoder(16#a9#)) OR
 					(reg_q286 AND symb_decoder(16#a8#)) OR
 					(reg_q286 AND symb_decoder(16#76#)) OR
 					(reg_q286 AND symb_decoder(16#00#)) OR
 					(reg_q286 AND symb_decoder(16#37#)) OR
 					(reg_q286 AND symb_decoder(16#bd#)) OR
 					(reg_q286 AND symb_decoder(16#f1#)) OR
 					(reg_q286 AND symb_decoder(16#17#)) OR
 					(reg_q286 AND symb_decoder(16#a0#)) OR
 					(reg_q286 AND symb_decoder(16#4a#)) OR
 					(reg_q286 AND symb_decoder(16#21#)) OR
 					(reg_q286 AND symb_decoder(16#8c#)) OR
 					(reg_q286 AND symb_decoder(16#0e#)) OR
 					(reg_q286 AND symb_decoder(16#4f#)) OR
 					(reg_q286 AND symb_decoder(16#22#)) OR
 					(reg_q286 AND symb_decoder(16#e9#)) OR
 					(reg_q286 AND symb_decoder(16#d0#)) OR
 					(reg_q286 AND symb_decoder(16#2a#)) OR
 					(reg_q286 AND symb_decoder(16#6b#)) OR
 					(reg_q286 AND symb_decoder(16#5f#)) OR
 					(reg_q286 AND symb_decoder(16#89#)) OR
 					(reg_q286 AND symb_decoder(16#e3#)) OR
 					(reg_q286 AND symb_decoder(16#fb#)) OR
 					(reg_q286 AND symb_decoder(16#14#)) OR
 					(reg_q286 AND symb_decoder(16#da#)) OR
 					(reg_q286 AND symb_decoder(16#7e#)) OR
 					(reg_q286 AND symb_decoder(16#6c#)) OR
 					(reg_q286 AND symb_decoder(16#ed#)) OR
 					(reg_q286 AND symb_decoder(16#62#)) OR
 					(reg_q286 AND symb_decoder(16#c1#)) OR
 					(reg_q286 AND symb_decoder(16#e6#)) OR
 					(reg_q286 AND symb_decoder(16#c9#)) OR
 					(reg_q286 AND symb_decoder(16#b1#)) OR
 					(reg_q286 AND symb_decoder(16#71#)) OR
 					(reg_q286 AND symb_decoder(16#cc#)) OR
 					(reg_q286 AND symb_decoder(16#1f#)) OR
 					(reg_q286 AND symb_decoder(16#0f#)) OR
 					(reg_q286 AND symb_decoder(16#2b#)) OR
 					(reg_q286 AND symb_decoder(16#8e#)) OR
 					(reg_q286 AND symb_decoder(16#3e#)) OR
 					(reg_q286 AND symb_decoder(16#e7#)) OR
 					(reg_q286 AND symb_decoder(16#2d#)) OR
 					(reg_q286 AND symb_decoder(16#f7#)) OR
 					(reg_q286 AND symb_decoder(16#56#)) OR
 					(reg_q286 AND symb_decoder(16#bb#)) OR
 					(reg_q286 AND symb_decoder(16#4b#)) OR
 					(reg_q286 AND symb_decoder(16#69#)) OR
 					(reg_q286 AND symb_decoder(16#5b#)) OR
 					(reg_q286 AND symb_decoder(16#47#)) OR
 					(reg_q286 AND symb_decoder(16#72#)) OR
 					(reg_q286 AND symb_decoder(16#df#)) OR
 					(reg_q286 AND symb_decoder(16#f6#)) OR
 					(reg_q286 AND symb_decoder(16#80#)) OR
 					(reg_q286 AND symb_decoder(16#30#)) OR
 					(reg_q286 AND symb_decoder(16#8f#)) OR
 					(reg_q286 AND symb_decoder(16#cf#)) OR
 					(reg_q286 AND symb_decoder(16#b8#)) OR
 					(reg_q286 AND symb_decoder(16#c6#)) OR
 					(reg_q286 AND symb_decoder(16#93#)) OR
 					(reg_q286 AND symb_decoder(16#91#)) OR
 					(reg_q286 AND symb_decoder(16#27#)) OR
 					(reg_q286 AND symb_decoder(16#65#)) OR
 					(reg_q286 AND symb_decoder(16#af#)) OR
 					(reg_q286 AND symb_decoder(16#ff#)) OR
 					(reg_q286 AND symb_decoder(16#2e#)) OR
 					(reg_q286 AND symb_decoder(16#3d#)) OR
 					(reg_q286 AND symb_decoder(16#2c#)) OR
 					(reg_q286 AND symb_decoder(16#51#)) OR
 					(reg_q286 AND symb_decoder(16#b6#)) OR
 					(reg_q286 AND symb_decoder(16#32#)) OR
 					(reg_q286 AND symb_decoder(16#b5#)) OR
 					(reg_q286 AND symb_decoder(16#5c#)) OR
 					(reg_q286 AND symb_decoder(16#de#)) OR
 					(reg_q286 AND symb_decoder(16#43#)) OR
 					(reg_q286 AND symb_decoder(16#3f#)) OR
 					(reg_q286 AND symb_decoder(16#01#)) OR
 					(reg_q286 AND symb_decoder(16#e4#)) OR
 					(reg_q286 AND symb_decoder(16#45#)) OR
 					(reg_q286 AND symb_decoder(16#f8#)) OR
 					(reg_q286 AND symb_decoder(16#cd#)) OR
 					(reg_q286 AND symb_decoder(16#b7#)) OR
 					(reg_q286 AND symb_decoder(16#5d#)) OR
 					(reg_q286 AND symb_decoder(16#c8#)) OR
 					(reg_q286 AND symb_decoder(16#99#)) OR
 					(reg_q286 AND symb_decoder(16#a5#)) OR
 					(reg_q286 AND symb_decoder(16#7b#)) OR
 					(reg_q286 AND symb_decoder(16#50#)) OR
 					(reg_q286 AND symb_decoder(16#ad#)) OR
 					(reg_q286 AND symb_decoder(16#05#)) OR
 					(reg_q286 AND symb_decoder(16#1c#)) OR
 					(reg_q286 AND symb_decoder(16#d7#)) OR
 					(reg_q286 AND symb_decoder(16#52#)) OR
 					(reg_q286 AND symb_decoder(16#87#)) OR
 					(reg_q286 AND symb_decoder(16#10#)) OR
 					(reg_q286 AND symb_decoder(16#5a#)) OR
 					(reg_q286 AND symb_decoder(16#54#)) OR
 					(reg_q286 AND symb_decoder(16#12#)) OR
 					(reg_q286 AND symb_decoder(16#09#)) OR
 					(reg_q286 AND symb_decoder(16#07#)) OR
 					(reg_q286 AND symb_decoder(16#a3#)) OR
 					(reg_q286 AND symb_decoder(16#15#)) OR
 					(reg_q286 AND symb_decoder(16#81#)) OR
 					(reg_q286 AND symb_decoder(16#18#)) OR
 					(reg_q286 AND symb_decoder(16#6f#)) OR
 					(reg_q286 AND symb_decoder(16#ea#)) OR
 					(reg_q286 AND symb_decoder(16#68#)) OR
 					(reg_q286 AND symb_decoder(16#48#)) OR
 					(reg_q286 AND symb_decoder(16#8a#)) OR
 					(reg_q286 AND symb_decoder(16#92#)) OR
 					(reg_q286 AND symb_decoder(16#85#)) OR
 					(reg_q286 AND symb_decoder(16#26#)) OR
 					(reg_q286 AND symb_decoder(16#f5#)) OR
 					(reg_q286 AND symb_decoder(16#06#)) OR
 					(reg_q286 AND symb_decoder(16#7d#)) OR
 					(reg_q286 AND symb_decoder(16#eb#)) OR
 					(reg_q286 AND symb_decoder(16#0c#)) OR
 					(reg_q286 AND symb_decoder(16#46#)) OR
 					(reg_q286 AND symb_decoder(16#ce#)) OR
 					(reg_q286 AND symb_decoder(16#78#)) OR
 					(reg_q286 AND symb_decoder(16#70#)) OR
 					(reg_q286 AND symb_decoder(16#3a#)) OR
 					(reg_q286 AND symb_decoder(16#33#)) OR
 					(reg_q286 AND symb_decoder(16#fd#)) OR
 					(reg_q286 AND symb_decoder(16#3b#)) OR
 					(reg_q286 AND symb_decoder(16#64#)) OR
 					(reg_q286 AND symb_decoder(16#6e#)) OR
 					(reg_q286 AND symb_decoder(16#f2#)) OR
 					(reg_q286 AND symb_decoder(16#ae#)) OR
 					(reg_q286 AND symb_decoder(16#ab#)) OR
 					(reg_q286 AND symb_decoder(16#23#)) OR
 					(reg_q286 AND symb_decoder(16#d3#)) OR
 					(reg_q286 AND symb_decoder(16#9d#)) OR
 					(reg_q286 AND symb_decoder(16#dd#)) OR
 					(reg_q286 AND symb_decoder(16#41#)) OR
 					(reg_q286 AND symb_decoder(16#a2#)) OR
 					(reg_q286 AND symb_decoder(16#e1#)) OR
 					(reg_q286 AND symb_decoder(16#24#)) OR
 					(reg_q286 AND symb_decoder(16#20#)) OR
 					(reg_q286 AND symb_decoder(16#1a#)) OR
 					(reg_q286 AND symb_decoder(16#c4#)) OR
 					(reg_q286 AND symb_decoder(16#58#)) OR
 					(reg_q286 AND symb_decoder(16#02#)) OR
 					(reg_q286 AND symb_decoder(16#34#)) OR
 					(reg_q286 AND symb_decoder(16#95#)) OR
 					(reg_q286 AND symb_decoder(16#31#)) OR
 					(reg_q286 AND symb_decoder(16#86#)) OR
 					(reg_q286 AND symb_decoder(16#cb#)) OR
 					(reg_q286 AND symb_decoder(16#a7#)) OR
 					(reg_q286 AND symb_decoder(16#2f#)) OR
 					(reg_q286 AND symb_decoder(16#6d#)) OR
 					(reg_q286 AND symb_decoder(16#aa#)) OR
 					(reg_q286 AND symb_decoder(16#e5#)) OR
 					(reg_q286 AND symb_decoder(16#1d#)) OR
 					(reg_q286 AND symb_decoder(16#d8#)) OR
 					(reg_q286 AND symb_decoder(16#83#)) OR
 					(reg_q286 AND symb_decoder(16#7a#)) OR
 					(reg_q286 AND symb_decoder(16#e2#)) OR
 					(reg_q286 AND symb_decoder(16#79#)) OR
 					(reg_q286 AND symb_decoder(16#44#)) OR
 					(reg_q286 AND symb_decoder(16#fc#)) OR
 					(reg_q286 AND symb_decoder(16#8d#)) OR
 					(reg_q286 AND symb_decoder(16#9c#)) OR
 					(reg_q286 AND symb_decoder(16#5e#));
reg_q286_init <= '0' ;
	p_reg_q286: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q286 <= reg_q286_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q286 <= reg_q286_init;
        else
          reg_q286 <= reg_q286_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1309_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1309 AND symb_decoder(16#ce#)) OR
 					(reg_q1309 AND symb_decoder(16#de#)) OR
 					(reg_q1309 AND symb_decoder(16#04#)) OR
 					(reg_q1309 AND symb_decoder(16#01#)) OR
 					(reg_q1309 AND symb_decoder(16#32#)) OR
 					(reg_q1309 AND symb_decoder(16#80#)) OR
 					(reg_q1309 AND symb_decoder(16#54#)) OR
 					(reg_q1309 AND symb_decoder(16#40#)) OR
 					(reg_q1309 AND symb_decoder(16#6c#)) OR
 					(reg_q1309 AND symb_decoder(16#a7#)) OR
 					(reg_q1309 AND symb_decoder(16#e0#)) OR
 					(reg_q1309 AND symb_decoder(16#8a#)) OR
 					(reg_q1309 AND symb_decoder(16#75#)) OR
 					(reg_q1309 AND symb_decoder(16#1e#)) OR
 					(reg_q1309 AND symb_decoder(16#62#)) OR
 					(reg_q1309 AND symb_decoder(16#9d#)) OR
 					(reg_q1309 AND symb_decoder(16#74#)) OR
 					(reg_q1309 AND symb_decoder(16#65#)) OR
 					(reg_q1309 AND symb_decoder(16#b8#)) OR
 					(reg_q1309 AND symb_decoder(16#9f#)) OR
 					(reg_q1309 AND symb_decoder(16#bb#)) OR
 					(reg_q1309 AND symb_decoder(16#0d#)) OR
 					(reg_q1309 AND symb_decoder(16#a1#)) OR
 					(reg_q1309 AND symb_decoder(16#64#)) OR
 					(reg_q1309 AND symb_decoder(16#f6#)) OR
 					(reg_q1309 AND symb_decoder(16#c5#)) OR
 					(reg_q1309 AND symb_decoder(16#33#)) OR
 					(reg_q1309 AND symb_decoder(16#d8#)) OR
 					(reg_q1309 AND symb_decoder(16#34#)) OR
 					(reg_q1309 AND symb_decoder(16#ab#)) OR
 					(reg_q1309 AND symb_decoder(16#d6#)) OR
 					(reg_q1309 AND symb_decoder(16#45#)) OR
 					(reg_q1309 AND symb_decoder(16#c4#)) OR
 					(reg_q1309 AND symb_decoder(16#6f#)) OR
 					(reg_q1309 AND symb_decoder(16#bd#)) OR
 					(reg_q1309 AND symb_decoder(16#36#)) OR
 					(reg_q1309 AND symb_decoder(16#51#)) OR
 					(reg_q1309 AND symb_decoder(16#be#)) OR
 					(reg_q1309 AND symb_decoder(16#58#)) OR
 					(reg_q1309 AND symb_decoder(16#0f#)) OR
 					(reg_q1309 AND symb_decoder(16#b7#)) OR
 					(reg_q1309 AND symb_decoder(16#7e#)) OR
 					(reg_q1309 AND symb_decoder(16#f9#)) OR
 					(reg_q1309 AND symb_decoder(16#d9#)) OR
 					(reg_q1309 AND symb_decoder(16#52#)) OR
 					(reg_q1309 AND symb_decoder(16#41#)) OR
 					(reg_q1309 AND symb_decoder(16#18#)) OR
 					(reg_q1309 AND symb_decoder(16#73#)) OR
 					(reg_q1309 AND symb_decoder(16#3a#)) OR
 					(reg_q1309 AND symb_decoder(16#15#)) OR
 					(reg_q1309 AND symb_decoder(16#1b#)) OR
 					(reg_q1309 AND symb_decoder(16#16#)) OR
 					(reg_q1309 AND symb_decoder(16#76#)) OR
 					(reg_q1309 AND symb_decoder(16#b9#)) OR
 					(reg_q1309 AND symb_decoder(16#10#)) OR
 					(reg_q1309 AND symb_decoder(16#c7#)) OR
 					(reg_q1309 AND symb_decoder(16#a6#)) OR
 					(reg_q1309 AND symb_decoder(16#a3#)) OR
 					(reg_q1309 AND symb_decoder(16#42#)) OR
 					(reg_q1309 AND symb_decoder(16#38#)) OR
 					(reg_q1309 AND symb_decoder(16#49#)) OR
 					(reg_q1309 AND symb_decoder(16#db#)) OR
 					(reg_q1309 AND symb_decoder(16#83#)) OR
 					(reg_q1309 AND symb_decoder(16#d2#)) OR
 					(reg_q1309 AND symb_decoder(16#78#)) OR
 					(reg_q1309 AND symb_decoder(16#aa#)) OR
 					(reg_q1309 AND symb_decoder(16#5b#)) OR
 					(reg_q1309 AND symb_decoder(16#f7#)) OR
 					(reg_q1309 AND symb_decoder(16#8f#)) OR
 					(reg_q1309 AND symb_decoder(16#09#)) OR
 					(reg_q1309 AND symb_decoder(16#5e#)) OR
 					(reg_q1309 AND symb_decoder(16#af#)) OR
 					(reg_q1309 AND symb_decoder(16#cf#)) OR
 					(reg_q1309 AND symb_decoder(16#cd#)) OR
 					(reg_q1309 AND symb_decoder(16#e5#)) OR
 					(reg_q1309 AND symb_decoder(16#97#)) OR
 					(reg_q1309 AND symb_decoder(16#d7#)) OR
 					(reg_q1309 AND symb_decoder(16#2b#)) OR
 					(reg_q1309 AND symb_decoder(16#37#)) OR
 					(reg_q1309 AND symb_decoder(16#8c#)) OR
 					(reg_q1309 AND symb_decoder(16#fd#)) OR
 					(reg_q1309 AND symb_decoder(16#17#)) OR
 					(reg_q1309 AND symb_decoder(16#7d#)) OR
 					(reg_q1309 AND symb_decoder(16#23#)) OR
 					(reg_q1309 AND symb_decoder(16#1a#)) OR
 					(reg_q1309 AND symb_decoder(16#da#)) OR
 					(reg_q1309 AND symb_decoder(16#70#)) OR
 					(reg_q1309 AND symb_decoder(16#96#)) OR
 					(reg_q1309 AND symb_decoder(16#1d#)) OR
 					(reg_q1309 AND symb_decoder(16#5d#)) OR
 					(reg_q1309 AND symb_decoder(16#ed#)) OR
 					(reg_q1309 AND symb_decoder(16#b5#)) OR
 					(reg_q1309 AND symb_decoder(16#c0#)) OR
 					(reg_q1309 AND symb_decoder(16#9b#)) OR
 					(reg_q1309 AND symb_decoder(16#06#)) OR
 					(reg_q1309 AND symb_decoder(16#5c#)) OR
 					(reg_q1309 AND symb_decoder(16#94#)) OR
 					(reg_q1309 AND symb_decoder(16#8b#)) OR
 					(reg_q1309 AND symb_decoder(16#4d#)) OR
 					(reg_q1309 AND symb_decoder(16#28#)) OR
 					(reg_q1309 AND symb_decoder(16#93#)) OR
 					(reg_q1309 AND symb_decoder(16#66#)) OR
 					(reg_q1309 AND symb_decoder(16#50#)) OR
 					(reg_q1309 AND symb_decoder(16#ee#)) OR
 					(reg_q1309 AND symb_decoder(16#88#)) OR
 					(reg_q1309 AND symb_decoder(16#46#)) OR
 					(reg_q1309 AND symb_decoder(16#c8#)) OR
 					(reg_q1309 AND symb_decoder(16#4e#)) OR
 					(reg_q1309 AND symb_decoder(16#56#)) OR
 					(reg_q1309 AND symb_decoder(16#ad#)) OR
 					(reg_q1309 AND symb_decoder(16#d3#)) OR
 					(reg_q1309 AND symb_decoder(16#07#)) OR
 					(reg_q1309 AND symb_decoder(16#cb#)) OR
 					(reg_q1309 AND symb_decoder(16#1f#)) OR
 					(reg_q1309 AND symb_decoder(16#02#)) OR
 					(reg_q1309 AND symb_decoder(16#a4#)) OR
 					(reg_q1309 AND symb_decoder(16#f4#)) OR
 					(reg_q1309 AND symb_decoder(16#21#)) OR
 					(reg_q1309 AND symb_decoder(16#44#)) OR
 					(reg_q1309 AND symb_decoder(16#82#)) OR
 					(reg_q1309 AND symb_decoder(16#ef#)) OR
 					(reg_q1309 AND symb_decoder(16#8d#)) OR
 					(reg_q1309 AND symb_decoder(16#c9#)) OR
 					(reg_q1309 AND symb_decoder(16#f8#)) OR
 					(reg_q1309 AND symb_decoder(16#89#)) OR
 					(reg_q1309 AND symb_decoder(16#5a#)) OR
 					(reg_q1309 AND symb_decoder(16#ca#)) OR
 					(reg_q1309 AND symb_decoder(16#e3#)) OR
 					(reg_q1309 AND symb_decoder(16#4b#)) OR
 					(reg_q1309 AND symb_decoder(16#61#)) OR
 					(reg_q1309 AND symb_decoder(16#b2#)) OR
 					(reg_q1309 AND symb_decoder(16#dd#)) OR
 					(reg_q1309 AND symb_decoder(16#91#)) OR
 					(reg_q1309 AND symb_decoder(16#57#)) OR
 					(reg_q1309 AND symb_decoder(16#c1#)) OR
 					(reg_q1309 AND symb_decoder(16#fb#)) OR
 					(reg_q1309 AND symb_decoder(16#e7#)) OR
 					(reg_q1309 AND symb_decoder(16#0b#)) OR
 					(reg_q1309 AND symb_decoder(16#cc#)) OR
 					(reg_q1309 AND symb_decoder(16#43#)) OR
 					(reg_q1309 AND symb_decoder(16#71#)) OR
 					(reg_q1309 AND symb_decoder(16#6a#)) OR
 					(reg_q1309 AND symb_decoder(16#35#)) OR
 					(reg_q1309 AND symb_decoder(16#e6#)) OR
 					(reg_q1309 AND symb_decoder(16#b0#)) OR
 					(reg_q1309 AND symb_decoder(16#fc#)) OR
 					(reg_q1309 AND symb_decoder(16#3d#)) OR
 					(reg_q1309 AND symb_decoder(16#3f#)) OR
 					(reg_q1309 AND symb_decoder(16#30#)) OR
 					(reg_q1309 AND symb_decoder(16#a9#)) OR
 					(reg_q1309 AND symb_decoder(16#13#)) OR
 					(reg_q1309 AND symb_decoder(16#ba#)) OR
 					(reg_q1309 AND symb_decoder(16#98#)) OR
 					(reg_q1309 AND symb_decoder(16#69#)) OR
 					(reg_q1309 AND symb_decoder(16#29#)) OR
 					(reg_q1309 AND symb_decoder(16#53#)) OR
 					(reg_q1309 AND symb_decoder(16#d0#)) OR
 					(reg_q1309 AND symb_decoder(16#bf#)) OR
 					(reg_q1309 AND symb_decoder(16#77#)) OR
 					(reg_q1309 AND symb_decoder(16#39#)) OR
 					(reg_q1309 AND symb_decoder(16#dc#)) OR
 					(reg_q1309 AND symb_decoder(16#b3#)) OR
 					(reg_q1309 AND symb_decoder(16#d4#)) OR
 					(reg_q1309 AND symb_decoder(16#2d#)) OR
 					(reg_q1309 AND symb_decoder(16#ff#)) OR
 					(reg_q1309 AND symb_decoder(16#7f#)) OR
 					(reg_q1309 AND symb_decoder(16#05#)) OR
 					(reg_q1309 AND symb_decoder(16#7b#)) OR
 					(reg_q1309 AND symb_decoder(16#f1#)) OR
 					(reg_q1309 AND symb_decoder(16#79#)) OR
 					(reg_q1309 AND symb_decoder(16#7c#)) OR
 					(reg_q1309 AND symb_decoder(16#bc#)) OR
 					(reg_q1309 AND symb_decoder(16#a5#)) OR
 					(reg_q1309 AND symb_decoder(16#9e#)) OR
 					(reg_q1309 AND symb_decoder(16#4c#)) OR
 					(reg_q1309 AND symb_decoder(16#eb#)) OR
 					(reg_q1309 AND symb_decoder(16#a8#)) OR
 					(reg_q1309 AND symb_decoder(16#5f#)) OR
 					(reg_q1309 AND symb_decoder(16#68#)) OR
 					(reg_q1309 AND symb_decoder(16#fe#)) OR
 					(reg_q1309 AND symb_decoder(16#47#)) OR
 					(reg_q1309 AND symb_decoder(16#86#)) OR
 					(reg_q1309 AND symb_decoder(16#0e#)) OR
 					(reg_q1309 AND symb_decoder(16#92#)) OR
 					(reg_q1309 AND symb_decoder(16#60#)) OR
 					(reg_q1309 AND symb_decoder(16#14#)) OR
 					(reg_q1309 AND symb_decoder(16#f0#)) OR
 					(reg_q1309 AND symb_decoder(16#9c#)) OR
 					(reg_q1309 AND symb_decoder(16#1c#)) OR
 					(reg_q1309 AND symb_decoder(16#2f#)) OR
 					(reg_q1309 AND symb_decoder(16#12#)) OR
 					(reg_q1309 AND symb_decoder(16#03#)) OR
 					(reg_q1309 AND symb_decoder(16#6b#)) OR
 					(reg_q1309 AND symb_decoder(16#e8#)) OR
 					(reg_q1309 AND symb_decoder(16#ec#)) OR
 					(reg_q1309 AND symb_decoder(16#72#)) OR
 					(reg_q1309 AND symb_decoder(16#11#)) OR
 					(reg_q1309 AND symb_decoder(16#d1#)) OR
 					(reg_q1309 AND symb_decoder(16#c2#)) OR
 					(reg_q1309 AND symb_decoder(16#20#)) OR
 					(reg_q1309 AND symb_decoder(16#0a#)) OR
 					(reg_q1309 AND symb_decoder(16#95#)) OR
 					(reg_q1309 AND symb_decoder(16#d5#)) OR
 					(reg_q1309 AND symb_decoder(16#2e#)) OR
 					(reg_q1309 AND symb_decoder(16#4f#)) OR
 					(reg_q1309 AND symb_decoder(16#59#)) OR
 					(reg_q1309 AND symb_decoder(16#87#)) OR
 					(reg_q1309 AND symb_decoder(16#a0#)) OR
 					(reg_q1309 AND symb_decoder(16#3b#)) OR
 					(reg_q1309 AND symb_decoder(16#84#)) OR
 					(reg_q1309 AND symb_decoder(16#63#)) OR
 					(reg_q1309 AND symb_decoder(16#fa#)) OR
 					(reg_q1309 AND symb_decoder(16#90#)) OR
 					(reg_q1309 AND symb_decoder(16#b1#)) OR
 					(reg_q1309 AND symb_decoder(16#e4#)) OR
 					(reg_q1309 AND symb_decoder(16#4a#)) OR
 					(reg_q1309 AND symb_decoder(16#6e#)) OR
 					(reg_q1309 AND symb_decoder(16#24#)) OR
 					(reg_q1309 AND symb_decoder(16#c3#)) OR
 					(reg_q1309 AND symb_decoder(16#0c#)) OR
 					(reg_q1309 AND symb_decoder(16#c6#)) OR
 					(reg_q1309 AND symb_decoder(16#08#)) OR
 					(reg_q1309 AND symb_decoder(16#a2#)) OR
 					(reg_q1309 AND symb_decoder(16#9a#)) OR
 					(reg_q1309 AND symb_decoder(16#19#)) OR
 					(reg_q1309 AND symb_decoder(16#81#)) OR
 					(reg_q1309 AND symb_decoder(16#e1#)) OR
 					(reg_q1309 AND symb_decoder(16#b4#)) OR
 					(reg_q1309 AND symb_decoder(16#25#)) OR
 					(reg_q1309 AND symb_decoder(16#85#)) OR
 					(reg_q1309 AND symb_decoder(16#f2#)) OR
 					(reg_q1309 AND symb_decoder(16#ae#)) OR
 					(reg_q1309 AND symb_decoder(16#67#)) OR
 					(reg_q1309 AND symb_decoder(16#ea#)) OR
 					(reg_q1309 AND symb_decoder(16#f3#)) OR
 					(reg_q1309 AND symb_decoder(16#b6#)) OR
 					(reg_q1309 AND symb_decoder(16#df#)) OR
 					(reg_q1309 AND symb_decoder(16#e2#)) OR
 					(reg_q1309 AND symb_decoder(16#2a#)) OR
 					(reg_q1309 AND symb_decoder(16#00#)) OR
 					(reg_q1309 AND symb_decoder(16#48#)) OR
 					(reg_q1309 AND symb_decoder(16#55#)) OR
 					(reg_q1309 AND symb_decoder(16#ac#)) OR
 					(reg_q1309 AND symb_decoder(16#3c#)) OR
 					(reg_q1309 AND symb_decoder(16#7a#)) OR
 					(reg_q1309 AND symb_decoder(16#6d#)) OR
 					(reg_q1309 AND symb_decoder(16#31#)) OR
 					(reg_q1309 AND symb_decoder(16#f5#)) OR
 					(reg_q1309 AND symb_decoder(16#8e#)) OR
 					(reg_q1309 AND symb_decoder(16#3e#)) OR
 					(reg_q1309 AND symb_decoder(16#26#)) OR
 					(reg_q1309 AND symb_decoder(16#2c#)) OR
 					(reg_q1309 AND symb_decoder(16#e9#)) OR
 					(reg_q1309 AND symb_decoder(16#27#)) OR
 					(reg_q1309 AND symb_decoder(16#99#)) OR
 					(reg_q1309 AND symb_decoder(16#22#));
reg_q1309_init <= '0' ;
	p_reg_q1309: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1309 <= reg_q1309_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1309 <= reg_q1309_init;
        else
          reg_q1309 <= reg_q1309_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2244_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q2244 AND symb_decoder(16#e0#)) OR
 					(reg_q2244 AND symb_decoder(16#f8#)) OR
 					(reg_q2244 AND symb_decoder(16#50#)) OR
 					(reg_q2244 AND symb_decoder(16#5a#)) OR
 					(reg_q2244 AND symb_decoder(16#f7#)) OR
 					(reg_q2244 AND symb_decoder(16#61#)) OR
 					(reg_q2244 AND symb_decoder(16#8e#)) OR
 					(reg_q2244 AND symb_decoder(16#05#)) OR
 					(reg_q2244 AND symb_decoder(16#16#)) OR
 					(reg_q2244 AND symb_decoder(16#8f#)) OR
 					(reg_q2244 AND symb_decoder(16#59#)) OR
 					(reg_q2244 AND symb_decoder(16#0c#)) OR
 					(reg_q2244 AND symb_decoder(16#02#)) OR
 					(reg_q2244 AND symb_decoder(16#54#)) OR
 					(reg_q2244 AND symb_decoder(16#36#)) OR
 					(reg_q2244 AND symb_decoder(16#8a#)) OR
 					(reg_q2244 AND symb_decoder(16#76#)) OR
 					(reg_q2244 AND symb_decoder(16#bc#)) OR
 					(reg_q2244 AND symb_decoder(16#c2#)) OR
 					(reg_q2244 AND symb_decoder(16#53#)) OR
 					(reg_q2244 AND symb_decoder(16#3f#)) OR
 					(reg_q2244 AND symb_decoder(16#fd#)) OR
 					(reg_q2244 AND symb_decoder(16#c4#)) OR
 					(reg_q2244 AND symb_decoder(16#bf#)) OR
 					(reg_q2244 AND symb_decoder(16#4b#)) OR
 					(reg_q2244 AND symb_decoder(16#bb#)) OR
 					(reg_q2244 AND symb_decoder(16#29#)) OR
 					(reg_q2244 AND symb_decoder(16#95#)) OR
 					(reg_q2244 AND symb_decoder(16#a6#)) OR
 					(reg_q2244 AND symb_decoder(16#b5#)) OR
 					(reg_q2244 AND symb_decoder(16#e9#)) OR
 					(reg_q2244 AND symb_decoder(16#fa#)) OR
 					(reg_q2244 AND symb_decoder(16#27#)) OR
 					(reg_q2244 AND symb_decoder(16#08#)) OR
 					(reg_q2244 AND symb_decoder(16#89#)) OR
 					(reg_q2244 AND symb_decoder(16#47#)) OR
 					(reg_q2244 AND symb_decoder(16#e5#)) OR
 					(reg_q2244 AND symb_decoder(16#af#)) OR
 					(reg_q2244 AND symb_decoder(16#0a#)) OR
 					(reg_q2244 AND symb_decoder(16#b2#)) OR
 					(reg_q2244 AND symb_decoder(16#a4#)) OR
 					(reg_q2244 AND symb_decoder(16#1d#)) OR
 					(reg_q2244 AND symb_decoder(16#85#)) OR
 					(reg_q2244 AND symb_decoder(16#b6#)) OR
 					(reg_q2244 AND symb_decoder(16#6d#)) OR
 					(reg_q2244 AND symb_decoder(16#10#)) OR
 					(reg_q2244 AND symb_decoder(16#23#)) OR
 					(reg_q2244 AND symb_decoder(16#c6#)) OR
 					(reg_q2244 AND symb_decoder(16#e7#)) OR
 					(reg_q2244 AND symb_decoder(16#0b#)) OR
 					(reg_q2244 AND symb_decoder(16#c0#)) OR
 					(reg_q2244 AND symb_decoder(16#ff#)) OR
 					(reg_q2244 AND symb_decoder(16#35#)) OR
 					(reg_q2244 AND symb_decoder(16#93#)) OR
 					(reg_q2244 AND symb_decoder(16#18#)) OR
 					(reg_q2244 AND symb_decoder(16#71#)) OR
 					(reg_q2244 AND symb_decoder(16#a3#)) OR
 					(reg_q2244 AND symb_decoder(16#1c#)) OR
 					(reg_q2244 AND symb_decoder(16#14#)) OR
 					(reg_q2244 AND symb_decoder(16#2a#)) OR
 					(reg_q2244 AND symb_decoder(16#7e#)) OR
 					(reg_q2244 AND symb_decoder(16#1e#)) OR
 					(reg_q2244 AND symb_decoder(16#a7#)) OR
 					(reg_q2244 AND symb_decoder(16#38#)) OR
 					(reg_q2244 AND symb_decoder(16#6e#)) OR
 					(reg_q2244 AND symb_decoder(16#40#)) OR
 					(reg_q2244 AND symb_decoder(16#8c#)) OR
 					(reg_q2244 AND symb_decoder(16#99#)) OR
 					(reg_q2244 AND symb_decoder(16#c8#)) OR
 					(reg_q2244 AND symb_decoder(16#c9#)) OR
 					(reg_q2244 AND symb_decoder(16#a8#)) OR
 					(reg_q2244 AND symb_decoder(16#13#)) OR
 					(reg_q2244 AND symb_decoder(16#f5#)) OR
 					(reg_q2244 AND symb_decoder(16#75#)) OR
 					(reg_q2244 AND symb_decoder(16#aa#)) OR
 					(reg_q2244 AND symb_decoder(16#11#)) OR
 					(reg_q2244 AND symb_decoder(16#1f#)) OR
 					(reg_q2244 AND symb_decoder(16#3b#)) OR
 					(reg_q2244 AND symb_decoder(16#65#)) OR
 					(reg_q2244 AND symb_decoder(16#3c#)) OR
 					(reg_q2244 AND symb_decoder(16#49#)) OR
 					(reg_q2244 AND symb_decoder(16#37#)) OR
 					(reg_q2244 AND symb_decoder(16#7d#)) OR
 					(reg_q2244 AND symb_decoder(16#84#)) OR
 					(reg_q2244 AND symb_decoder(16#30#)) OR
 					(reg_q2244 AND symb_decoder(16#cd#)) OR
 					(reg_q2244 AND symb_decoder(16#31#)) OR
 					(reg_q2244 AND symb_decoder(16#d1#)) OR
 					(reg_q2244 AND symb_decoder(16#78#)) OR
 					(reg_q2244 AND symb_decoder(16#ed#)) OR
 					(reg_q2244 AND symb_decoder(16#6c#)) OR
 					(reg_q2244 AND symb_decoder(16#c5#)) OR
 					(reg_q2244 AND symb_decoder(16#83#)) OR
 					(reg_q2244 AND symb_decoder(16#9f#)) OR
 					(reg_q2244 AND symb_decoder(16#f1#)) OR
 					(reg_q2244 AND symb_decoder(16#ac#)) OR
 					(reg_q2244 AND symb_decoder(16#ab#)) OR
 					(reg_q2244 AND symb_decoder(16#d2#)) OR
 					(reg_q2244 AND symb_decoder(16#6b#)) OR
 					(reg_q2244 AND symb_decoder(16#c7#)) OR
 					(reg_q2244 AND symb_decoder(16#60#)) OR
 					(reg_q2244 AND symb_decoder(16#ca#)) OR
 					(reg_q2244 AND symb_decoder(16#2c#)) OR
 					(reg_q2244 AND symb_decoder(16#9a#)) OR
 					(reg_q2244 AND symb_decoder(16#06#)) OR
 					(reg_q2244 AND symb_decoder(16#7c#)) OR
 					(reg_q2244 AND symb_decoder(16#79#)) OR
 					(reg_q2244 AND symb_decoder(16#a2#)) OR
 					(reg_q2244 AND symb_decoder(16#2d#)) OR
 					(reg_q2244 AND symb_decoder(16#d3#)) OR
 					(reg_q2244 AND symb_decoder(16#7f#)) OR
 					(reg_q2244 AND symb_decoder(16#e1#)) OR
 					(reg_q2244 AND symb_decoder(16#24#)) OR
 					(reg_q2244 AND symb_decoder(16#17#)) OR
 					(reg_q2244 AND symb_decoder(16#dd#)) OR
 					(reg_q2244 AND symb_decoder(16#00#)) OR
 					(reg_q2244 AND symb_decoder(16#ad#)) OR
 					(reg_q2244 AND symb_decoder(16#2b#)) OR
 					(reg_q2244 AND symb_decoder(16#c1#)) OR
 					(reg_q2244 AND symb_decoder(16#6f#)) OR
 					(reg_q2244 AND symb_decoder(16#07#)) OR
 					(reg_q2244 AND symb_decoder(16#ba#)) OR
 					(reg_q2244 AND symb_decoder(16#fe#)) OR
 					(reg_q2244 AND symb_decoder(16#eb#)) OR
 					(reg_q2244 AND symb_decoder(16#f6#)) OR
 					(reg_q2244 AND symb_decoder(16#d6#)) OR
 					(reg_q2244 AND symb_decoder(16#f2#)) OR
 					(reg_q2244 AND symb_decoder(16#f4#)) OR
 					(reg_q2244 AND symb_decoder(16#94#)) OR
 					(reg_q2244 AND symb_decoder(16#0f#)) OR
 					(reg_q2244 AND symb_decoder(16#0d#)) OR
 					(reg_q2244 AND symb_decoder(16#e4#)) OR
 					(reg_q2244 AND symb_decoder(16#0e#)) OR
 					(reg_q2244 AND symb_decoder(16#cb#)) OR
 					(reg_q2244 AND symb_decoder(16#48#)) OR
 					(reg_q2244 AND symb_decoder(16#34#)) OR
 					(reg_q2244 AND symb_decoder(16#70#)) OR
 					(reg_q2244 AND symb_decoder(16#03#)) OR
 					(reg_q2244 AND symb_decoder(16#4d#)) OR
 					(reg_q2244 AND symb_decoder(16#15#)) OR
 					(reg_q2244 AND symb_decoder(16#ae#)) OR
 					(reg_q2244 AND symb_decoder(16#33#)) OR
 					(reg_q2244 AND symb_decoder(16#4c#)) OR
 					(reg_q2244 AND symb_decoder(16#28#)) OR
 					(reg_q2244 AND symb_decoder(16#be#)) OR
 					(reg_q2244 AND symb_decoder(16#a1#)) OR
 					(reg_q2244 AND symb_decoder(16#d5#)) OR
 					(reg_q2244 AND symb_decoder(16#7b#)) OR
 					(reg_q2244 AND symb_decoder(16#97#)) OR
 					(reg_q2244 AND symb_decoder(16#20#)) OR
 					(reg_q2244 AND symb_decoder(16#63#)) OR
 					(reg_q2244 AND symb_decoder(16#f0#)) OR
 					(reg_q2244 AND symb_decoder(16#f9#)) OR
 					(reg_q2244 AND symb_decoder(16#98#)) OR
 					(reg_q2244 AND symb_decoder(16#df#)) OR
 					(reg_q2244 AND symb_decoder(16#b8#)) OR
 					(reg_q2244 AND symb_decoder(16#74#)) OR
 					(reg_q2244 AND symb_decoder(16#96#)) OR
 					(reg_q2244 AND symb_decoder(16#68#)) OR
 					(reg_q2244 AND symb_decoder(16#b7#)) OR
 					(reg_q2244 AND symb_decoder(16#46#)) OR
 					(reg_q2244 AND symb_decoder(16#3a#)) OR
 					(reg_q2244 AND symb_decoder(16#f3#)) OR
 					(reg_q2244 AND symb_decoder(16#2f#)) OR
 					(reg_q2244 AND symb_decoder(16#26#)) OR
 					(reg_q2244 AND symb_decoder(16#dc#)) OR
 					(reg_q2244 AND symb_decoder(16#55#)) OR
 					(reg_q2244 AND symb_decoder(16#cf#)) OR
 					(reg_q2244 AND symb_decoder(16#77#)) OR
 					(reg_q2244 AND symb_decoder(16#b0#)) OR
 					(reg_q2244 AND symb_decoder(16#db#)) OR
 					(reg_q2244 AND symb_decoder(16#58#)) OR
 					(reg_q2244 AND symb_decoder(16#44#)) OR
 					(reg_q2244 AND symb_decoder(16#3d#)) OR
 					(reg_q2244 AND symb_decoder(16#80#)) OR
 					(reg_q2244 AND symb_decoder(16#04#)) OR
 					(reg_q2244 AND symb_decoder(16#d7#)) OR
 					(reg_q2244 AND symb_decoder(16#b1#)) OR
 					(reg_q2244 AND symb_decoder(16#5e#)) OR
 					(reg_q2244 AND symb_decoder(16#72#)) OR
 					(reg_q2244 AND symb_decoder(16#52#)) OR
 					(reg_q2244 AND symb_decoder(16#73#)) OR
 					(reg_q2244 AND symb_decoder(16#d4#)) OR
 					(reg_q2244 AND symb_decoder(16#b4#)) OR
 					(reg_q2244 AND symb_decoder(16#5d#)) OR
 					(reg_q2244 AND symb_decoder(16#1b#)) OR
 					(reg_q2244 AND symb_decoder(16#32#)) OR
 					(reg_q2244 AND symb_decoder(16#21#)) OR
 					(reg_q2244 AND symb_decoder(16#90#)) OR
 					(reg_q2244 AND symb_decoder(16#6a#)) OR
 					(reg_q2244 AND symb_decoder(16#ee#)) OR
 					(reg_q2244 AND symb_decoder(16#b3#)) OR
 					(reg_q2244 AND symb_decoder(16#3e#)) OR
 					(reg_q2244 AND symb_decoder(16#9d#)) OR
 					(reg_q2244 AND symb_decoder(16#8b#)) OR
 					(reg_q2244 AND symb_decoder(16#62#)) OR
 					(reg_q2244 AND symb_decoder(16#bd#)) OR
 					(reg_q2244 AND symb_decoder(16#b9#)) OR
 					(reg_q2244 AND symb_decoder(16#5f#)) OR
 					(reg_q2244 AND symb_decoder(16#12#)) OR
 					(reg_q2244 AND symb_decoder(16#ea#)) OR
 					(reg_q2244 AND symb_decoder(16#e2#)) OR
 					(reg_q2244 AND symb_decoder(16#57#)) OR
 					(reg_q2244 AND symb_decoder(16#66#)) OR
 					(reg_q2244 AND symb_decoder(16#ec#)) OR
 					(reg_q2244 AND symb_decoder(16#fb#)) OR
 					(reg_q2244 AND symb_decoder(16#67#)) OR
 					(reg_q2244 AND symb_decoder(16#19#)) OR
 					(reg_q2244 AND symb_decoder(16#86#)) OR
 					(reg_q2244 AND symb_decoder(16#56#)) OR
 					(reg_q2244 AND symb_decoder(16#5b#)) OR
 					(reg_q2244 AND symb_decoder(16#69#)) OR
 					(reg_q2244 AND symb_decoder(16#ef#)) OR
 					(reg_q2244 AND symb_decoder(16#4a#)) OR
 					(reg_q2244 AND symb_decoder(16#da#)) OR
 					(reg_q2244 AND symb_decoder(16#e6#)) OR
 					(reg_q2244 AND symb_decoder(16#43#)) OR
 					(reg_q2244 AND symb_decoder(16#51#)) OR
 					(reg_q2244 AND symb_decoder(16#ce#)) OR
 					(reg_q2244 AND symb_decoder(16#fc#)) OR
 					(reg_q2244 AND symb_decoder(16#81#)) OR
 					(reg_q2244 AND symb_decoder(16#82#)) OR
 					(reg_q2244 AND symb_decoder(16#88#)) OR
 					(reg_q2244 AND symb_decoder(16#de#)) OR
 					(reg_q2244 AND symb_decoder(16#8d#)) OR
 					(reg_q2244 AND symb_decoder(16#9c#)) OR
 					(reg_q2244 AND symb_decoder(16#41#)) OR
 					(reg_q2244 AND symb_decoder(16#d9#)) OR
 					(reg_q2244 AND symb_decoder(16#45#)) OR
 					(reg_q2244 AND symb_decoder(16#cc#)) OR
 					(reg_q2244 AND symb_decoder(16#c3#)) OR
 					(reg_q2244 AND symb_decoder(16#7a#)) OR
 					(reg_q2244 AND symb_decoder(16#d0#)) OR
 					(reg_q2244 AND symb_decoder(16#39#)) OR
 					(reg_q2244 AND symb_decoder(16#09#)) OR
 					(reg_q2244 AND symb_decoder(16#a9#)) OR
 					(reg_q2244 AND symb_decoder(16#2e#)) OR
 					(reg_q2244 AND symb_decoder(16#87#)) OR
 					(reg_q2244 AND symb_decoder(16#01#)) OR
 					(reg_q2244 AND symb_decoder(16#4e#)) OR
 					(reg_q2244 AND symb_decoder(16#9b#)) OR
 					(reg_q2244 AND symb_decoder(16#d8#)) OR
 					(reg_q2244 AND symb_decoder(16#22#)) OR
 					(reg_q2244 AND symb_decoder(16#91#)) OR
 					(reg_q2244 AND symb_decoder(16#42#)) OR
 					(reg_q2244 AND symb_decoder(16#a5#)) OR
 					(reg_q2244 AND symb_decoder(16#64#)) OR
 					(reg_q2244 AND symb_decoder(16#1a#)) OR
 					(reg_q2244 AND symb_decoder(16#92#)) OR
 					(reg_q2244 AND symb_decoder(16#e8#)) OR
 					(reg_q2244 AND symb_decoder(16#25#)) OR
 					(reg_q2244 AND symb_decoder(16#e3#)) OR
 					(reg_q2244 AND symb_decoder(16#9e#)) OR
 					(reg_q2244 AND symb_decoder(16#a0#)) OR
 					(reg_q2244 AND symb_decoder(16#4f#)) OR
 					(reg_q2244 AND symb_decoder(16#5c#));
reg_q2244_init <= '0' ;
	p_reg_q2244: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2244 <= reg_q2244_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2244 <= reg_q2244_init;
        else
          reg_q2244 <= reg_q2244_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph15

reg_q1682_in <= (reg_q1672 AND symb_decoder(16#a9#)) OR
 					(reg_q1672 AND symb_decoder(16#66#)) OR
 					(reg_q1672 AND symb_decoder(16#ae#)) OR
 					(reg_q1672 AND symb_decoder(16#69#)) OR
 					(reg_q1672 AND symb_decoder(16#71#)) OR
 					(reg_q1672 AND symb_decoder(16#d3#)) OR
 					(reg_q1672 AND symb_decoder(16#a0#)) OR
 					(reg_q1672 AND symb_decoder(16#91#)) OR
 					(reg_q1672 AND symb_decoder(16#a3#)) OR
 					(reg_q1672 AND symb_decoder(16#d4#)) OR
 					(reg_q1672 AND symb_decoder(16#da#)) OR
 					(reg_q1672 AND symb_decoder(16#8d#)) OR
 					(reg_q1672 AND symb_decoder(16#a5#)) OR
 					(reg_q1672 AND symb_decoder(16#72#)) OR
 					(reg_q1672 AND symb_decoder(16#1d#)) OR
 					(reg_q1672 AND symb_decoder(16#ce#)) OR
 					(reg_q1672 AND symb_decoder(16#20#)) OR
 					(reg_q1672 AND symb_decoder(16#2b#)) OR
 					(reg_q1672 AND symb_decoder(16#35#)) OR
 					(reg_q1672 AND symb_decoder(16#aa#)) OR
 					(reg_q1672 AND symb_decoder(16#32#)) OR
 					(reg_q1672 AND symb_decoder(16#e0#)) OR
 					(reg_q1672 AND symb_decoder(16#eb#)) OR
 					(reg_q1672 AND symb_decoder(16#9c#)) OR
 					(reg_q1672 AND symb_decoder(16#b6#)) OR
 					(reg_q1672 AND symb_decoder(16#53#)) OR
 					(reg_q1672 AND symb_decoder(16#39#)) OR
 					(reg_q1672 AND symb_decoder(16#b5#)) OR
 					(reg_q1672 AND symb_decoder(16#67#)) OR
 					(reg_q1672 AND symb_decoder(16#05#)) OR
 					(reg_q1672 AND symb_decoder(16#42#)) OR
 					(reg_q1672 AND symb_decoder(16#c8#)) OR
 					(reg_q1672 AND symb_decoder(16#b9#)) OR
 					(reg_q1672 AND symb_decoder(16#0f#)) OR
 					(reg_q1672 AND symb_decoder(16#19#)) OR
 					(reg_q1672 AND symb_decoder(16#95#)) OR
 					(reg_q1672 AND symb_decoder(16#5f#)) OR
 					(reg_q1672 AND symb_decoder(16#af#)) OR
 					(reg_q1672 AND symb_decoder(16#3b#)) OR
 					(reg_q1672 AND symb_decoder(16#ba#)) OR
 					(reg_q1672 AND symb_decoder(16#76#)) OR
 					(reg_q1672 AND symb_decoder(16#d9#)) OR
 					(reg_q1672 AND symb_decoder(16#fb#)) OR
 					(reg_q1672 AND symb_decoder(16#96#)) OR
 					(reg_q1672 AND symb_decoder(16#93#)) OR
 					(reg_q1672 AND symb_decoder(16#f3#)) OR
 					(reg_q1672 AND symb_decoder(16#bb#)) OR
 					(reg_q1672 AND symb_decoder(16#5c#)) OR
 					(reg_q1672 AND symb_decoder(16#6c#)) OR
 					(reg_q1672 AND symb_decoder(16#cc#)) OR
 					(reg_q1672 AND symb_decoder(16#56#)) OR
 					(reg_q1672 AND symb_decoder(16#f0#)) OR
 					(reg_q1672 AND symb_decoder(16#50#)) OR
 					(reg_q1672 AND symb_decoder(16#bf#)) OR
 					(reg_q1672 AND symb_decoder(16#41#)) OR
 					(reg_q1672 AND symb_decoder(16#8e#)) OR
 					(reg_q1672 AND symb_decoder(16#14#)) OR
 					(reg_q1672 AND symb_decoder(16#79#)) OR
 					(reg_q1672 AND symb_decoder(16#00#)) OR
 					(reg_q1672 AND symb_decoder(16#44#)) OR
 					(reg_q1672 AND symb_decoder(16#37#)) OR
 					(reg_q1672 AND symb_decoder(16#43#)) OR
 					(reg_q1672 AND symb_decoder(16#b0#)) OR
 					(reg_q1672 AND symb_decoder(16#c2#)) OR
 					(reg_q1672 AND symb_decoder(16#ef#)) OR
 					(reg_q1672 AND symb_decoder(16#12#)) OR
 					(reg_q1672 AND symb_decoder(16#52#)) OR
 					(reg_q1672 AND symb_decoder(16#01#)) OR
 					(reg_q1672 AND symb_decoder(16#ca#)) OR
 					(reg_q1672 AND symb_decoder(16#a7#)) OR
 					(reg_q1672 AND symb_decoder(16#ee#)) OR
 					(reg_q1672 AND symb_decoder(16#09#)) OR
 					(reg_q1672 AND symb_decoder(16#89#)) OR
 					(reg_q1672 AND symb_decoder(16#fa#)) OR
 					(reg_q1672 AND symb_decoder(16#c4#)) OR
 					(reg_q1672 AND symb_decoder(16#03#)) OR
 					(reg_q1672 AND symb_decoder(16#80#)) OR
 					(reg_q1672 AND symb_decoder(16#fc#)) OR
 					(reg_q1672 AND symb_decoder(16#8b#)) OR
 					(reg_q1672 AND symb_decoder(16#27#)) OR
 					(reg_q1672 AND symb_decoder(16#9b#)) OR
 					(reg_q1672 AND symb_decoder(16#23#)) OR
 					(reg_q1672 AND symb_decoder(16#e8#)) OR
 					(reg_q1672 AND symb_decoder(16#2e#)) OR
 					(reg_q1672 AND symb_decoder(16#f7#)) OR
 					(reg_q1672 AND symb_decoder(16#7c#)) OR
 					(reg_q1672 AND symb_decoder(16#9a#)) OR
 					(reg_q1672 AND symb_decoder(16#cf#)) OR
 					(reg_q1672 AND symb_decoder(16#22#)) OR
 					(reg_q1672 AND symb_decoder(16#d2#)) OR
 					(reg_q1672 AND symb_decoder(16#9e#)) OR
 					(reg_q1672 AND symb_decoder(16#e7#)) OR
 					(reg_q1672 AND symb_decoder(16#d8#)) OR
 					(reg_q1672 AND symb_decoder(16#6d#)) OR
 					(reg_q1672 AND symb_decoder(16#6f#)) OR
 					(reg_q1672 AND symb_decoder(16#f4#)) OR
 					(reg_q1672 AND symb_decoder(16#33#)) OR
 					(reg_q1672 AND symb_decoder(16#8f#)) OR
 					(reg_q1672 AND symb_decoder(16#51#)) OR
 					(reg_q1672 AND symb_decoder(16#d1#)) OR
 					(reg_q1672 AND symb_decoder(16#99#)) OR
 					(reg_q1672 AND symb_decoder(16#ec#)) OR
 					(reg_q1672 AND symb_decoder(16#c7#)) OR
 					(reg_q1672 AND symb_decoder(16#55#)) OR
 					(reg_q1672 AND symb_decoder(16#ac#)) OR
 					(reg_q1672 AND symb_decoder(16#a1#)) OR
 					(reg_q1672 AND symb_decoder(16#dd#)) OR
 					(reg_q1672 AND symb_decoder(16#5b#)) OR
 					(reg_q1672 AND symb_decoder(16#06#)) OR
 					(reg_q1672 AND symb_decoder(16#c1#)) OR
 					(reg_q1672 AND symb_decoder(16#74#)) OR
 					(reg_q1672 AND symb_decoder(16#a2#)) OR
 					(reg_q1672 AND symb_decoder(16#21#)) OR
 					(reg_q1672 AND symb_decoder(16#f5#)) OR
 					(reg_q1672 AND symb_decoder(16#92#)) OR
 					(reg_q1672 AND symb_decoder(16#73#)) OR
 					(reg_q1672 AND symb_decoder(16#86#)) OR
 					(reg_q1672 AND symb_decoder(16#d0#)) OR
 					(reg_q1672 AND symb_decoder(16#cd#)) OR
 					(reg_q1672 AND symb_decoder(16#81#)) OR
 					(reg_q1672 AND symb_decoder(16#04#)) OR
 					(reg_q1672 AND symb_decoder(16#8c#)) OR
 					(reg_q1672 AND symb_decoder(16#2f#)) OR
 					(reg_q1672 AND symb_decoder(16#c0#)) OR
 					(reg_q1672 AND symb_decoder(16#7d#)) OR
 					(reg_q1672 AND symb_decoder(16#2a#)) OR
 					(reg_q1672 AND symb_decoder(16#4e#)) OR
 					(reg_q1672 AND symb_decoder(16#45#)) OR
 					(reg_q1672 AND symb_decoder(16#1a#)) OR
 					(reg_q1672 AND symb_decoder(16#84#)) OR
 					(reg_q1672 AND symb_decoder(16#59#)) OR
 					(reg_q1672 AND symb_decoder(16#a6#)) OR
 					(reg_q1672 AND symb_decoder(16#11#)) OR
 					(reg_q1672 AND symb_decoder(16#7a#)) OR
 					(reg_q1672 AND symb_decoder(16#1c#)) OR
 					(reg_q1672 AND symb_decoder(16#64#)) OR
 					(reg_q1672 AND symb_decoder(16#61#)) OR
 					(reg_q1672 AND symb_decoder(16#b8#)) OR
 					(reg_q1672 AND symb_decoder(16#6b#)) OR
 					(reg_q1672 AND symb_decoder(16#db#)) OR
 					(reg_q1672 AND symb_decoder(16#5d#)) OR
 					(reg_q1672 AND symb_decoder(16#77#)) OR
 					(reg_q1672 AND symb_decoder(16#c3#)) OR
 					(reg_q1672 AND symb_decoder(16#0c#)) OR
 					(reg_q1672 AND symb_decoder(16#85#)) OR
 					(reg_q1672 AND symb_decoder(16#8a#)) OR
 					(reg_q1672 AND symb_decoder(16#6e#)) OR
 					(reg_q1672 AND symb_decoder(16#57#)) OR
 					(reg_q1672 AND symb_decoder(16#4f#)) OR
 					(reg_q1672 AND symb_decoder(16#ea#)) OR
 					(reg_q1672 AND symb_decoder(16#bd#)) OR
 					(reg_q1672 AND symb_decoder(16#5a#)) OR
 					(reg_q1672 AND symb_decoder(16#68#)) OR
 					(reg_q1672 AND symb_decoder(16#65#)) OR
 					(reg_q1672 AND symb_decoder(16#17#)) OR
 					(reg_q1672 AND symb_decoder(16#4a#)) OR
 					(reg_q1672 AND symb_decoder(16#88#)) OR
 					(reg_q1672 AND symb_decoder(16#d5#)) OR
 					(reg_q1672 AND symb_decoder(16#f1#)) OR
 					(reg_q1672 AND symb_decoder(16#b4#)) OR
 					(reg_q1672 AND symb_decoder(16#3d#)) OR
 					(reg_q1672 AND symb_decoder(16#4d#)) OR
 					(reg_q1672 AND symb_decoder(16#fd#)) OR
 					(reg_q1672 AND symb_decoder(16#3f#)) OR
 					(reg_q1672 AND symb_decoder(16#f8#)) OR
 					(reg_q1672 AND symb_decoder(16#e9#)) OR
 					(reg_q1672 AND symb_decoder(16#38#)) OR
 					(reg_q1672 AND symb_decoder(16#83#)) OR
 					(reg_q1672 AND symb_decoder(16#9f#)) OR
 					(reg_q1672 AND symb_decoder(16#15#)) OR
 					(reg_q1672 AND symb_decoder(16#f6#)) OR
 					(reg_q1672 AND symb_decoder(16#0b#)) OR
 					(reg_q1672 AND symb_decoder(16#16#)) OR
 					(reg_q1672 AND symb_decoder(16#75#)) OR
 					(reg_q1672 AND symb_decoder(16#24#)) OR
 					(reg_q1672 AND symb_decoder(16#62#)) OR
 					(reg_q1672 AND symb_decoder(16#58#)) OR
 					(reg_q1672 AND symb_decoder(16#7f#)) OR
 					(reg_q1672 AND symb_decoder(16#be#)) OR
 					(reg_q1672 AND symb_decoder(16#90#)) OR
 					(reg_q1672 AND symb_decoder(16#10#)) OR
 					(reg_q1672 AND symb_decoder(16#48#)) OR
 					(reg_q1672 AND symb_decoder(16#e1#)) OR
 					(reg_q1672 AND symb_decoder(16#08#)) OR
 					(reg_q1672 AND symb_decoder(16#d6#)) OR
 					(reg_q1672 AND symb_decoder(16#07#)) OR
 					(reg_q1672 AND symb_decoder(16#bc#)) OR
 					(reg_q1672 AND symb_decoder(16#26#)) OR
 					(reg_q1672 AND symb_decoder(16#63#)) OR
 					(reg_q1672 AND symb_decoder(16#0e#)) OR
 					(reg_q1672 AND symb_decoder(16#e5#)) OR
 					(reg_q1672 AND symb_decoder(16#28#)) OR
 					(reg_q1672 AND symb_decoder(16#13#)) OR
 					(reg_q1672 AND symb_decoder(16#1f#)) OR
 					(reg_q1672 AND symb_decoder(16#cb#)) OR
 					(reg_q1672 AND symb_decoder(16#1e#)) OR
 					(reg_q1672 AND symb_decoder(16#1b#)) OR
 					(reg_q1672 AND symb_decoder(16#7e#)) OR
 					(reg_q1672 AND symb_decoder(16#4b#)) OR
 					(reg_q1672 AND symb_decoder(16#31#)) OR
 					(reg_q1672 AND symb_decoder(16#60#)) OR
 					(reg_q1672 AND symb_decoder(16#30#)) OR
 					(reg_q1672 AND symb_decoder(16#4c#)) OR
 					(reg_q1672 AND symb_decoder(16#18#)) OR
 					(reg_q1672 AND symb_decoder(16#36#)) OR
 					(reg_q1672 AND symb_decoder(16#c5#)) OR
 					(reg_q1672 AND symb_decoder(16#9d#)) OR
 					(reg_q1672 AND symb_decoder(16#47#)) OR
 					(reg_q1672 AND symb_decoder(16#fe#)) OR
 					(reg_q1672 AND symb_decoder(16#3a#)) OR
 					(reg_q1672 AND symb_decoder(16#d7#)) OR
 					(reg_q1672 AND symb_decoder(16#2c#)) OR
 					(reg_q1672 AND symb_decoder(16#49#)) OR
 					(reg_q1672 AND symb_decoder(16#7b#)) OR
 					(reg_q1672 AND symb_decoder(16#ad#)) OR
 					(reg_q1672 AND symb_decoder(16#54#)) OR
 					(reg_q1672 AND symb_decoder(16#b2#)) OR
 					(reg_q1672 AND symb_decoder(16#3e#)) OR
 					(reg_q1672 AND symb_decoder(16#70#)) OR
 					(reg_q1672 AND symb_decoder(16#b1#)) OR
 					(reg_q1672 AND symb_decoder(16#6a#)) OR
 					(reg_q1672 AND symb_decoder(16#f2#)) OR
 					(reg_q1672 AND symb_decoder(16#3c#)) OR
 					(reg_q1672 AND symb_decoder(16#ed#)) OR
 					(reg_q1672 AND symb_decoder(16#40#)) OR
 					(reg_q1672 AND symb_decoder(16#e4#)) OR
 					(reg_q1672 AND symb_decoder(16#dc#)) OR
 					(reg_q1672 AND symb_decoder(16#34#)) OR
 					(reg_q1672 AND symb_decoder(16#e3#)) OR
 					(reg_q1672 AND symb_decoder(16#2d#)) OR
 					(reg_q1672 AND symb_decoder(16#f9#)) OR
 					(reg_q1672 AND symb_decoder(16#5e#)) OR
 					(reg_q1672 AND symb_decoder(16#29#)) OR
 					(reg_q1672 AND symb_decoder(16#ab#)) OR
 					(reg_q1672 AND symb_decoder(16#02#)) OR
 					(reg_q1672 AND symb_decoder(16#e2#)) OR
 					(reg_q1672 AND symb_decoder(16#97#)) OR
 					(reg_q1672 AND symb_decoder(16#c9#)) OR
 					(reg_q1672 AND symb_decoder(16#a4#)) OR
 					(reg_q1672 AND symb_decoder(16#ff#)) OR
 					(reg_q1672 AND symb_decoder(16#de#)) OR
 					(reg_q1672 AND symb_decoder(16#82#)) OR
 					(reg_q1672 AND symb_decoder(16#c6#)) OR
 					(reg_q1672 AND symb_decoder(16#25#)) OR
 					(reg_q1672 AND symb_decoder(16#98#)) OR
 					(reg_q1672 AND symb_decoder(16#78#)) OR
 					(reg_q1672 AND symb_decoder(16#df#)) OR
 					(reg_q1672 AND symb_decoder(16#46#)) OR
 					(reg_q1672 AND symb_decoder(16#b7#)) OR
 					(reg_q1672 AND symb_decoder(16#b3#)) OR
 					(reg_q1672 AND symb_decoder(16#e6#)) OR
 					(reg_q1672 AND symb_decoder(16#87#)) OR
 					(reg_q1672 AND symb_decoder(16#94#)) OR
 					(reg_q1672 AND symb_decoder(16#a8#)) OR
 					(reg_q1682 AND symb_decoder(16#30#)) OR
 					(reg_q1682 AND symb_decoder(16#6e#)) OR
 					(reg_q1682 AND symb_decoder(16#1b#)) OR
 					(reg_q1682 AND symb_decoder(16#68#)) OR
 					(reg_q1682 AND symb_decoder(16#97#)) OR
 					(reg_q1682 AND symb_decoder(16#13#)) OR
 					(reg_q1682 AND symb_decoder(16#c6#)) OR
 					(reg_q1682 AND symb_decoder(16#62#)) OR
 					(reg_q1682 AND symb_decoder(16#d9#)) OR
 					(reg_q1682 AND symb_decoder(16#0e#)) OR
 					(reg_q1682 AND symb_decoder(16#81#)) OR
 					(reg_q1682 AND symb_decoder(16#a6#)) OR
 					(reg_q1682 AND symb_decoder(16#fc#)) OR
 					(reg_q1682 AND symb_decoder(16#de#)) OR
 					(reg_q1682 AND symb_decoder(16#0b#)) OR
 					(reg_q1682 AND symb_decoder(16#29#)) OR
 					(reg_q1682 AND symb_decoder(16#cb#)) OR
 					(reg_q1682 AND symb_decoder(16#e8#)) OR
 					(reg_q1682 AND symb_decoder(16#24#)) OR
 					(reg_q1682 AND symb_decoder(16#46#)) OR
 					(reg_q1682 AND symb_decoder(16#18#)) OR
 					(reg_q1682 AND symb_decoder(16#83#)) OR
 					(reg_q1682 AND symb_decoder(16#a5#)) OR
 					(reg_q1682 AND symb_decoder(16#45#)) OR
 					(reg_q1682 AND symb_decoder(16#5e#)) OR
 					(reg_q1682 AND symb_decoder(16#41#)) OR
 					(reg_q1682 AND symb_decoder(16#ff#)) OR
 					(reg_q1682 AND symb_decoder(16#bb#)) OR
 					(reg_q1682 AND symb_decoder(16#99#)) OR
 					(reg_q1682 AND symb_decoder(16#6a#)) OR
 					(reg_q1682 AND symb_decoder(16#7c#)) OR
 					(reg_q1682 AND symb_decoder(16#3c#)) OR
 					(reg_q1682 AND symb_decoder(16#da#)) OR
 					(reg_q1682 AND symb_decoder(16#79#)) OR
 					(reg_q1682 AND symb_decoder(16#71#)) OR
 					(reg_q1682 AND symb_decoder(16#4d#)) OR
 					(reg_q1682 AND symb_decoder(16#f1#)) OR
 					(reg_q1682 AND symb_decoder(16#9a#)) OR
 					(reg_q1682 AND symb_decoder(16#a2#)) OR
 					(reg_q1682 AND symb_decoder(16#54#)) OR
 					(reg_q1682 AND symb_decoder(16#36#)) OR
 					(reg_q1682 AND symb_decoder(16#57#)) OR
 					(reg_q1682 AND symb_decoder(16#21#)) OR
 					(reg_q1682 AND symb_decoder(16#1d#)) OR
 					(reg_q1682 AND symb_decoder(16#a9#)) OR
 					(reg_q1682 AND symb_decoder(16#0c#)) OR
 					(reg_q1682 AND symb_decoder(16#7a#)) OR
 					(reg_q1682 AND symb_decoder(16#c7#)) OR
 					(reg_q1682 AND symb_decoder(16#26#)) OR
 					(reg_q1682 AND symb_decoder(16#f3#)) OR
 					(reg_q1682 AND symb_decoder(16#02#)) OR
 					(reg_q1682 AND symb_decoder(16#a7#)) OR
 					(reg_q1682 AND symb_decoder(16#af#)) OR
 					(reg_q1682 AND symb_decoder(16#69#)) OR
 					(reg_q1682 AND symb_decoder(16#85#)) OR
 					(reg_q1682 AND symb_decoder(16#a0#)) OR
 					(reg_q1682 AND symb_decoder(16#c0#)) OR
 					(reg_q1682 AND symb_decoder(16#e4#)) OR
 					(reg_q1682 AND symb_decoder(16#01#)) OR
 					(reg_q1682 AND symb_decoder(16#f8#)) OR
 					(reg_q1682 AND symb_decoder(16#05#)) OR
 					(reg_q1682 AND symb_decoder(16#48#)) OR
 					(reg_q1682 AND symb_decoder(16#7f#)) OR
 					(reg_q1682 AND symb_decoder(16#9d#)) OR
 					(reg_q1682 AND symb_decoder(16#df#)) OR
 					(reg_q1682 AND symb_decoder(16#8b#)) OR
 					(reg_q1682 AND symb_decoder(16#53#)) OR
 					(reg_q1682 AND symb_decoder(16#e0#)) OR
 					(reg_q1682 AND symb_decoder(16#f0#)) OR
 					(reg_q1682 AND symb_decoder(16#b5#)) OR
 					(reg_q1682 AND symb_decoder(16#04#)) OR
 					(reg_q1682 AND symb_decoder(16#10#)) OR
 					(reg_q1682 AND symb_decoder(16#c8#)) OR
 					(reg_q1682 AND symb_decoder(16#08#)) OR
 					(reg_q1682 AND symb_decoder(16#4c#)) OR
 					(reg_q1682 AND symb_decoder(16#a1#)) OR
 					(reg_q1682 AND symb_decoder(16#d2#)) OR
 					(reg_q1682 AND symb_decoder(16#5b#)) OR
 					(reg_q1682 AND symb_decoder(16#c9#)) OR
 					(reg_q1682 AND symb_decoder(16#1a#)) OR
 					(reg_q1682 AND symb_decoder(16#d4#)) OR
 					(reg_q1682 AND symb_decoder(16#db#)) OR
 					(reg_q1682 AND symb_decoder(16#e5#)) OR
 					(reg_q1682 AND symb_decoder(16#06#)) OR
 					(reg_q1682 AND symb_decoder(16#16#)) OR
 					(reg_q1682 AND symb_decoder(16#dd#)) OR
 					(reg_q1682 AND symb_decoder(16#7b#)) OR
 					(reg_q1682 AND symb_decoder(16#4b#)) OR
 					(reg_q1682 AND symb_decoder(16#76#)) OR
 					(reg_q1682 AND symb_decoder(16#f7#)) OR
 					(reg_q1682 AND symb_decoder(16#fb#)) OR
 					(reg_q1682 AND symb_decoder(16#17#)) OR
 					(reg_q1682 AND symb_decoder(16#34#)) OR
 					(reg_q1682 AND symb_decoder(16#cd#)) OR
 					(reg_q1682 AND symb_decoder(16#3e#)) OR
 					(reg_q1682 AND symb_decoder(16#c2#)) OR
 					(reg_q1682 AND symb_decoder(16#ac#)) OR
 					(reg_q1682 AND symb_decoder(16#fd#)) OR
 					(reg_q1682 AND symb_decoder(16#ae#)) OR
 					(reg_q1682 AND symb_decoder(16#2e#)) OR
 					(reg_q1682 AND symb_decoder(16#5f#)) OR
 					(reg_q1682 AND symb_decoder(16#1c#)) OR
 					(reg_q1682 AND symb_decoder(16#66#)) OR
 					(reg_q1682 AND symb_decoder(16#cc#)) OR
 					(reg_q1682 AND symb_decoder(16#d6#)) OR
 					(reg_q1682 AND symb_decoder(16#38#)) OR
 					(reg_q1682 AND symb_decoder(16#bf#)) OR
 					(reg_q1682 AND symb_decoder(16#e9#)) OR
 					(reg_q1682 AND symb_decoder(16#72#)) OR
 					(reg_q1682 AND symb_decoder(16#ef#)) OR
 					(reg_q1682 AND symb_decoder(16#9c#)) OR
 					(reg_q1682 AND symb_decoder(16#8e#)) OR
 					(reg_q1682 AND symb_decoder(16#93#)) OR
 					(reg_q1682 AND symb_decoder(16#6f#)) OR
 					(reg_q1682 AND symb_decoder(16#90#)) OR
 					(reg_q1682 AND symb_decoder(16#52#)) OR
 					(reg_q1682 AND symb_decoder(16#22#)) OR
 					(reg_q1682 AND symb_decoder(16#25#)) OR
 					(reg_q1682 AND symb_decoder(16#07#)) OR
 					(reg_q1682 AND symb_decoder(16#c3#)) OR
 					(reg_q1682 AND symb_decoder(16#00#)) OR
 					(reg_q1682 AND symb_decoder(16#fe#)) OR
 					(reg_q1682 AND symb_decoder(16#2f#)) OR
 					(reg_q1682 AND symb_decoder(16#73#)) OR
 					(reg_q1682 AND symb_decoder(16#95#)) OR
 					(reg_q1682 AND symb_decoder(16#4a#)) OR
 					(reg_q1682 AND symb_decoder(16#51#)) OR
 					(reg_q1682 AND symb_decoder(16#42#)) OR
 					(reg_q1682 AND symb_decoder(16#6d#)) OR
 					(reg_q1682 AND symb_decoder(16#1f#)) OR
 					(reg_q1682 AND symb_decoder(16#ab#)) OR
 					(reg_q1682 AND symb_decoder(16#67#)) OR
 					(reg_q1682 AND symb_decoder(16#43#)) OR
 					(reg_q1682 AND symb_decoder(16#87#)) OR
 					(reg_q1682 AND symb_decoder(16#b6#)) OR
 					(reg_q1682 AND symb_decoder(16#2a#)) OR
 					(reg_q1682 AND symb_decoder(16#ed#)) OR
 					(reg_q1682 AND symb_decoder(16#58#)) OR
 					(reg_q1682 AND symb_decoder(16#84#)) OR
 					(reg_q1682 AND symb_decoder(16#f5#)) OR
 					(reg_q1682 AND symb_decoder(16#e6#)) OR
 					(reg_q1682 AND symb_decoder(16#50#)) OR
 					(reg_q1682 AND symb_decoder(16#4f#)) OR
 					(reg_q1682 AND symb_decoder(16#e2#)) OR
 					(reg_q1682 AND symb_decoder(16#d1#)) OR
 					(reg_q1682 AND symb_decoder(16#7e#)) OR
 					(reg_q1682 AND symb_decoder(16#5d#)) OR
 					(reg_q1682 AND symb_decoder(16#f6#)) OR
 					(reg_q1682 AND symb_decoder(16#37#)) OR
 					(reg_q1682 AND symb_decoder(16#d0#)) OR
 					(reg_q1682 AND symb_decoder(16#ba#)) OR
 					(reg_q1682 AND symb_decoder(16#7d#)) OR
 					(reg_q1682 AND symb_decoder(16#09#)) OR
 					(reg_q1682 AND symb_decoder(16#49#)) OR
 					(reg_q1682 AND symb_decoder(16#3d#)) OR
 					(reg_q1682 AND symb_decoder(16#d8#)) OR
 					(reg_q1682 AND symb_decoder(16#ce#)) OR
 					(reg_q1682 AND symb_decoder(16#80#)) OR
 					(reg_q1682 AND symb_decoder(16#11#)) OR
 					(reg_q1682 AND symb_decoder(16#a8#)) OR
 					(reg_q1682 AND symb_decoder(16#bd#)) OR
 					(reg_q1682 AND symb_decoder(16#cf#)) OR
 					(reg_q1682 AND symb_decoder(16#91#)) OR
 					(reg_q1682 AND symb_decoder(16#03#)) OR
 					(reg_q1682 AND symb_decoder(16#98#)) OR
 					(reg_q1682 AND symb_decoder(16#14#)) OR
 					(reg_q1682 AND symb_decoder(16#a4#)) OR
 					(reg_q1682 AND symb_decoder(16#b7#)) OR
 					(reg_q1682 AND symb_decoder(16#ea#)) OR
 					(reg_q1682 AND symb_decoder(16#e3#)) OR
 					(reg_q1682 AND symb_decoder(16#d5#)) OR
 					(reg_q1682 AND symb_decoder(16#f4#)) OR
 					(reg_q1682 AND symb_decoder(16#c4#)) OR
 					(reg_q1682 AND symb_decoder(16#b9#)) OR
 					(reg_q1682 AND symb_decoder(16#3a#)) OR
 					(reg_q1682 AND symb_decoder(16#96#)) OR
 					(reg_q1682 AND symb_decoder(16#40#)) OR
 					(reg_q1682 AND symb_decoder(16#20#)) OR
 					(reg_q1682 AND symb_decoder(16#55#)) OR
 					(reg_q1682 AND symb_decoder(16#28#)) OR
 					(reg_q1682 AND symb_decoder(16#b1#)) OR
 					(reg_q1682 AND symb_decoder(16#b2#)) OR
 					(reg_q1682 AND symb_decoder(16#6b#)) OR
 					(reg_q1682 AND symb_decoder(16#59#)) OR
 					(reg_q1682 AND symb_decoder(16#39#)) OR
 					(reg_q1682 AND symb_decoder(16#35#)) OR
 					(reg_q1682 AND symb_decoder(16#47#)) OR
 					(reg_q1682 AND symb_decoder(16#33#)) OR
 					(reg_q1682 AND symb_decoder(16#aa#)) OR
 					(reg_q1682 AND symb_decoder(16#9f#)) OR
 					(reg_q1682 AND symb_decoder(16#9b#)) OR
 					(reg_q1682 AND symb_decoder(16#3b#)) OR
 					(reg_q1682 AND symb_decoder(16#75#)) OR
 					(reg_q1682 AND symb_decoder(16#3f#)) OR
 					(reg_q1682 AND symb_decoder(16#92#)) OR
 					(reg_q1682 AND symb_decoder(16#be#)) OR
 					(reg_q1682 AND symb_decoder(16#32#)) OR
 					(reg_q1682 AND symb_decoder(16#1e#)) OR
 					(reg_q1682 AND symb_decoder(16#86#)) OR
 					(reg_q1682 AND symb_decoder(16#78#)) OR
 					(reg_q1682 AND symb_decoder(16#a3#)) OR
 					(reg_q1682 AND symb_decoder(16#64#)) OR
 					(reg_q1682 AND symb_decoder(16#b4#)) OR
 					(reg_q1682 AND symb_decoder(16#8f#)) OR
 					(reg_q1682 AND symb_decoder(16#44#)) OR
 					(reg_q1682 AND symb_decoder(16#2b#)) OR
 					(reg_q1682 AND symb_decoder(16#d3#)) OR
 					(reg_q1682 AND symb_decoder(16#eb#)) OR
 					(reg_q1682 AND symb_decoder(16#bc#)) OR
 					(reg_q1682 AND symb_decoder(16#ca#)) OR
 					(reg_q1682 AND symb_decoder(16#f9#)) OR
 					(reg_q1682 AND symb_decoder(16#5c#)) OR
 					(reg_q1682 AND symb_decoder(16#60#)) OR
 					(reg_q1682 AND symb_decoder(16#27#)) OR
 					(reg_q1682 AND symb_decoder(16#89#)) OR
 					(reg_q1682 AND symb_decoder(16#4e#)) OR
 					(reg_q1682 AND symb_decoder(16#23#)) OR
 					(reg_q1682 AND symb_decoder(16#74#)) OR
 					(reg_q1682 AND symb_decoder(16#b8#)) OR
 					(reg_q1682 AND symb_decoder(16#65#)) OR
 					(reg_q1682 AND symb_decoder(16#c1#)) OR
 					(reg_q1682 AND symb_decoder(16#b3#)) OR
 					(reg_q1682 AND symb_decoder(16#ee#)) OR
 					(reg_q1682 AND symb_decoder(16#b0#)) OR
 					(reg_q1682 AND symb_decoder(16#d7#)) OR
 					(reg_q1682 AND symb_decoder(16#12#)) OR
 					(reg_q1682 AND symb_decoder(16#77#)) OR
 					(reg_q1682 AND symb_decoder(16#15#)) OR
 					(reg_q1682 AND symb_decoder(16#9e#)) OR
 					(reg_q1682 AND symb_decoder(16#c5#)) OR
 					(reg_q1682 AND symb_decoder(16#61#)) OR
 					(reg_q1682 AND symb_decoder(16#8c#)) OR
 					(reg_q1682 AND symb_decoder(16#82#)) OR
 					(reg_q1682 AND symb_decoder(16#19#)) OR
 					(reg_q1682 AND symb_decoder(16#dc#)) OR
 					(reg_q1682 AND symb_decoder(16#56#)) OR
 					(reg_q1682 AND symb_decoder(16#ec#)) OR
 					(reg_q1682 AND symb_decoder(16#5a#)) OR
 					(reg_q1682 AND symb_decoder(16#f2#)) OR
 					(reg_q1682 AND symb_decoder(16#2d#)) OR
 					(reg_q1682 AND symb_decoder(16#e1#)) OR
 					(reg_q1682 AND symb_decoder(16#0f#)) OR
 					(reg_q1682 AND symb_decoder(16#8d#)) OR
 					(reg_q1682 AND symb_decoder(16#70#)) OR
 					(reg_q1682 AND symb_decoder(16#88#)) OR
 					(reg_q1682 AND symb_decoder(16#31#)) OR
 					(reg_q1682 AND symb_decoder(16#94#)) OR
 					(reg_q1682 AND symb_decoder(16#ad#)) OR
 					(reg_q1682 AND symb_decoder(16#e7#)) OR
 					(reg_q1682 AND symb_decoder(16#8a#)) OR
 					(reg_q1682 AND symb_decoder(16#63#)) OR
 					(reg_q1682 AND symb_decoder(16#2c#)) OR
 					(reg_q1682 AND symb_decoder(16#fa#)) OR
 					(reg_q1682 AND symb_decoder(16#6c#));
reg_q2625_in <= (reg_q2623 AND symb_decoder(16#42#)) OR
 					(reg_q2623 AND symb_decoder(16#a5#)) OR
 					(reg_q2623 AND symb_decoder(16#f2#)) OR
 					(reg_q2623 AND symb_decoder(16#65#)) OR
 					(reg_q2623 AND symb_decoder(16#e5#)) OR
 					(reg_q2623 AND symb_decoder(16#e1#)) OR
 					(reg_q2623 AND symb_decoder(16#1e#)) OR
 					(reg_q2623 AND symb_decoder(16#3a#)) OR
 					(reg_q2623 AND symb_decoder(16#47#)) OR
 					(reg_q2623 AND symb_decoder(16#4f#)) OR
 					(reg_q2623 AND symb_decoder(16#b0#)) OR
 					(reg_q2623 AND symb_decoder(16#72#)) OR
 					(reg_q2623 AND symb_decoder(16#40#)) OR
 					(reg_q2623 AND symb_decoder(16#15#)) OR
 					(reg_q2623 AND symb_decoder(16#cb#)) OR
 					(reg_q2623 AND symb_decoder(16#1c#)) OR
 					(reg_q2623 AND symb_decoder(16#e2#)) OR
 					(reg_q2623 AND symb_decoder(16#79#)) OR
 					(reg_q2623 AND symb_decoder(16#bd#)) OR
 					(reg_q2623 AND symb_decoder(16#7f#)) OR
 					(reg_q2623 AND symb_decoder(16#9b#)) OR
 					(reg_q2623 AND symb_decoder(16#bc#)) OR
 					(reg_q2623 AND symb_decoder(16#ae#)) OR
 					(reg_q2623 AND symb_decoder(16#2f#)) OR
 					(reg_q2623 AND symb_decoder(16#71#)) OR
 					(reg_q2623 AND symb_decoder(16#17#)) OR
 					(reg_q2623 AND symb_decoder(16#13#)) OR
 					(reg_q2623 AND symb_decoder(16#02#)) OR
 					(reg_q2623 AND symb_decoder(16#16#)) OR
 					(reg_q2623 AND symb_decoder(16#dc#)) OR
 					(reg_q2623 AND symb_decoder(16#2d#)) OR
 					(reg_q2623 AND symb_decoder(16#a2#)) OR
 					(reg_q2623 AND symb_decoder(16#b7#)) OR
 					(reg_q2623 AND symb_decoder(16#e9#)) OR
 					(reg_q2623 AND symb_decoder(16#5e#)) OR
 					(reg_q2623 AND symb_decoder(16#c2#)) OR
 					(reg_q2623 AND symb_decoder(16#d4#)) OR
 					(reg_q2623 AND symb_decoder(16#4d#)) OR
 					(reg_q2623 AND symb_decoder(16#7a#)) OR
 					(reg_q2623 AND symb_decoder(16#a1#)) OR
 					(reg_q2623 AND symb_decoder(16#3d#)) OR
 					(reg_q2623 AND symb_decoder(16#59#)) OR
 					(reg_q2623 AND symb_decoder(16#9a#)) OR
 					(reg_q2623 AND symb_decoder(16#82#)) OR
 					(reg_q2623 AND symb_decoder(16#ec#)) OR
 					(reg_q2623 AND symb_decoder(16#8a#)) OR
 					(reg_q2623 AND symb_decoder(16#98#)) OR
 					(reg_q2623 AND symb_decoder(16#fa#)) OR
 					(reg_q2623 AND symb_decoder(16#ad#)) OR
 					(reg_q2623 AND symb_decoder(16#ce#)) OR
 					(reg_q2623 AND symb_decoder(16#0a#)) OR
 					(reg_q2623 AND symb_decoder(16#d8#)) OR
 					(reg_q2623 AND symb_decoder(16#3b#)) OR
 					(reg_q2623 AND symb_decoder(16#12#)) OR
 					(reg_q2623 AND symb_decoder(16#90#)) OR
 					(reg_q2623 AND symb_decoder(16#f7#)) OR
 					(reg_q2623 AND symb_decoder(16#b2#)) OR
 					(reg_q2623 AND symb_decoder(16#ff#)) OR
 					(reg_q2623 AND symb_decoder(16#94#)) OR
 					(reg_q2623 AND symb_decoder(16#d3#)) OR
 					(reg_q2623 AND symb_decoder(16#0d#)) OR
 					(reg_q2623 AND symb_decoder(16#ca#)) OR
 					(reg_q2623 AND symb_decoder(16#3f#)) OR
 					(reg_q2623 AND symb_decoder(16#f6#)) OR
 					(reg_q2623 AND symb_decoder(16#da#)) OR
 					(reg_q2623 AND symb_decoder(16#f1#)) OR
 					(reg_q2623 AND symb_decoder(16#db#)) OR
 					(reg_q2623 AND symb_decoder(16#b6#)) OR
 					(reg_q2623 AND symb_decoder(16#5d#)) OR
 					(reg_q2623 AND symb_decoder(16#7b#)) OR
 					(reg_q2623 AND symb_decoder(16#ea#)) OR
 					(reg_q2623 AND symb_decoder(16#de#)) OR
 					(reg_q2623 AND symb_decoder(16#bf#)) OR
 					(reg_q2623 AND symb_decoder(16#ba#)) OR
 					(reg_q2623 AND symb_decoder(16#33#)) OR
 					(reg_q2623 AND symb_decoder(16#29#)) OR
 					(reg_q2623 AND symb_decoder(16#d6#)) OR
 					(reg_q2623 AND symb_decoder(16#fc#)) OR
 					(reg_q2623 AND symb_decoder(16#4a#)) OR
 					(reg_q2623 AND symb_decoder(16#1d#)) OR
 					(reg_q2623 AND symb_decoder(16#f8#)) OR
 					(reg_q2623 AND symb_decoder(16#37#)) OR
 					(reg_q2623 AND symb_decoder(16#9c#)) OR
 					(reg_q2623 AND symb_decoder(16#31#)) OR
 					(reg_q2623 AND symb_decoder(16#0e#)) OR
 					(reg_q2623 AND symb_decoder(16#5c#)) OR
 					(reg_q2623 AND symb_decoder(16#c8#)) OR
 					(reg_q2623 AND symb_decoder(16#04#)) OR
 					(reg_q2623 AND symb_decoder(16#4c#)) OR
 					(reg_q2623 AND symb_decoder(16#e3#)) OR
 					(reg_q2623 AND symb_decoder(16#dd#)) OR
 					(reg_q2623 AND symb_decoder(16#89#)) OR
 					(reg_q2623 AND symb_decoder(16#fb#)) OR
 					(reg_q2623 AND symb_decoder(16#63#)) OR
 					(reg_q2623 AND symb_decoder(16#36#)) OR
 					(reg_q2623 AND symb_decoder(16#66#)) OR
 					(reg_q2623 AND symb_decoder(16#a8#)) OR
 					(reg_q2623 AND symb_decoder(16#60#)) OR
 					(reg_q2623 AND symb_decoder(16#27#)) OR
 					(reg_q2623 AND symb_decoder(16#34#)) OR
 					(reg_q2623 AND symb_decoder(16#e4#)) OR
 					(reg_q2623 AND symb_decoder(16#4e#)) OR
 					(reg_q2623 AND symb_decoder(16#a0#)) OR
 					(reg_q2623 AND symb_decoder(16#e7#)) OR
 					(reg_q2623 AND symb_decoder(16#6c#)) OR
 					(reg_q2623 AND symb_decoder(16#84#)) OR
 					(reg_q2623 AND symb_decoder(16#be#)) OR
 					(reg_q2623 AND symb_decoder(16#9f#)) OR
 					(reg_q2623 AND symb_decoder(16#10#)) OR
 					(reg_q2623 AND symb_decoder(16#44#)) OR
 					(reg_q2623 AND symb_decoder(16#7c#)) OR
 					(reg_q2623 AND symb_decoder(16#52#)) OR
 					(reg_q2623 AND symb_decoder(16#92#)) OR
 					(reg_q2623 AND symb_decoder(16#35#)) OR
 					(reg_q2623 AND symb_decoder(16#c1#)) OR
 					(reg_q2623 AND symb_decoder(16#32#)) OR
 					(reg_q2623 AND symb_decoder(16#a7#)) OR
 					(reg_q2623 AND symb_decoder(16#af#)) OR
 					(reg_q2623 AND symb_decoder(16#81#)) OR
 					(reg_q2623 AND symb_decoder(16#43#)) OR
 					(reg_q2623 AND symb_decoder(16#55#)) OR
 					(reg_q2623 AND symb_decoder(16#ed#)) OR
 					(reg_q2623 AND symb_decoder(16#05#)) OR
 					(reg_q2623 AND symb_decoder(16#ee#)) OR
 					(reg_q2623 AND symb_decoder(16#22#)) OR
 					(reg_q2623 AND symb_decoder(16#06#)) OR
 					(reg_q2623 AND symb_decoder(16#b3#)) OR
 					(reg_q2623 AND symb_decoder(16#95#)) OR
 					(reg_q2623 AND symb_decoder(16#0c#)) OR
 					(reg_q2623 AND symb_decoder(16#e6#)) OR
 					(reg_q2623 AND symb_decoder(16#67#)) OR
 					(reg_q2623 AND symb_decoder(16#c7#)) OR
 					(reg_q2623 AND symb_decoder(16#7e#)) OR
 					(reg_q2623 AND symb_decoder(16#54#)) OR
 					(reg_q2623 AND symb_decoder(16#b9#)) OR
 					(reg_q2623 AND symb_decoder(16#8c#)) OR
 					(reg_q2623 AND symb_decoder(16#48#)) OR
 					(reg_q2623 AND symb_decoder(16#30#)) OR
 					(reg_q2623 AND symb_decoder(16#99#)) OR
 					(reg_q2623 AND symb_decoder(16#c4#)) OR
 					(reg_q2623 AND symb_decoder(16#7d#)) OR
 					(reg_q2623 AND symb_decoder(16#87#)) OR
 					(reg_q2623 AND symb_decoder(16#6b#)) OR
 					(reg_q2623 AND symb_decoder(16#0f#)) OR
 					(reg_q2623 AND symb_decoder(16#d7#)) OR
 					(reg_q2623 AND symb_decoder(16#6e#)) OR
 					(reg_q2623 AND symb_decoder(16#b8#)) OR
 					(reg_q2623 AND symb_decoder(16#1f#)) OR
 					(reg_q2623 AND symb_decoder(16#9d#)) OR
 					(reg_q2623 AND symb_decoder(16#24#)) OR
 					(reg_q2623 AND symb_decoder(16#80#)) OR
 					(reg_q2623 AND symb_decoder(16#2c#)) OR
 					(reg_q2623 AND symb_decoder(16#39#)) OR
 					(reg_q2623 AND symb_decoder(16#58#)) OR
 					(reg_q2623 AND symb_decoder(16#45#)) OR
 					(reg_q2623 AND symb_decoder(16#c9#)) OR
 					(reg_q2623 AND symb_decoder(16#91#)) OR
 					(reg_q2623 AND symb_decoder(16#6d#)) OR
 					(reg_q2623 AND symb_decoder(16#5f#)) OR
 					(reg_q2623 AND symb_decoder(16#5a#)) OR
 					(reg_q2623 AND symb_decoder(16#74#)) OR
 					(reg_q2623 AND symb_decoder(16#64#)) OR
 					(reg_q2623 AND symb_decoder(16#93#)) OR
 					(reg_q2623 AND symb_decoder(16#fd#)) OR
 					(reg_q2623 AND symb_decoder(16#19#)) OR
 					(reg_q2623 AND symb_decoder(16#f5#)) OR
 					(reg_q2623 AND symb_decoder(16#e8#)) OR
 					(reg_q2623 AND symb_decoder(16#26#)) OR
 					(reg_q2623 AND symb_decoder(16#f3#)) OR
 					(reg_q2623 AND symb_decoder(16#61#)) OR
 					(reg_q2623 AND symb_decoder(16#cd#)) OR
 					(reg_q2623 AND symb_decoder(16#f0#)) OR
 					(reg_q2623 AND symb_decoder(16#b5#)) OR
 					(reg_q2623 AND symb_decoder(16#21#)) OR
 					(reg_q2623 AND symb_decoder(16#11#)) OR
 					(reg_q2623 AND symb_decoder(16#83#)) OR
 					(reg_q2623 AND symb_decoder(16#86#)) OR
 					(reg_q2623 AND symb_decoder(16#d9#)) OR
 					(reg_q2623 AND symb_decoder(16#df#)) OR
 					(reg_q2623 AND symb_decoder(16#85#)) OR
 					(reg_q2623 AND symb_decoder(16#38#)) OR
 					(reg_q2623 AND symb_decoder(16#53#)) OR
 					(reg_q2623 AND symb_decoder(16#2e#)) OR
 					(reg_q2623 AND symb_decoder(16#28#)) OR
 					(reg_q2623 AND symb_decoder(16#69#)) OR
 					(reg_q2623 AND symb_decoder(16#ef#)) OR
 					(reg_q2623 AND symb_decoder(16#aa#)) OR
 					(reg_q2623 AND symb_decoder(16#97#)) OR
 					(reg_q2623 AND symb_decoder(16#a6#)) OR
 					(reg_q2623 AND symb_decoder(16#3e#)) OR
 					(reg_q2623 AND symb_decoder(16#8d#)) OR
 					(reg_q2623 AND symb_decoder(16#4b#)) OR
 					(reg_q2623 AND symb_decoder(16#78#)) OR
 					(reg_q2623 AND symb_decoder(16#e0#)) OR
 					(reg_q2623 AND symb_decoder(16#c0#)) OR
 					(reg_q2623 AND symb_decoder(16#41#)) OR
 					(reg_q2623 AND symb_decoder(16#23#)) OR
 					(reg_q2623 AND symb_decoder(16#f4#)) OR
 					(reg_q2623 AND symb_decoder(16#25#)) OR
 					(reg_q2623 AND symb_decoder(16#ac#)) OR
 					(reg_q2623 AND symb_decoder(16#46#)) OR
 					(reg_q2623 AND symb_decoder(16#fe#)) OR
 					(reg_q2623 AND symb_decoder(16#d1#)) OR
 					(reg_q2623 AND symb_decoder(16#c6#)) OR
 					(reg_q2623 AND symb_decoder(16#50#)) OR
 					(reg_q2623 AND symb_decoder(16#88#)) OR
 					(reg_q2623 AND symb_decoder(16#00#)) OR
 					(reg_q2623 AND symb_decoder(16#20#)) OR
 					(reg_q2623 AND symb_decoder(16#d5#)) OR
 					(reg_q2623 AND symb_decoder(16#75#)) OR
 					(reg_q2623 AND symb_decoder(16#08#)) OR
 					(reg_q2623 AND symb_decoder(16#77#)) OR
 					(reg_q2623 AND symb_decoder(16#ab#)) OR
 					(reg_q2623 AND symb_decoder(16#9e#)) OR
 					(reg_q2623 AND symb_decoder(16#5b#)) OR
 					(reg_q2623 AND symb_decoder(16#70#)) OR
 					(reg_q2623 AND symb_decoder(16#0b#)) OR
 					(reg_q2623 AND symb_decoder(16#8b#)) OR
 					(reg_q2623 AND symb_decoder(16#eb#)) OR
 					(reg_q2623 AND symb_decoder(16#cf#)) OR
 					(reg_q2623 AND symb_decoder(16#bb#)) OR
 					(reg_q2623 AND symb_decoder(16#18#)) OR
 					(reg_q2623 AND symb_decoder(16#d0#)) OR
 					(reg_q2623 AND symb_decoder(16#62#)) OR
 					(reg_q2623 AND symb_decoder(16#c3#)) OR
 					(reg_q2623 AND symb_decoder(16#09#)) OR
 					(reg_q2623 AND symb_decoder(16#51#)) OR
 					(reg_q2623 AND symb_decoder(16#2b#)) OR
 					(reg_q2623 AND symb_decoder(16#c5#)) OR
 					(reg_q2623 AND symb_decoder(16#73#)) OR
 					(reg_q2623 AND symb_decoder(16#03#)) OR
 					(reg_q2623 AND symb_decoder(16#1a#)) OR
 					(reg_q2623 AND symb_decoder(16#07#)) OR
 					(reg_q2623 AND symb_decoder(16#6a#)) OR
 					(reg_q2623 AND symb_decoder(16#b4#)) OR
 					(reg_q2623 AND symb_decoder(16#6f#)) OR
 					(reg_q2623 AND symb_decoder(16#14#)) OR
 					(reg_q2623 AND symb_decoder(16#f9#)) OR
 					(reg_q2623 AND symb_decoder(16#56#)) OR
 					(reg_q2623 AND symb_decoder(16#a3#)) OR
 					(reg_q2623 AND symb_decoder(16#b1#)) OR
 					(reg_q2623 AND symb_decoder(16#a9#)) OR
 					(reg_q2623 AND symb_decoder(16#49#)) OR
 					(reg_q2623 AND symb_decoder(16#68#)) OR
 					(reg_q2623 AND symb_decoder(16#a4#)) OR
 					(reg_q2623 AND symb_decoder(16#1b#)) OR
 					(reg_q2623 AND symb_decoder(16#76#)) OR
 					(reg_q2623 AND symb_decoder(16#8e#)) OR
 					(reg_q2623 AND symb_decoder(16#01#)) OR
 					(reg_q2623 AND symb_decoder(16#3c#)) OR
 					(reg_q2623 AND symb_decoder(16#d2#)) OR
 					(reg_q2623 AND symb_decoder(16#96#)) OR
 					(reg_q2623 AND symb_decoder(16#cc#)) OR
 					(reg_q2623 AND symb_decoder(16#2a#)) OR
 					(reg_q2623 AND symb_decoder(16#8f#)) OR
 					(reg_q2623 AND symb_decoder(16#57#));
reg_q499_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q498 AND symb_decoder(16#73#)) OR
 					(reg_q498 AND symb_decoder(16#53#));
reg_q663_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q662 AND symb_decoder(16#0c#)) OR
 					(reg_q662 AND symb_decoder(16#0a#)) OR
 					(reg_q662 AND symb_decoder(16#20#)) OR
 					(reg_q662 AND symb_decoder(16#09#)) OR
 					(reg_q662 AND symb_decoder(16#0d#));
reg_q520_in <= (reg_q518 AND symb_decoder(16#69#)) OR
 					(reg_q518 AND symb_decoder(16#49#));
reg_q667_in <= (reg_q665 AND symb_decoder(16#72#)) OR
 					(reg_q665 AND symb_decoder(16#52#));
reg_q101_in <= (reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q100 AND symb_decoder(16#70#)) OR
 					(reg_q100 AND symb_decoder(16#50#));
reg_q1206_in <= (reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q1205 AND symb_decoder(16#76#)) OR
 					(reg_q1205 AND symb_decoder(16#56#));
reg_q1978_in <= (reg_q2757 AND symb_decoder(16#2f#));
reg_q30_in <= (reg_q28 AND symb_decoder(16#57#)) OR
 					(reg_q28 AND symb_decoder(16#77#));
reg_q1063_in <= (reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q1062 AND symb_decoder(16#54#)) OR
 					(reg_q1062 AND symb_decoder(16#74#));
reg_fullgraph15_init <= "0000";

reg_fullgraph15_sel <= "00000" & reg_q1063_in & reg_q30_in & reg_q1978_in & reg_q1206_in & reg_q101_in & reg_q667_in & reg_q520_in & reg_q663_in & reg_q499_in & reg_q2625_in & reg_q1682_in;

	--coder fullgraph15
with reg_fullgraph15_sel select
reg_fullgraph15_in <=
	"0001" when "0000000000000001",
	"0010" when "0000000000000010",
	"0011" when "0000000000000100",
	"0100" when "0000000000001000",
	"0101" when "0000000000010000",
	"0110" when "0000000000100000",
	"0111" when "0000000001000000",
	"1000" when "0000000010000000",
	"1001" when "0000000100000000",
	"1010" when "0000001000000000",
	"1011" when "0000010000000000",
	"0000" when others;
 --end coder

	p_reg_fullgraph15: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph15 <= reg_fullgraph15_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph15 <= reg_fullgraph15_init;
        else
          reg_fullgraph15 <= reg_fullgraph15_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph15

		reg_q1682 <= '1' when reg_fullgraph15 = "0001" else '0'; 
		reg_q2625 <= '1' when reg_fullgraph15 = "0010" else '0'; 
		reg_q499 <= '1' when reg_fullgraph15 = "0011" else '0'; 
		reg_q663 <= '1' when reg_fullgraph15 = "0100" else '0'; 
		reg_q520 <= '1' when reg_fullgraph15 = "0101" else '0'; 
		reg_q667 <= '1' when reg_fullgraph15 = "0110" else '0'; 
		reg_q101 <= '1' when reg_fullgraph15 = "0111" else '0'; 
		reg_q1206 <= '1' when reg_fullgraph15 = "1000" else '0'; 
		reg_q1978 <= '1' when reg_fullgraph15 = "1001" else '0'; 
		reg_q30 <= '1' when reg_fullgraph15 = "1010" else '0'; 
		reg_q1063 <= '1' when reg_fullgraph15 = "1011" else '0'; 
--end decoder 

reg_q945_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q945 AND symb_decoder(16#d2#)) OR
 					(reg_q945 AND symb_decoder(16#d5#)) OR
 					(reg_q945 AND symb_decoder(16#6c#)) OR
 					(reg_q945 AND symb_decoder(16#64#)) OR
 					(reg_q945 AND symb_decoder(16#74#)) OR
 					(reg_q945 AND symb_decoder(16#3e#)) OR
 					(reg_q945 AND symb_decoder(16#f2#)) OR
 					(reg_q945 AND symb_decoder(16#85#)) OR
 					(reg_q945 AND symb_decoder(16#b7#)) OR
 					(reg_q945 AND symb_decoder(16#93#)) OR
 					(reg_q945 AND symb_decoder(16#e6#)) OR
 					(reg_q945 AND symb_decoder(16#eb#)) OR
 					(reg_q945 AND symb_decoder(16#55#)) OR
 					(reg_q945 AND symb_decoder(16#07#)) OR
 					(reg_q945 AND symb_decoder(16#77#)) OR
 					(reg_q945 AND symb_decoder(16#df#)) OR
 					(reg_q945 AND symb_decoder(16#5e#)) OR
 					(reg_q945 AND symb_decoder(16#50#)) OR
 					(reg_q945 AND symb_decoder(16#4a#)) OR
 					(reg_q945 AND symb_decoder(16#ba#)) OR
 					(reg_q945 AND symb_decoder(16#29#)) OR
 					(reg_q945 AND symb_decoder(16#ae#)) OR
 					(reg_q945 AND symb_decoder(16#92#)) OR
 					(reg_q945 AND symb_decoder(16#e4#)) OR
 					(reg_q945 AND symb_decoder(16#65#)) OR
 					(reg_q945 AND symb_decoder(16#7b#)) OR
 					(reg_q945 AND symb_decoder(16#66#)) OR
 					(reg_q945 AND symb_decoder(16#cd#)) OR
 					(reg_q945 AND symb_decoder(16#c4#)) OR
 					(reg_q945 AND symb_decoder(16#8d#)) OR
 					(reg_q945 AND symb_decoder(16#9c#)) OR
 					(reg_q945 AND symb_decoder(16#62#)) OR
 					(reg_q945 AND symb_decoder(16#2a#)) OR
 					(reg_q945 AND symb_decoder(16#ec#)) OR
 					(reg_q945 AND symb_decoder(16#41#)) OR
 					(reg_q945 AND symb_decoder(16#76#)) OR
 					(reg_q945 AND symb_decoder(16#ef#)) OR
 					(reg_q945 AND symb_decoder(16#91#)) OR
 					(reg_q945 AND symb_decoder(16#fa#)) OR
 					(reg_q945 AND symb_decoder(16#23#)) OR
 					(reg_q945 AND symb_decoder(16#ad#)) OR
 					(reg_q945 AND symb_decoder(16#30#)) OR
 					(reg_q945 AND symb_decoder(16#e9#)) OR
 					(reg_q945 AND symb_decoder(16#5a#)) OR
 					(reg_q945 AND symb_decoder(16#49#)) OR
 					(reg_q945 AND symb_decoder(16#0a#)) OR
 					(reg_q945 AND symb_decoder(16#78#)) OR
 					(reg_q945 AND symb_decoder(16#67#)) OR
 					(reg_q945 AND symb_decoder(16#a8#)) OR
 					(reg_q945 AND symb_decoder(16#18#)) OR
 					(reg_q945 AND symb_decoder(16#fb#)) OR
 					(reg_q945 AND symb_decoder(16#d4#)) OR
 					(reg_q945 AND symb_decoder(16#cc#)) OR
 					(reg_q945 AND symb_decoder(16#ab#)) OR
 					(reg_q945 AND symb_decoder(16#60#)) OR
 					(reg_q945 AND symb_decoder(16#2e#)) OR
 					(reg_q945 AND symb_decoder(16#1e#)) OR
 					(reg_q945 AND symb_decoder(16#38#)) OR
 					(reg_q945 AND symb_decoder(16#72#)) OR
 					(reg_q945 AND symb_decoder(16#75#)) OR
 					(reg_q945 AND symb_decoder(16#3d#)) OR
 					(reg_q945 AND symb_decoder(16#95#)) OR
 					(reg_q945 AND symb_decoder(16#09#)) OR
 					(reg_q945 AND symb_decoder(16#89#)) OR
 					(reg_q945 AND symb_decoder(16#f7#)) OR
 					(reg_q945 AND symb_decoder(16#45#)) OR
 					(reg_q945 AND symb_decoder(16#c8#)) OR
 					(reg_q945 AND symb_decoder(16#73#)) OR
 					(reg_q945 AND symb_decoder(16#44#)) OR
 					(reg_q945 AND symb_decoder(16#4f#)) OR
 					(reg_q945 AND symb_decoder(16#da#)) OR
 					(reg_q945 AND symb_decoder(16#8b#)) OR
 					(reg_q945 AND symb_decoder(16#08#)) OR
 					(reg_q945 AND symb_decoder(16#1f#)) OR
 					(reg_q945 AND symb_decoder(16#ed#)) OR
 					(reg_q945 AND symb_decoder(16#cf#)) OR
 					(reg_q945 AND symb_decoder(16#dd#)) OR
 					(reg_q945 AND symb_decoder(16#80#)) OR
 					(reg_q945 AND symb_decoder(16#97#)) OR
 					(reg_q945 AND symb_decoder(16#3c#)) OR
 					(reg_q945 AND symb_decoder(16#c0#)) OR
 					(reg_q945 AND symb_decoder(16#a3#)) OR
 					(reg_q945 AND symb_decoder(16#3a#)) OR
 					(reg_q945 AND symb_decoder(16#fe#)) OR
 					(reg_q945 AND symb_decoder(16#52#)) OR
 					(reg_q945 AND symb_decoder(16#02#)) OR
 					(reg_q945 AND symb_decoder(16#43#)) OR
 					(reg_q945 AND symb_decoder(16#42#)) OR
 					(reg_q945 AND symb_decoder(16#01#)) OR
 					(reg_q945 AND symb_decoder(16#15#)) OR
 					(reg_q945 AND symb_decoder(16#4c#)) OR
 					(reg_q945 AND symb_decoder(16#9a#)) OR
 					(reg_q945 AND symb_decoder(16#79#)) OR
 					(reg_q945 AND symb_decoder(16#96#)) OR
 					(reg_q945 AND symb_decoder(16#54#)) OR
 					(reg_q945 AND symb_decoder(16#84#)) OR
 					(reg_q945 AND symb_decoder(16#d7#)) OR
 					(reg_q945 AND symb_decoder(16#f1#)) OR
 					(reg_q945 AND symb_decoder(16#06#)) OR
 					(reg_q945 AND symb_decoder(16#56#)) OR
 					(reg_q945 AND symb_decoder(16#3f#)) OR
 					(reg_q945 AND symb_decoder(16#27#)) OR
 					(reg_q945 AND symb_decoder(16#c7#)) OR
 					(reg_q945 AND symb_decoder(16#8f#)) OR
 					(reg_q945 AND symb_decoder(16#6e#)) OR
 					(reg_q945 AND symb_decoder(16#f4#)) OR
 					(reg_q945 AND symb_decoder(16#10#)) OR
 					(reg_q945 AND symb_decoder(16#20#)) OR
 					(reg_q945 AND symb_decoder(16#48#)) OR
 					(reg_q945 AND symb_decoder(16#e2#)) OR
 					(reg_q945 AND symb_decoder(16#c6#)) OR
 					(reg_q945 AND symb_decoder(16#9d#)) OR
 					(reg_q945 AND symb_decoder(16#0c#)) OR
 					(reg_q945 AND symb_decoder(16#f6#)) OR
 					(reg_q945 AND symb_decoder(16#31#)) OR
 					(reg_q945 AND symb_decoder(16#a4#)) OR
 					(reg_q945 AND symb_decoder(16#d9#)) OR
 					(reg_q945 AND symb_decoder(16#a6#)) OR
 					(reg_q945 AND symb_decoder(16#a5#)) OR
 					(reg_q945 AND symb_decoder(16#9e#)) OR
 					(reg_q945 AND symb_decoder(16#e5#)) OR
 					(reg_q945 AND symb_decoder(16#0f#)) OR
 					(reg_q945 AND symb_decoder(16#de#)) OR
 					(reg_q945 AND symb_decoder(16#39#)) OR
 					(reg_q945 AND symb_decoder(16#c5#)) OR
 					(reg_q945 AND symb_decoder(16#1a#)) OR
 					(reg_q945 AND symb_decoder(16#81#)) OR
 					(reg_q945 AND symb_decoder(16#70#)) OR
 					(reg_q945 AND symb_decoder(16#12#)) OR
 					(reg_q945 AND symb_decoder(16#05#)) OR
 					(reg_q945 AND symb_decoder(16#37#)) OR
 					(reg_q945 AND symb_decoder(16#fc#)) OR
 					(reg_q945 AND symb_decoder(16#b9#)) OR
 					(reg_q945 AND symb_decoder(16#be#)) OR
 					(reg_q945 AND symb_decoder(16#d6#)) OR
 					(reg_q945 AND symb_decoder(16#03#)) OR
 					(reg_q945 AND symb_decoder(16#bd#)) OR
 					(reg_q945 AND symb_decoder(16#bb#)) OR
 					(reg_q945 AND symb_decoder(16#b6#)) OR
 					(reg_q945 AND symb_decoder(16#22#)) OR
 					(reg_q945 AND symb_decoder(16#ff#)) OR
 					(reg_q945 AND symb_decoder(16#57#)) OR
 					(reg_q945 AND symb_decoder(16#c3#)) OR
 					(reg_q945 AND symb_decoder(16#8e#)) OR
 					(reg_q945 AND symb_decoder(16#d1#)) OR
 					(reg_q945 AND symb_decoder(16#28#)) OR
 					(reg_q945 AND symb_decoder(16#21#)) OR
 					(reg_q945 AND symb_decoder(16#ce#)) OR
 					(reg_q945 AND symb_decoder(16#7a#)) OR
 					(reg_q945 AND symb_decoder(16#94#)) OR
 					(reg_q945 AND symb_decoder(16#98#)) OR
 					(reg_q945 AND symb_decoder(16#b2#)) OR
 					(reg_q945 AND symb_decoder(16#0e#)) OR
 					(reg_q945 AND symb_decoder(16#2c#)) OR
 					(reg_q945 AND symb_decoder(16#3b#)) OR
 					(reg_q945 AND symb_decoder(16#e0#)) OR
 					(reg_q945 AND symb_decoder(16#c2#)) OR
 					(reg_q945 AND symb_decoder(16#46#)) OR
 					(reg_q945 AND symb_decoder(16#af#)) OR
 					(reg_q945 AND symb_decoder(16#8c#)) OR
 					(reg_q945 AND symb_decoder(16#63#)) OR
 					(reg_q945 AND symb_decoder(16#53#)) OR
 					(reg_q945 AND symb_decoder(16#69#)) OR
 					(reg_q945 AND symb_decoder(16#6d#)) OR
 					(reg_q945 AND symb_decoder(16#6f#)) OR
 					(reg_q945 AND symb_decoder(16#cb#)) OR
 					(reg_q945 AND symb_decoder(16#71#)) OR
 					(reg_q945 AND symb_decoder(16#1b#)) OR
 					(reg_q945 AND symb_decoder(16#25#)) OR
 					(reg_q945 AND symb_decoder(16#f8#)) OR
 					(reg_q945 AND symb_decoder(16#34#)) OR
 					(reg_q945 AND symb_decoder(16#32#)) OR
 					(reg_q945 AND symb_decoder(16#d0#)) OR
 					(reg_q945 AND symb_decoder(16#59#)) OR
 					(reg_q945 AND symb_decoder(16#4e#)) OR
 					(reg_q945 AND symb_decoder(16#e8#)) OR
 					(reg_q945 AND symb_decoder(16#36#)) OR
 					(reg_q945 AND symb_decoder(16#88#)) OR
 					(reg_q945 AND symb_decoder(16#e1#)) OR
 					(reg_q945 AND symb_decoder(16#17#)) OR
 					(reg_q945 AND symb_decoder(16#86#)) OR
 					(reg_q945 AND symb_decoder(16#26#)) OR
 					(reg_q945 AND symb_decoder(16#5d#)) OR
 					(reg_q945 AND symb_decoder(16#0b#)) OR
 					(reg_q945 AND symb_decoder(16#68#)) OR
 					(reg_q945 AND symb_decoder(16#1d#)) OR
 					(reg_q945 AND symb_decoder(16#b4#)) OR
 					(reg_q945 AND symb_decoder(16#7f#)) OR
 					(reg_q945 AND symb_decoder(16#fd#)) OR
 					(reg_q945 AND symb_decoder(16#e7#)) OR
 					(reg_q945 AND symb_decoder(16#a7#)) OR
 					(reg_q945 AND symb_decoder(16#13#)) OR
 					(reg_q945 AND symb_decoder(16#f3#)) OR
 					(reg_q945 AND symb_decoder(16#dc#)) OR
 					(reg_q945 AND symb_decoder(16#f9#)) OR
 					(reg_q945 AND symb_decoder(16#14#)) OR
 					(reg_q945 AND symb_decoder(16#b0#)) OR
 					(reg_q945 AND symb_decoder(16#90#)) OR
 					(reg_q945 AND symb_decoder(16#7d#)) OR
 					(reg_q945 AND symb_decoder(16#6b#)) OR
 					(reg_q945 AND symb_decoder(16#ac#)) OR
 					(reg_q945 AND symb_decoder(16#99#)) OR
 					(reg_q945 AND symb_decoder(16#82#)) OR
 					(reg_q945 AND symb_decoder(16#0d#)) OR
 					(reg_q945 AND symb_decoder(16#4d#)) OR
 					(reg_q945 AND symb_decoder(16#b3#)) OR
 					(reg_q945 AND symb_decoder(16#11#)) OR
 					(reg_q945 AND symb_decoder(16#a2#)) OR
 					(reg_q945 AND symb_decoder(16#bf#)) OR
 					(reg_q945 AND symb_decoder(16#a0#)) OR
 					(reg_q945 AND symb_decoder(16#19#)) OR
 					(reg_q945 AND symb_decoder(16#58#)) OR
 					(reg_q945 AND symb_decoder(16#1c#)) OR
 					(reg_q945 AND symb_decoder(16#35#)) OR
 					(reg_q945 AND symb_decoder(16#5c#)) OR
 					(reg_q945 AND symb_decoder(16#b1#)) OR
 					(reg_q945 AND symb_decoder(16#8a#)) OR
 					(reg_q945 AND symb_decoder(16#c9#)) OR
 					(reg_q945 AND symb_decoder(16#16#)) OR
 					(reg_q945 AND symb_decoder(16#db#)) OR
 					(reg_q945 AND symb_decoder(16#61#)) OR
 					(reg_q945 AND symb_decoder(16#9f#)) OR
 					(reg_q945 AND symb_decoder(16#2d#)) OR
 					(reg_q945 AND symb_decoder(16#ea#)) OR
 					(reg_q945 AND symb_decoder(16#40#)) OR
 					(reg_q945 AND symb_decoder(16#5f#)) OR
 					(reg_q945 AND symb_decoder(16#b5#)) OR
 					(reg_q945 AND symb_decoder(16#e3#)) OR
 					(reg_q945 AND symb_decoder(16#6a#)) OR
 					(reg_q945 AND symb_decoder(16#00#)) OR
 					(reg_q945 AND symb_decoder(16#83#)) OR
 					(reg_q945 AND symb_decoder(16#ee#)) OR
 					(reg_q945 AND symb_decoder(16#b8#)) OR
 					(reg_q945 AND symb_decoder(16#4b#)) OR
 					(reg_q945 AND symb_decoder(16#c1#)) OR
 					(reg_q945 AND symb_decoder(16#5b#)) OR
 					(reg_q945 AND symb_decoder(16#24#)) OR
 					(reg_q945 AND symb_decoder(16#f5#)) OR
 					(reg_q945 AND symb_decoder(16#7e#)) OR
 					(reg_q945 AND symb_decoder(16#04#)) OR
 					(reg_q945 AND symb_decoder(16#47#)) OR
 					(reg_q945 AND symb_decoder(16#a9#)) OR
 					(reg_q945 AND symb_decoder(16#a1#)) OR
 					(reg_q945 AND symb_decoder(16#d3#)) OR
 					(reg_q945 AND symb_decoder(16#ca#)) OR
 					(reg_q945 AND symb_decoder(16#33#)) OR
 					(reg_q945 AND symb_decoder(16#9b#)) OR
 					(reg_q945 AND symb_decoder(16#f0#)) OR
 					(reg_q945 AND symb_decoder(16#7c#)) OR
 					(reg_q945 AND symb_decoder(16#bc#)) OR
 					(reg_q945 AND symb_decoder(16#2b#)) OR
 					(reg_q945 AND symb_decoder(16#51#)) OR
 					(reg_q945 AND symb_decoder(16#aa#)) OR
 					(reg_q945 AND symb_decoder(16#87#)) OR
 					(reg_q945 AND symb_decoder(16#2f#)) OR
 					(reg_q945 AND symb_decoder(16#d8#));
reg_q945_init <= '0' ;
	p_reg_q945: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q945 <= reg_q945_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q945 <= reg_q945_init;
        else
          reg_q945 <= reg_q945_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2554_in <= (reg_q2526 AND symb_decoder(16#ff#)) OR
 					(reg_q2526 AND symb_decoder(16#6d#)) OR
 					(reg_q2526 AND symb_decoder(16#24#)) OR
 					(reg_q2526 AND symb_decoder(16#20#)) OR
 					(reg_q2526 AND symb_decoder(16#8e#)) OR
 					(reg_q2526 AND symb_decoder(16#70#)) OR
 					(reg_q2526 AND symb_decoder(16#62#)) OR
 					(reg_q2526 AND symb_decoder(16#a1#)) OR
 					(reg_q2526 AND symb_decoder(16#0b#)) OR
 					(reg_q2526 AND symb_decoder(16#6c#)) OR
 					(reg_q2526 AND symb_decoder(16#e6#)) OR
 					(reg_q2526 AND symb_decoder(16#07#)) OR
 					(reg_q2526 AND symb_decoder(16#89#)) OR
 					(reg_q2526 AND symb_decoder(16#46#)) OR
 					(reg_q2526 AND symb_decoder(16#60#)) OR
 					(reg_q2526 AND symb_decoder(16#c1#)) OR
 					(reg_q2526 AND symb_decoder(16#90#)) OR
 					(reg_q2526 AND symb_decoder(16#86#)) OR
 					(reg_q2526 AND symb_decoder(16#6e#)) OR
 					(reg_q2526 AND symb_decoder(16#82#)) OR
 					(reg_q2526 AND symb_decoder(16#32#)) OR
 					(reg_q2526 AND symb_decoder(16#22#)) OR
 					(reg_q2526 AND symb_decoder(16#17#)) OR
 					(reg_q2526 AND symb_decoder(16#ae#)) OR
 					(reg_q2526 AND symb_decoder(16#71#)) OR
 					(reg_q2526 AND symb_decoder(16#c2#)) OR
 					(reg_q2526 AND symb_decoder(16#ba#)) OR
 					(reg_q2526 AND symb_decoder(16#51#)) OR
 					(reg_q2526 AND symb_decoder(16#95#)) OR
 					(reg_q2526 AND symb_decoder(16#8d#)) OR
 					(reg_q2526 AND symb_decoder(16#18#)) OR
 					(reg_q2526 AND symb_decoder(16#97#)) OR
 					(reg_q2526 AND symb_decoder(16#cc#)) OR
 					(reg_q2526 AND symb_decoder(16#a5#)) OR
 					(reg_q2526 AND symb_decoder(16#ea#)) OR
 					(reg_q2526 AND symb_decoder(16#aa#)) OR
 					(reg_q2526 AND symb_decoder(16#74#)) OR
 					(reg_q2526 AND symb_decoder(16#d8#)) OR
 					(reg_q2526 AND symb_decoder(16#b2#)) OR
 					(reg_q2526 AND symb_decoder(16#fa#)) OR
 					(reg_q2526 AND symb_decoder(16#69#)) OR
 					(reg_q2526 AND symb_decoder(16#48#)) OR
 					(reg_q2526 AND symb_decoder(16#25#)) OR
 					(reg_q2526 AND symb_decoder(16#1f#)) OR
 					(reg_q2526 AND symb_decoder(16#ca#)) OR
 					(reg_q2526 AND symb_decoder(16#7c#)) OR
 					(reg_q2526 AND symb_decoder(16#49#)) OR
 					(reg_q2526 AND symb_decoder(16#92#)) OR
 					(reg_q2526 AND symb_decoder(16#e7#)) OR
 					(reg_q2526 AND symb_decoder(16#12#)) OR
 					(reg_q2526 AND symb_decoder(16#2e#)) OR
 					(reg_q2526 AND symb_decoder(16#59#)) OR
 					(reg_q2526 AND symb_decoder(16#73#)) OR
 					(reg_q2526 AND symb_decoder(16#4d#)) OR
 					(reg_q2526 AND symb_decoder(16#0a#)) OR
 					(reg_q2526 AND symb_decoder(16#6f#)) OR
 					(reg_q2526 AND symb_decoder(16#a7#)) OR
 					(reg_q2526 AND symb_decoder(16#7f#)) OR
 					(reg_q2526 AND symb_decoder(16#5b#)) OR
 					(reg_q2526 AND symb_decoder(16#1e#)) OR
 					(reg_q2526 AND symb_decoder(16#ab#)) OR
 					(reg_q2526 AND symb_decoder(16#dc#)) OR
 					(reg_q2526 AND symb_decoder(16#bc#)) OR
 					(reg_q2526 AND symb_decoder(16#a8#)) OR
 					(reg_q2526 AND symb_decoder(16#fc#)) OR
 					(reg_q2526 AND symb_decoder(16#45#)) OR
 					(reg_q2526 AND symb_decoder(16#78#)) OR
 					(reg_q2526 AND symb_decoder(16#58#)) OR
 					(reg_q2526 AND symb_decoder(16#3a#)) OR
 					(reg_q2526 AND symb_decoder(16#66#)) OR
 					(reg_q2526 AND symb_decoder(16#42#)) OR
 					(reg_q2526 AND symb_decoder(16#b7#)) OR
 					(reg_q2526 AND symb_decoder(16#27#)) OR
 					(reg_q2526 AND symb_decoder(16#f0#)) OR
 					(reg_q2526 AND symb_decoder(16#e2#)) OR
 					(reg_q2526 AND symb_decoder(16#c7#)) OR
 					(reg_q2526 AND symb_decoder(16#91#)) OR
 					(reg_q2526 AND symb_decoder(16#88#)) OR
 					(reg_q2526 AND symb_decoder(16#85#)) OR
 					(reg_q2526 AND symb_decoder(16#0c#)) OR
 					(reg_q2526 AND symb_decoder(16#2b#)) OR
 					(reg_q2526 AND symb_decoder(16#2d#)) OR
 					(reg_q2526 AND symb_decoder(16#d2#)) OR
 					(reg_q2526 AND symb_decoder(16#b4#)) OR
 					(reg_q2526 AND symb_decoder(16#ce#)) OR
 					(reg_q2526 AND symb_decoder(16#df#)) OR
 					(reg_q2526 AND symb_decoder(16#9d#)) OR
 					(reg_q2526 AND symb_decoder(16#cf#)) OR
 					(reg_q2526 AND symb_decoder(16#d3#)) OR
 					(reg_q2526 AND symb_decoder(16#a6#)) OR
 					(reg_q2526 AND symb_decoder(16#00#)) OR
 					(reg_q2526 AND symb_decoder(16#3c#)) OR
 					(reg_q2526 AND symb_decoder(16#c5#)) OR
 					(reg_q2526 AND symb_decoder(16#bd#)) OR
 					(reg_q2526 AND symb_decoder(16#4c#)) OR
 					(reg_q2526 AND symb_decoder(16#10#)) OR
 					(reg_q2526 AND symb_decoder(16#84#)) OR
 					(reg_q2526 AND symb_decoder(16#1b#)) OR
 					(reg_q2526 AND symb_decoder(16#65#)) OR
 					(reg_q2526 AND symb_decoder(16#a4#)) OR
 					(reg_q2526 AND symb_decoder(16#23#)) OR
 					(reg_q2526 AND symb_decoder(16#3b#)) OR
 					(reg_q2526 AND symb_decoder(16#31#)) OR
 					(reg_q2526 AND symb_decoder(16#52#)) OR
 					(reg_q2526 AND symb_decoder(16#50#)) OR
 					(reg_q2526 AND symb_decoder(16#bb#)) OR
 					(reg_q2526 AND symb_decoder(16#a0#)) OR
 					(reg_q2526 AND symb_decoder(16#53#)) OR
 					(reg_q2526 AND symb_decoder(16#68#)) OR
 					(reg_q2526 AND symb_decoder(16#30#)) OR
 					(reg_q2526 AND symb_decoder(16#b0#)) OR
 					(reg_q2526 AND symb_decoder(16#1c#)) OR
 					(reg_q2526 AND symb_decoder(16#03#)) OR
 					(reg_q2526 AND symb_decoder(16#09#)) OR
 					(reg_q2526 AND symb_decoder(16#40#)) OR
 					(reg_q2526 AND symb_decoder(16#4a#)) OR
 					(reg_q2526 AND symb_decoder(16#f7#)) OR
 					(reg_q2526 AND symb_decoder(16#d7#)) OR
 					(reg_q2526 AND symb_decoder(16#7a#)) OR
 					(reg_q2526 AND symb_decoder(16#08#)) OR
 					(reg_q2526 AND symb_decoder(16#36#)) OR
 					(reg_q2526 AND symb_decoder(16#c8#)) OR
 					(reg_q2526 AND symb_decoder(16#9a#)) OR
 					(reg_q2526 AND symb_decoder(16#a9#)) OR
 					(reg_q2526 AND symb_decoder(16#83#)) OR
 					(reg_q2526 AND symb_decoder(16#be#)) OR
 					(reg_q2526 AND symb_decoder(16#6a#)) OR
 					(reg_q2526 AND symb_decoder(16#b6#)) OR
 					(reg_q2526 AND symb_decoder(16#c0#)) OR
 					(reg_q2526 AND symb_decoder(16#9e#)) OR
 					(reg_q2526 AND symb_decoder(16#38#)) OR
 					(reg_q2526 AND symb_decoder(16#f2#)) OR
 					(reg_q2526 AND symb_decoder(16#a3#)) OR
 					(reg_q2526 AND symb_decoder(16#34#)) OR
 					(reg_q2526 AND symb_decoder(16#57#)) OR
 					(reg_q2526 AND symb_decoder(16#11#)) OR
 					(reg_q2526 AND symb_decoder(16#81#)) OR
 					(reg_q2526 AND symb_decoder(16#99#)) OR
 					(reg_q2526 AND symb_decoder(16#21#)) OR
 					(reg_q2526 AND symb_decoder(16#26#)) OR
 					(reg_q2526 AND symb_decoder(16#af#)) OR
 					(reg_q2526 AND symb_decoder(16#7b#)) OR
 					(reg_q2526 AND symb_decoder(16#c6#)) OR
 					(reg_q2526 AND symb_decoder(16#8b#)) OR
 					(reg_q2526 AND symb_decoder(16#94#)) OR
 					(reg_q2526 AND symb_decoder(16#1a#)) OR
 					(reg_q2526 AND symb_decoder(16#02#)) OR
 					(reg_q2526 AND symb_decoder(16#96#)) OR
 					(reg_q2526 AND symb_decoder(16#33#)) OR
 					(reg_q2526 AND symb_decoder(16#d1#)) OR
 					(reg_q2526 AND symb_decoder(16#61#)) OR
 					(reg_q2526 AND symb_decoder(16#2c#)) OR
 					(reg_q2526 AND symb_decoder(16#39#)) OR
 					(reg_q2526 AND symb_decoder(16#35#)) OR
 					(reg_q2526 AND symb_decoder(16#d6#)) OR
 					(reg_q2526 AND symb_decoder(16#5a#)) OR
 					(reg_q2526 AND symb_decoder(16#3e#)) OR
 					(reg_q2526 AND symb_decoder(16#f8#)) OR
 					(reg_q2526 AND symb_decoder(16#16#)) OR
 					(reg_q2526 AND symb_decoder(16#06#)) OR
 					(reg_q2526 AND symb_decoder(16#f9#)) OR
 					(reg_q2526 AND symb_decoder(16#6b#)) OR
 					(reg_q2526 AND symb_decoder(16#01#)) OR
 					(reg_q2526 AND symb_decoder(16#0f#)) OR
 					(reg_q2526 AND symb_decoder(16#cb#)) OR
 					(reg_q2526 AND symb_decoder(16#47#)) OR
 					(reg_q2526 AND symb_decoder(16#dd#)) OR
 					(reg_q2526 AND symb_decoder(16#5f#)) OR
 					(reg_q2526 AND symb_decoder(16#e4#)) OR
 					(reg_q2526 AND symb_decoder(16#f4#)) OR
 					(reg_q2526 AND symb_decoder(16#d4#)) OR
 					(reg_q2526 AND symb_decoder(16#ec#)) OR
 					(reg_q2526 AND symb_decoder(16#e9#)) OR
 					(reg_q2526 AND symb_decoder(16#37#)) OR
 					(reg_q2526 AND symb_decoder(16#c4#)) OR
 					(reg_q2526 AND symb_decoder(16#d5#)) OR
 					(reg_q2526 AND symb_decoder(16#e3#)) OR
 					(reg_q2526 AND symb_decoder(16#4e#)) OR
 					(reg_q2526 AND symb_decoder(16#b3#)) OR
 					(reg_q2526 AND symb_decoder(16#b5#)) OR
 					(reg_q2526 AND symb_decoder(16#4b#)) OR
 					(reg_q2526 AND symb_decoder(16#15#)) OR
 					(reg_q2526 AND symb_decoder(16#fb#)) OR
 					(reg_q2526 AND symb_decoder(16#28#)) OR
 					(reg_q2526 AND symb_decoder(16#bf#)) OR
 					(reg_q2526 AND symb_decoder(16#1d#)) OR
 					(reg_q2526 AND symb_decoder(16#ad#)) OR
 					(reg_q2526 AND symb_decoder(16#19#)) OR
 					(reg_q2526 AND symb_decoder(16#7e#)) OR
 					(reg_q2526 AND symb_decoder(16#14#)) OR
 					(reg_q2526 AND symb_decoder(16#8a#)) OR
 					(reg_q2526 AND symb_decoder(16#9f#)) OR
 					(reg_q2526 AND symb_decoder(16#98#)) OR
 					(reg_q2526 AND symb_decoder(16#fd#)) OR
 					(reg_q2526 AND symb_decoder(16#e0#)) OR
 					(reg_q2526 AND symb_decoder(16#4f#)) OR
 					(reg_q2526 AND symb_decoder(16#5e#)) OR
 					(reg_q2526 AND symb_decoder(16#54#)) OR
 					(reg_q2526 AND symb_decoder(16#3d#)) OR
 					(reg_q2526 AND symb_decoder(16#c3#)) OR
 					(reg_q2526 AND symb_decoder(16#93#)) OR
 					(reg_q2526 AND symb_decoder(16#f5#)) OR
 					(reg_q2526 AND symb_decoder(16#0d#)) OR
 					(reg_q2526 AND symb_decoder(16#44#)) OR
 					(reg_q2526 AND symb_decoder(16#db#)) OR
 					(reg_q2526 AND symb_decoder(16#0e#)) OR
 					(reg_q2526 AND symb_decoder(16#87#)) OR
 					(reg_q2526 AND symb_decoder(16#de#)) OR
 					(reg_q2526 AND symb_decoder(16#67#)) OR
 					(reg_q2526 AND symb_decoder(16#64#)) OR
 					(reg_q2526 AND symb_decoder(16#ac#)) OR
 					(reg_q2526 AND symb_decoder(16#c9#)) OR
 					(reg_q2526 AND symb_decoder(16#2a#)) OR
 					(reg_q2526 AND symb_decoder(16#f1#)) OR
 					(reg_q2526 AND symb_decoder(16#fe#)) OR
 					(reg_q2526 AND symb_decoder(16#ed#)) OR
 					(reg_q2526 AND symb_decoder(16#05#)) OR
 					(reg_q2526 AND symb_decoder(16#cd#)) OR
 					(reg_q2526 AND symb_decoder(16#d0#)) OR
 					(reg_q2526 AND symb_decoder(16#29#)) OR
 					(reg_q2526 AND symb_decoder(16#2f#)) OR
 					(reg_q2526 AND symb_decoder(16#5d#)) OR
 					(reg_q2526 AND symb_decoder(16#a2#)) OR
 					(reg_q2526 AND symb_decoder(16#eb#)) OR
 					(reg_q2526 AND symb_decoder(16#41#)) OR
 					(reg_q2526 AND symb_decoder(16#63#)) OR
 					(reg_q2526 AND symb_decoder(16#75#)) OR
 					(reg_q2526 AND symb_decoder(16#5c#)) OR
 					(reg_q2526 AND symb_decoder(16#e5#)) OR
 					(reg_q2526 AND symb_decoder(16#da#)) OR
 					(reg_q2526 AND symb_decoder(16#13#)) OR
 					(reg_q2526 AND symb_decoder(16#b9#)) OR
 					(reg_q2526 AND symb_decoder(16#3f#)) OR
 					(reg_q2526 AND symb_decoder(16#9c#)) OR
 					(reg_q2526 AND symb_decoder(16#f3#)) OR
 					(reg_q2526 AND symb_decoder(16#ef#)) OR
 					(reg_q2526 AND symb_decoder(16#77#)) OR
 					(reg_q2526 AND symb_decoder(16#8c#)) OR
 					(reg_q2526 AND symb_decoder(16#04#)) OR
 					(reg_q2526 AND symb_decoder(16#e8#)) OR
 					(reg_q2526 AND symb_decoder(16#43#)) OR
 					(reg_q2526 AND symb_decoder(16#d9#)) OR
 					(reg_q2526 AND symb_decoder(16#56#)) OR
 					(reg_q2526 AND symb_decoder(16#8f#)) OR
 					(reg_q2526 AND symb_decoder(16#f6#)) OR
 					(reg_q2526 AND symb_decoder(16#7d#)) OR
 					(reg_q2526 AND symb_decoder(16#79#)) OR
 					(reg_q2526 AND symb_decoder(16#9b#)) OR
 					(reg_q2526 AND symb_decoder(16#e1#)) OR
 					(reg_q2526 AND symb_decoder(16#76#)) OR
 					(reg_q2526 AND symb_decoder(16#b8#)) OR
 					(reg_q2526 AND symb_decoder(16#ee#)) OR
 					(reg_q2526 AND symb_decoder(16#b1#)) OR
 					(reg_q2526 AND symb_decoder(16#72#)) OR
 					(reg_q2526 AND symb_decoder(16#55#)) OR
 					(reg_q2526 AND symb_decoder(16#80#)) OR
 					(reg_q2554 AND symb_decoder(16#33#)) OR
 					(reg_q2554 AND symb_decoder(16#77#)) OR
 					(reg_q2554 AND symb_decoder(16#6e#)) OR
 					(reg_q2554 AND symb_decoder(16#bc#)) OR
 					(reg_q2554 AND symb_decoder(16#7f#)) OR
 					(reg_q2554 AND symb_decoder(16#e4#)) OR
 					(reg_q2554 AND symb_decoder(16#5d#)) OR
 					(reg_q2554 AND symb_decoder(16#35#)) OR
 					(reg_q2554 AND symb_decoder(16#d5#)) OR
 					(reg_q2554 AND symb_decoder(16#27#)) OR
 					(reg_q2554 AND symb_decoder(16#2b#)) OR
 					(reg_q2554 AND symb_decoder(16#dd#)) OR
 					(reg_q2554 AND symb_decoder(16#ba#)) OR
 					(reg_q2554 AND symb_decoder(16#c9#)) OR
 					(reg_q2554 AND symb_decoder(16#c8#)) OR
 					(reg_q2554 AND symb_decoder(16#08#)) OR
 					(reg_q2554 AND symb_decoder(16#b6#)) OR
 					(reg_q2554 AND symb_decoder(16#85#)) OR
 					(reg_q2554 AND symb_decoder(16#f3#)) OR
 					(reg_q2554 AND symb_decoder(16#ec#)) OR
 					(reg_q2554 AND symb_decoder(16#20#)) OR
 					(reg_q2554 AND symb_decoder(16#83#)) OR
 					(reg_q2554 AND symb_decoder(16#fa#)) OR
 					(reg_q2554 AND symb_decoder(16#56#)) OR
 					(reg_q2554 AND symb_decoder(16#d4#)) OR
 					(reg_q2554 AND symb_decoder(16#21#)) OR
 					(reg_q2554 AND symb_decoder(16#29#)) OR
 					(reg_q2554 AND symb_decoder(16#88#)) OR
 					(reg_q2554 AND symb_decoder(16#81#)) OR
 					(reg_q2554 AND symb_decoder(16#1d#)) OR
 					(reg_q2554 AND symb_decoder(16#98#)) OR
 					(reg_q2554 AND symb_decoder(16#aa#)) OR
 					(reg_q2554 AND symb_decoder(16#af#)) OR
 					(reg_q2554 AND symb_decoder(16#10#)) OR
 					(reg_q2554 AND symb_decoder(16#9f#)) OR
 					(reg_q2554 AND symb_decoder(16#3d#)) OR
 					(reg_q2554 AND symb_decoder(16#06#)) OR
 					(reg_q2554 AND symb_decoder(16#97#)) OR
 					(reg_q2554 AND symb_decoder(16#05#)) OR
 					(reg_q2554 AND symb_decoder(16#5e#)) OR
 					(reg_q2554 AND symb_decoder(16#e5#)) OR
 					(reg_q2554 AND symb_decoder(16#5a#)) OR
 					(reg_q2554 AND symb_decoder(16#b8#)) OR
 					(reg_q2554 AND symb_decoder(16#64#)) OR
 					(reg_q2554 AND symb_decoder(16#50#)) OR
 					(reg_q2554 AND symb_decoder(16#69#)) OR
 					(reg_q2554 AND symb_decoder(16#1c#)) OR
 					(reg_q2554 AND symb_decoder(16#9d#)) OR
 					(reg_q2554 AND symb_decoder(16#c6#)) OR
 					(reg_q2554 AND symb_decoder(16#99#)) OR
 					(reg_q2554 AND symb_decoder(16#0b#)) OR
 					(reg_q2554 AND symb_decoder(16#cd#)) OR
 					(reg_q2554 AND symb_decoder(16#19#)) OR
 					(reg_q2554 AND symb_decoder(16#4c#)) OR
 					(reg_q2554 AND symb_decoder(16#c4#)) OR
 					(reg_q2554 AND symb_decoder(16#76#)) OR
 					(reg_q2554 AND symb_decoder(16#f7#)) OR
 					(reg_q2554 AND symb_decoder(16#45#)) OR
 					(reg_q2554 AND symb_decoder(16#86#)) OR
 					(reg_q2554 AND symb_decoder(16#30#)) OR
 					(reg_q2554 AND symb_decoder(16#d9#)) OR
 					(reg_q2554 AND symb_decoder(16#3f#)) OR
 					(reg_q2554 AND symb_decoder(16#f8#)) OR
 					(reg_q2554 AND symb_decoder(16#13#)) OR
 					(reg_q2554 AND symb_decoder(16#5b#)) OR
 					(reg_q2554 AND symb_decoder(16#41#)) OR
 					(reg_q2554 AND symb_decoder(16#1b#)) OR
 					(reg_q2554 AND symb_decoder(16#32#)) OR
 					(reg_q2554 AND symb_decoder(16#31#)) OR
 					(reg_q2554 AND symb_decoder(16#09#)) OR
 					(reg_q2554 AND symb_decoder(16#3e#)) OR
 					(reg_q2554 AND symb_decoder(16#18#)) OR
 					(reg_q2554 AND symb_decoder(16#e2#)) OR
 					(reg_q2554 AND symb_decoder(16#c5#)) OR
 					(reg_q2554 AND symb_decoder(16#59#)) OR
 					(reg_q2554 AND symb_decoder(16#4e#)) OR
 					(reg_q2554 AND symb_decoder(16#91#)) OR
 					(reg_q2554 AND symb_decoder(16#9e#)) OR
 					(reg_q2554 AND symb_decoder(16#da#)) OR
 					(reg_q2554 AND symb_decoder(16#04#)) OR
 					(reg_q2554 AND symb_decoder(16#dc#)) OR
 					(reg_q2554 AND symb_decoder(16#01#)) OR
 					(reg_q2554 AND symb_decoder(16#e6#)) OR
 					(reg_q2554 AND symb_decoder(16#d7#)) OR
 					(reg_q2554 AND symb_decoder(16#6a#)) OR
 					(reg_q2554 AND symb_decoder(16#6d#)) OR
 					(reg_q2554 AND symb_decoder(16#70#)) OR
 					(reg_q2554 AND symb_decoder(16#a6#)) OR
 					(reg_q2554 AND symb_decoder(16#fd#)) OR
 					(reg_q2554 AND symb_decoder(16#c2#)) OR
 					(reg_q2554 AND symb_decoder(16#b5#)) OR
 					(reg_q2554 AND symb_decoder(16#ea#)) OR
 					(reg_q2554 AND symb_decoder(16#46#)) OR
 					(reg_q2554 AND symb_decoder(16#e0#)) OR
 					(reg_q2554 AND symb_decoder(16#df#)) OR
 					(reg_q2554 AND symb_decoder(16#93#)) OR
 					(reg_q2554 AND symb_decoder(16#a2#)) OR
 					(reg_q2554 AND symb_decoder(16#17#)) OR
 					(reg_q2554 AND symb_decoder(16#94#)) OR
 					(reg_q2554 AND symb_decoder(16#ee#)) OR
 					(reg_q2554 AND symb_decoder(16#57#)) OR
 					(reg_q2554 AND symb_decoder(16#c7#)) OR
 					(reg_q2554 AND symb_decoder(16#90#)) OR
 					(reg_q2554 AND symb_decoder(16#82#)) OR
 					(reg_q2554 AND symb_decoder(16#bb#)) OR
 					(reg_q2554 AND symb_decoder(16#02#)) OR
 					(reg_q2554 AND symb_decoder(16#0c#)) OR
 					(reg_q2554 AND symb_decoder(16#3c#)) OR
 					(reg_q2554 AND symb_decoder(16#4b#)) OR
 					(reg_q2554 AND symb_decoder(16#e8#)) OR
 					(reg_q2554 AND symb_decoder(16#53#)) OR
 					(reg_q2554 AND symb_decoder(16#f4#)) OR
 					(reg_q2554 AND symb_decoder(16#63#)) OR
 					(reg_q2554 AND symb_decoder(16#b1#)) OR
 					(reg_q2554 AND symb_decoder(16#f1#)) OR
 					(reg_q2554 AND symb_decoder(16#75#)) OR
 					(reg_q2554 AND symb_decoder(16#58#)) OR
 					(reg_q2554 AND symb_decoder(16#a9#)) OR
 					(reg_q2554 AND symb_decoder(16#d6#)) OR
 					(reg_q2554 AND symb_decoder(16#96#)) OR
 					(reg_q2554 AND symb_decoder(16#1a#)) OR
 					(reg_q2554 AND symb_decoder(16#a5#)) OR
 					(reg_q2554 AND symb_decoder(16#bd#)) OR
 					(reg_q2554 AND symb_decoder(16#c3#)) OR
 					(reg_q2554 AND symb_decoder(16#de#)) OR
 					(reg_q2554 AND symb_decoder(16#66#)) OR
 					(reg_q2554 AND symb_decoder(16#cc#)) OR
 					(reg_q2554 AND symb_decoder(16#3b#)) OR
 					(reg_q2554 AND symb_decoder(16#47#)) OR
 					(reg_q2554 AND symb_decoder(16#1e#)) OR
 					(reg_q2554 AND symb_decoder(16#5f#)) OR
 					(reg_q2554 AND symb_decoder(16#f2#)) OR
 					(reg_q2554 AND symb_decoder(16#d2#)) OR
 					(reg_q2554 AND symb_decoder(16#7c#)) OR
 					(reg_q2554 AND symb_decoder(16#ae#)) OR
 					(reg_q2554 AND symb_decoder(16#a7#)) OR
 					(reg_q2554 AND symb_decoder(16#49#)) OR
 					(reg_q2554 AND symb_decoder(16#ff#)) OR
 					(reg_q2554 AND symb_decoder(16#11#)) OR
 					(reg_q2554 AND symb_decoder(16#ad#)) OR
 					(reg_q2554 AND symb_decoder(16#ca#)) OR
 					(reg_q2554 AND symb_decoder(16#b9#)) OR
 					(reg_q2554 AND symb_decoder(16#0a#)) OR
 					(reg_q2554 AND symb_decoder(16#f0#)) OR
 					(reg_q2554 AND symb_decoder(16#37#)) OR
 					(reg_q2554 AND symb_decoder(16#fc#)) OR
 					(reg_q2554 AND symb_decoder(16#d1#)) OR
 					(reg_q2554 AND symb_decoder(16#fe#)) OR
 					(reg_q2554 AND symb_decoder(16#8a#)) OR
 					(reg_q2554 AND symb_decoder(16#14#)) OR
 					(reg_q2554 AND symb_decoder(16#ce#)) OR
 					(reg_q2554 AND symb_decoder(16#d0#)) OR
 					(reg_q2554 AND symb_decoder(16#60#)) OR
 					(reg_q2554 AND symb_decoder(16#62#)) OR
 					(reg_q2554 AND symb_decoder(16#72#)) OR
 					(reg_q2554 AND symb_decoder(16#d3#)) OR
 					(reg_q2554 AND symb_decoder(16#b0#)) OR
 					(reg_q2554 AND symb_decoder(16#36#)) OR
 					(reg_q2554 AND symb_decoder(16#b2#)) OR
 					(reg_q2554 AND symb_decoder(16#2f#)) OR
 					(reg_q2554 AND symb_decoder(16#26#)) OR
 					(reg_q2554 AND symb_decoder(16#07#)) OR
 					(reg_q2554 AND symb_decoder(16#52#)) OR
 					(reg_q2554 AND symb_decoder(16#a1#)) OR
 					(reg_q2554 AND symb_decoder(16#95#)) OR
 					(reg_q2554 AND symb_decoder(16#bf#)) OR
 					(reg_q2554 AND symb_decoder(16#9c#)) OR
 					(reg_q2554 AND symb_decoder(16#22#)) OR
 					(reg_q2554 AND symb_decoder(16#78#)) OR
 					(reg_q2554 AND symb_decoder(16#e7#)) OR
 					(reg_q2554 AND symb_decoder(16#8d#)) OR
 					(reg_q2554 AND symb_decoder(16#79#)) OR
 					(reg_q2554 AND symb_decoder(16#7a#)) OR
 					(reg_q2554 AND symb_decoder(16#cb#)) OR
 					(reg_q2554 AND symb_decoder(16#be#)) OR
 					(reg_q2554 AND symb_decoder(16#7b#)) OR
 					(reg_q2554 AND symb_decoder(16#9a#)) OR
 					(reg_q2554 AND symb_decoder(16#34#)) OR
 					(reg_q2554 AND symb_decoder(16#84#)) OR
 					(reg_q2554 AND symb_decoder(16#65#)) OR
 					(reg_q2554 AND symb_decoder(16#6f#)) OR
 					(reg_q2554 AND symb_decoder(16#2a#)) OR
 					(reg_q2554 AND symb_decoder(16#89#)) OR
 					(reg_q2554 AND symb_decoder(16#23#)) OR
 					(reg_q2554 AND symb_decoder(16#03#)) OR
 					(reg_q2554 AND symb_decoder(16#a0#)) OR
 					(reg_q2554 AND symb_decoder(16#68#)) OR
 					(reg_q2554 AND symb_decoder(16#a4#)) OR
 					(reg_q2554 AND symb_decoder(16#15#)) OR
 					(reg_q2554 AND symb_decoder(16#6c#)) OR
 					(reg_q2554 AND symb_decoder(16#ab#)) OR
 					(reg_q2554 AND symb_decoder(16#2c#)) OR
 					(reg_q2554 AND symb_decoder(16#f9#)) OR
 					(reg_q2554 AND symb_decoder(16#54#)) OR
 					(reg_q2554 AND symb_decoder(16#9b#)) OR
 					(reg_q2554 AND symb_decoder(16#ef#)) OR
 					(reg_q2554 AND symb_decoder(16#25#)) OR
 					(reg_q2554 AND symb_decoder(16#e1#)) OR
 					(reg_q2554 AND symb_decoder(16#4a#)) OR
 					(reg_q2554 AND symb_decoder(16#e3#)) OR
 					(reg_q2554 AND symb_decoder(16#2e#)) OR
 					(reg_q2554 AND symb_decoder(16#5c#)) OR
 					(reg_q2554 AND symb_decoder(16#43#)) OR
 					(reg_q2554 AND symb_decoder(16#c0#)) OR
 					(reg_q2554 AND symb_decoder(16#b3#)) OR
 					(reg_q2554 AND symb_decoder(16#48#)) OR
 					(reg_q2554 AND symb_decoder(16#f6#)) OR
 					(reg_q2554 AND symb_decoder(16#92#)) OR
 					(reg_q2554 AND symb_decoder(16#7d#)) OR
 					(reg_q2554 AND symb_decoder(16#16#)) OR
 					(reg_q2554 AND symb_decoder(16#38#)) OR
 					(reg_q2554 AND symb_decoder(16#80#)) OR
 					(reg_q2554 AND symb_decoder(16#4d#)) OR
 					(reg_q2554 AND symb_decoder(16#eb#)) OR
 					(reg_q2554 AND symb_decoder(16#8e#)) OR
 					(reg_q2554 AND symb_decoder(16#a3#)) OR
 					(reg_q2554 AND symb_decoder(16#44#)) OR
 					(reg_q2554 AND symb_decoder(16#00#)) OR
 					(reg_q2554 AND symb_decoder(16#55#)) OR
 					(reg_q2554 AND symb_decoder(16#ed#)) OR
 					(reg_q2554 AND symb_decoder(16#7e#)) OR
 					(reg_q2554 AND symb_decoder(16#1f#)) OR
 					(reg_q2554 AND symb_decoder(16#db#)) OR
 					(reg_q2554 AND symb_decoder(16#a8#)) OR
 					(reg_q2554 AND symb_decoder(16#42#)) OR
 					(reg_q2554 AND symb_decoder(16#39#)) OR
 					(reg_q2554 AND symb_decoder(16#4f#)) OR
 					(reg_q2554 AND symb_decoder(16#8b#)) OR
 					(reg_q2554 AND symb_decoder(16#ac#)) OR
 					(reg_q2554 AND symb_decoder(16#40#)) OR
 					(reg_q2554 AND symb_decoder(16#8f#)) OR
 					(reg_q2554 AND symb_decoder(16#0e#)) OR
 					(reg_q2554 AND symb_decoder(16#61#)) OR
 					(reg_q2554 AND symb_decoder(16#87#)) OR
 					(reg_q2554 AND symb_decoder(16#cf#)) OR
 					(reg_q2554 AND symb_decoder(16#e9#)) OR
 					(reg_q2554 AND symb_decoder(16#b7#)) OR
 					(reg_q2554 AND symb_decoder(16#71#)) OR
 					(reg_q2554 AND symb_decoder(16#c1#)) OR
 					(reg_q2554 AND symb_decoder(16#6b#)) OR
 					(reg_q2554 AND symb_decoder(16#2d#)) OR
 					(reg_q2554 AND symb_decoder(16#0f#)) OR
 					(reg_q2554 AND symb_decoder(16#24#)) OR
 					(reg_q2554 AND symb_decoder(16#8c#)) OR
 					(reg_q2554 AND symb_decoder(16#f5#)) OR
 					(reg_q2554 AND symb_decoder(16#12#)) OR
 					(reg_q2554 AND symb_decoder(16#73#)) OR
 					(reg_q2554 AND symb_decoder(16#67#)) OR
 					(reg_q2554 AND symb_decoder(16#fb#)) OR
 					(reg_q2554 AND symb_decoder(16#0d#)) OR
 					(reg_q2554 AND symb_decoder(16#51#)) OR
 					(reg_q2554 AND symb_decoder(16#28#)) OR
 					(reg_q2554 AND symb_decoder(16#b4#)) OR
 					(reg_q2554 AND symb_decoder(16#d8#)) OR
 					(reg_q2554 AND symb_decoder(16#3a#)) OR
 					(reg_q2554 AND symb_decoder(16#74#));
reg_q2554_init <= '0' ;
	p_reg_q2554: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2554 <= reg_q2554_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2554 <= reg_q2554_init;
        else
          reg_q2554 <= reg_q2554_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1479_in <= (reg_q1479 AND symb_decoder(16#2a#)) OR
 					(reg_q1479 AND symb_decoder(16#7e#)) OR
 					(reg_q1479 AND symb_decoder(16#50#)) OR
 					(reg_q1479 AND symb_decoder(16#5a#)) OR
 					(reg_q1479 AND symb_decoder(16#3e#)) OR
 					(reg_q1479 AND symb_decoder(16#9d#)) OR
 					(reg_q1479 AND symb_decoder(16#8b#)) OR
 					(reg_q1479 AND symb_decoder(16#f6#)) OR
 					(reg_q1479 AND symb_decoder(16#bd#)) OR
 					(reg_q1479 AND symb_decoder(16#f2#)) OR
 					(reg_q1479 AND symb_decoder(16#12#)) OR
 					(reg_q1479 AND symb_decoder(16#ea#)) OR
 					(reg_q1479 AND symb_decoder(16#0c#)) OR
 					(reg_q1479 AND symb_decoder(16#02#)) OR
 					(reg_q1479 AND symb_decoder(16#70#)) OR
 					(reg_q1479 AND symb_decoder(16#33#)) OR
 					(reg_q1479 AND symb_decoder(16#d5#)) OR
 					(reg_q1479 AND symb_decoder(16#4a#)) OR
 					(reg_q1479 AND symb_decoder(16#63#)) OR
 					(reg_q1479 AND symb_decoder(16#bf#)) OR
 					(reg_q1479 AND symb_decoder(16#7d#)) OR
 					(reg_q1479 AND symb_decoder(16#84#)) OR
 					(reg_q1479 AND symb_decoder(16#41#)) OR
 					(reg_q1479 AND symb_decoder(16#30#)) OR
 					(reg_q1479 AND symb_decoder(16#74#)) OR
 					(reg_q1479 AND symb_decoder(16#96#)) OR
 					(reg_q1479 AND symb_decoder(16#3a#)) OR
 					(reg_q1479 AND symb_decoder(16#f3#)) OR
 					(reg_q1479 AND symb_decoder(16#89#)) OR
 					(reg_q1479 AND symb_decoder(16#e5#)) OR
 					(reg_q1479 AND symb_decoder(16#26#)) OR
 					(reg_q1479 AND symb_decoder(16#b2#)) OR
 					(reg_q1479 AND symb_decoder(16#c7#)) OR
 					(reg_q1479 AND symb_decoder(16#a4#)) OR
 					(reg_q1479 AND symb_decoder(16#1d#)) OR
 					(reg_q1479 AND symb_decoder(16#2c#)) OR
 					(reg_q1479 AND symb_decoder(16#06#)) OR
 					(reg_q1479 AND symb_decoder(16#58#)) OR
 					(reg_q1479 AND symb_decoder(16#91#)) OR
 					(reg_q1479 AND symb_decoder(16#a5#)) OR
 					(reg_q1479 AND symb_decoder(16#04#)) OR
 					(reg_q1479 AND symb_decoder(16#0a#)) OR
 					(reg_q1479 AND symb_decoder(16#52#)) OR
 					(reg_q1479 AND symb_decoder(16#e3#)) OR
 					(reg_q1479 AND symb_decoder(16#e1#)) OR
 					(reg_q1479 AND symb_decoder(16#35#)) OR
 					(reg_q1479 AND symb_decoder(16#dd#)) OR
 					(reg_q1479 AND symb_decoder(16#93#)) OR
 					(reg_q1479 AND symb_decoder(16#32#)) OR
 					(reg_q1479 AND symb_decoder(16#a3#)) OR
 					(reg_q1479 AND symb_decoder(16#2b#)) OR
 					(reg_q1479 AND symb_decoder(16#1c#)) OR
 					(reg_q1479 AND symb_decoder(16#e0#)) OR
 					(reg_q1479 AND symb_decoder(16#ba#)) OR
 					(reg_q1479 AND symb_decoder(16#a7#)) OR
 					(reg_q1479 AND symb_decoder(16#ee#)) OR
 					(reg_q1479 AND symb_decoder(16#6e#)) OR
 					(reg_q1479 AND symb_decoder(16#40#)) OR
 					(reg_q1479 AND symb_decoder(16#99#)) OR
 					(reg_q1479 AND symb_decoder(16#d6#)) OR
 					(reg_q1479 AND symb_decoder(16#94#)) OR
 					(reg_q1479 AND symb_decoder(16#5f#)) OR
 					(reg_q1479 AND symb_decoder(16#34#)) OR
 					(reg_q1479 AND symb_decoder(16#59#)) OR
 					(reg_q1479 AND symb_decoder(16#e2#)) OR
 					(reg_q1479 AND symb_decoder(16#f5#)) OR
 					(reg_q1479 AND symb_decoder(16#46#)) OR
 					(reg_q1479 AND symb_decoder(16#66#)) OR
 					(reg_q1479 AND symb_decoder(16#19#)) OR
 					(reg_q1479 AND symb_decoder(16#11#)) OR
 					(reg_q1479 AND symb_decoder(16#86#)) OR
 					(reg_q1479 AND symb_decoder(16#03#)) OR
 					(reg_q1479 AND symb_decoder(16#54#)) OR
 					(reg_q1479 AND symb_decoder(16#15#)) OR
 					(reg_q1479 AND symb_decoder(16#36#)) OR
 					(reg_q1479 AND symb_decoder(16#56#)) OR
 					(reg_q1479 AND symb_decoder(16#76#)) OR
 					(reg_q1479 AND symb_decoder(16#a1#)) OR
 					(reg_q1479 AND symb_decoder(16#c2#)) OR
 					(reg_q1479 AND symb_decoder(16#97#)) OR
 					(reg_q1479 AND symb_decoder(16#49#)) OR
 					(reg_q1479 AND symb_decoder(16#53#)) OR
 					(reg_q1479 AND symb_decoder(16#e6#)) OR
 					(reg_q1479 AND symb_decoder(16#43#)) OR
 					(reg_q1479 AND symb_decoder(16#fd#)) OR
 					(reg_q1479 AND symb_decoder(16#20#)) OR
 					(reg_q1479 AND symb_decoder(16#c4#)) OR
 					(reg_q1479 AND symb_decoder(16#ce#)) OR
 					(reg_q1479 AND symb_decoder(16#bb#)) OR
 					(reg_q1479 AND symb_decoder(16#29#)) OR
 					(reg_q1479 AND symb_decoder(16#98#)) OR
 					(reg_q1479 AND symb_decoder(16#95#)) OR
 					(reg_q1479 AND symb_decoder(16#a6#)) OR
 					(reg_q1479 AND symb_decoder(16#b8#)) OR
 					(reg_q1479 AND symb_decoder(16#8d#)) OR
 					(reg_q1479 AND symb_decoder(16#cd#)) OR
 					(reg_q1479 AND symb_decoder(16#fa#)) OR
 					(reg_q1479 AND symb_decoder(16#c3#)) OR
 					(reg_q1479 AND symb_decoder(16#d1#)) OR
 					(reg_q1479 AND symb_decoder(16#b7#)) OR
 					(reg_q1479 AND symb_decoder(16#7a#)) OR
 					(reg_q1479 AND symb_decoder(16#39#)) OR
 					(reg_q1479 AND symb_decoder(16#6c#)) OR
 					(reg_q1479 AND symb_decoder(16#08#)) OR
 					(reg_q1479 AND symb_decoder(16#2f#)) OR
 					(reg_q1479 AND symb_decoder(16#af#)) OR
 					(reg_q1479 AND symb_decoder(16#83#)) OR
 					(reg_q1479 AND symb_decoder(16#a9#)) OR
 					(reg_q1479 AND symb_decoder(16#dc#)) OR
 					(reg_q1479 AND symb_decoder(16#f1#)) OR
 					(reg_q1479 AND symb_decoder(16#2e#)) OR
 					(reg_q1479 AND symb_decoder(16#77#)) OR
 					(reg_q1479 AND symb_decoder(16#87#)) OR
 					(reg_q1479 AND symb_decoder(16#60#)) OR
 					(reg_q1479 AND symb_decoder(16#85#)) OR
 					(reg_q1479 AND symb_decoder(16#9a#)) OR
 					(reg_q1479 AND symb_decoder(16#7c#)) OR
 					(reg_q1479 AND symb_decoder(16#d8#)) OR
 					(reg_q1479 AND symb_decoder(16#a2#)) OR
 					(reg_q1479 AND symb_decoder(16#64#)) OR
 					(reg_q1479 AND symb_decoder(16#2d#)) OR
 					(reg_q1479 AND symb_decoder(16#e7#)) OR
 					(reg_q1479 AND symb_decoder(16#0b#)) OR
 					(reg_q1479 AND symb_decoder(16#c0#)) OR
 					(reg_q1479 AND symb_decoder(16#ff#)) OR
 					(reg_q1479 AND symb_decoder(16#24#)) OR
 					(reg_q1479 AND symb_decoder(16#5d#)) OR
 					(reg_q1479 AND symb_decoder(16#1b#)) OR
 					(reg_q1479 AND symb_decoder(16#c1#)) OR
 					(reg_q1479 AND symb_decoder(16#4f#)) OR
 					(reg_q1479 AND symb_decoder(16#6f#)) OR
 					(reg_q1479 AND symb_decoder(16#5c#)) OR
 					(reg_q1479 AND symb_decoder(16#f7#)) OR
 					(reg_q1479 AND symb_decoder(16#38#)) OR
 					(reg_q1479 AND symb_decoder(16#61#)) OR
 					(reg_q1479 AND symb_decoder(16#b3#)) OR
 					(reg_q1479 AND symb_decoder(16#62#)) OR
 					(reg_q1479 AND symb_decoder(16#b9#)) OR
 					(reg_q1479 AND symb_decoder(16#f4#)) OR
 					(reg_q1479 AND symb_decoder(16#16#)) OR
 					(reg_q1479 AND symb_decoder(16#8f#)) OR
 					(reg_q1479 AND symb_decoder(16#c8#)) OR
 					(reg_q1479 AND symb_decoder(16#0d#)) OR
 					(reg_q1479 AND symb_decoder(16#e4#)) OR
 					(reg_q1479 AND symb_decoder(16#0e#)) OR
 					(reg_q1479 AND symb_decoder(16#cb#)) OR
 					(reg_q1479 AND symb_decoder(16#13#)) OR
 					(reg_q1479 AND symb_decoder(16#57#)) OR
 					(reg_q1479 AND symb_decoder(16#ec#)) OR
 					(reg_q1479 AND symb_decoder(16#4d#)) OR
 					(reg_q1479 AND symb_decoder(16#1f#)) OR
 					(reg_q1479 AND symb_decoder(16#3b#)) OR
 					(reg_q1479 AND symb_decoder(16#5b#)) OR
 					(reg_q1479 AND symb_decoder(16#bc#)) OR
 					(reg_q1479 AND symb_decoder(16#be#)) OR
 					(reg_q1479 AND symb_decoder(16#ef#)) OR
 					(reg_q1479 AND symb_decoder(16#37#)) OR
 					(reg_q1479 AND symb_decoder(16#de#)) OR
 					(reg_q1479 AND symb_decoder(16#df#)) OR
 					(reg_q1479 AND symb_decoder(16#9c#)) OR
 					(reg_q1479 AND symb_decoder(16#b5#)) OR
 					(reg_q1479 AND symb_decoder(16#e9#)) OR
 					(reg_q1479 AND symb_decoder(16#d9#)) OR
 					(reg_q1479 AND symb_decoder(16#45#)) OR
 					(reg_q1479 AND symb_decoder(16#cc#)) OR
 					(reg_q1479 AND symb_decoder(16#31#)) OR
 					(reg_q1479 AND symb_decoder(16#68#)) OR
 					(reg_q1479 AND symb_decoder(16#78#)) OR
 					(reg_q1479 AND symb_decoder(16#ed#)) OR
 					(reg_q1479 AND symb_decoder(16#d0#)) OR
 					(reg_q1479 AND symb_decoder(16#27#)) OR
 					(reg_q1479 AND symb_decoder(16#c5#)) OR
 					(reg_q1479 AND symb_decoder(16#47#)) OR
 					(reg_q1479 AND symb_decoder(16#cf#)) OR
 					(reg_q1479 AND symb_decoder(16#d2#)) OR
 					(reg_q1479 AND symb_decoder(16#6b#)) OR
 					(reg_q1479 AND symb_decoder(16#01#)) OR
 					(reg_q1479 AND symb_decoder(16#ca#)) OR
 					(reg_q1479 AND symb_decoder(16#4e#)) OR
 					(reg_q1479 AND symb_decoder(16#b6#)) OR
 					(reg_q1479 AND symb_decoder(16#6d#)) OR
 					(reg_q1479 AND symb_decoder(16#10#)) OR
 					(reg_q1479 AND symb_decoder(16#44#)) OR
 					(reg_q1479 AND symb_decoder(16#79#)) OR
 					(reg_q1479 AND symb_decoder(16#3d#)) OR
 					(reg_q1479 AND symb_decoder(16#c6#)) OR
 					(reg_q1479 AND symb_decoder(16#80#)) OR
 					(reg_q1479 AND symb_decoder(16#d7#)) OR
 					(reg_q1479 AND symb_decoder(16#1a#)) OR
 					(reg_q1479 AND symb_decoder(16#b1#)) OR
 					(reg_q1479 AND symb_decoder(16#7f#)) OR
 					(reg_q1479 AND symb_decoder(16#73#)) OR
 					(reg_q1479 AND symb_decoder(16#d4#)) OR
 					(reg_q1479 AND symb_decoder(16#17#)) OR
 					(reg_q1479 AND symb_decoder(16#b4#)) OR
 					(reg_q1479 AND symb_decoder(16#00#)) OR
 					(reg_q1479 AND symb_decoder(16#18#)) OR
 					(reg_q1479 AND symb_decoder(16#71#)) OR
 					(reg_q1479 AND symb_decoder(16#21#)) OR
 					(reg_q1479 AND symb_decoder(16#07#)) OR
 					(reg_q1479 AND symb_decoder(16#6a#)) OR
 					(reg_q1479 AND symb_decoder(16#f8#)) OR
 					(reg_q1479 AND symb_decoder(16#1e#)) OR
 					(reg_q1479 AND symb_decoder(16#8e#)) OR
 					(reg_q1479 AND symb_decoder(16#fe#)) OR
 					(reg_q1479 AND symb_decoder(16#eb#)) OR
 					(reg_q1479 AND symb_decoder(16#8c#)) OR
 					(reg_q1479 AND symb_decoder(16#05#)) OR
 					(reg_q1479 AND symb_decoder(16#0f#)) OR
 					(reg_q1479 AND symb_decoder(16#c9#)) OR
 					(reg_q1479 AND symb_decoder(16#a8#)) OR
 					(reg_q1479 AND symb_decoder(16#48#)) OR
 					(reg_q1479 AND symb_decoder(16#75#)) OR
 					(reg_q1479 AND symb_decoder(16#fb#)) OR
 					(reg_q1479 AND symb_decoder(16#67#)) OR
 					(reg_q1479 AND symb_decoder(16#aa#)) OR
 					(reg_q1479 AND symb_decoder(16#ae#)) OR
 					(reg_q1479 AND symb_decoder(16#65#)) OR
 					(reg_q1479 AND symb_decoder(16#8a#)) OR
 					(reg_q1479 AND symb_decoder(16#4c#)) OR
 					(reg_q1479 AND symb_decoder(16#28#)) OR
 					(reg_q1479 AND symb_decoder(16#69#)) OR
 					(reg_q1479 AND symb_decoder(16#7b#)) OR
 					(reg_q1479 AND symb_decoder(16#3c#)) OR
 					(reg_q1479 AND symb_decoder(16#da#)) OR
 					(reg_q1479 AND symb_decoder(16#3f#)) OR
 					(reg_q1479 AND symb_decoder(16#51#)) OR
 					(reg_q1479 AND symb_decoder(16#4b#)) OR
 					(reg_q1479 AND symb_decoder(16#fc#)) OR
 					(reg_q1479 AND symb_decoder(16#f0#)) OR
 					(reg_q1479 AND symb_decoder(16#f9#)) OR
 					(reg_q1479 AND symb_decoder(16#81#)) OR
 					(reg_q1479 AND symb_decoder(16#82#)) OR
 					(reg_q1479 AND symb_decoder(16#88#)) OR
 					(reg_q1479 AND symb_decoder(16#09#)) OR
 					(reg_q1479 AND symb_decoder(16#9f#)) OR
 					(reg_q1479 AND symb_decoder(16#55#)) OR
 					(reg_q1479 AND symb_decoder(16#ac#)) OR
 					(reg_q1479 AND symb_decoder(16#ab#)) OR
 					(reg_q1479 AND symb_decoder(16#b0#)) OR
 					(reg_q1479 AND symb_decoder(16#db#)) OR
 					(reg_q1479 AND symb_decoder(16#9b#)) OR
 					(reg_q1479 AND symb_decoder(16#22#)) OR
 					(reg_q1479 AND symb_decoder(16#23#)) OR
 					(reg_q1479 AND symb_decoder(16#42#)) OR
 					(reg_q1479 AND symb_decoder(16#d3#)) OR
 					(reg_q1479 AND symb_decoder(16#5e#)) OR
 					(reg_q1479 AND symb_decoder(16#92#)) OR
 					(reg_q1479 AND symb_decoder(16#72#)) OR
 					(reg_q1479 AND symb_decoder(16#e8#)) OR
 					(reg_q1479 AND symb_decoder(16#25#)) OR
 					(reg_q1479 AND symb_decoder(16#9e#)) OR
 					(reg_q1479 AND symb_decoder(16#ad#)) OR
 					(reg_q1479 AND symb_decoder(16#90#)) OR
 					(reg_q1479 AND symb_decoder(16#a0#)) OR
 					(reg_q1479 AND symb_decoder(16#14#)) OR
 					(reg_q1443 AND symb_decoder(16#38#)) OR
 					(reg_q1443 AND symb_decoder(16#6a#)) OR
 					(reg_q1443 AND symb_decoder(16#ec#)) OR
 					(reg_q1443 AND symb_decoder(16#5c#)) OR
 					(reg_q1443 AND symb_decoder(16#a5#)) OR
 					(reg_q1443 AND symb_decoder(16#09#)) OR
 					(reg_q1443 AND symb_decoder(16#f6#)) OR
 					(reg_q1443 AND symb_decoder(16#8b#)) OR
 					(reg_q1443 AND symb_decoder(16#41#)) OR
 					(reg_q1443 AND symb_decoder(16#8f#)) OR
 					(reg_q1443 AND symb_decoder(16#71#)) OR
 					(reg_q1443 AND symb_decoder(16#a7#)) OR
 					(reg_q1443 AND symb_decoder(16#6d#)) OR
 					(reg_q1443 AND symb_decoder(16#39#)) OR
 					(reg_q1443 AND symb_decoder(16#ad#)) OR
 					(reg_q1443 AND symb_decoder(16#83#)) OR
 					(reg_q1443 AND symb_decoder(16#b3#)) OR
 					(reg_q1443 AND symb_decoder(16#5b#)) OR
 					(reg_q1443 AND symb_decoder(16#ce#)) OR
 					(reg_q1443 AND symb_decoder(16#e7#)) OR
 					(reg_q1443 AND symb_decoder(16#8a#)) OR
 					(reg_q1443 AND symb_decoder(16#04#)) OR
 					(reg_q1443 AND symb_decoder(16#d9#)) OR
 					(reg_q1443 AND symb_decoder(16#5a#)) OR
 					(reg_q1443 AND symb_decoder(16#fb#)) OR
 					(reg_q1443 AND symb_decoder(16#52#)) OR
 					(reg_q1443 AND symb_decoder(16#a6#)) OR
 					(reg_q1443 AND symb_decoder(16#e9#)) OR
 					(reg_q1443 AND symb_decoder(16#df#)) OR
 					(reg_q1443 AND symb_decoder(16#d6#)) OR
 					(reg_q1443 AND symb_decoder(16#81#)) OR
 					(reg_q1443 AND symb_decoder(16#e5#)) OR
 					(reg_q1443 AND symb_decoder(16#4f#)) OR
 					(reg_q1443 AND symb_decoder(16#eb#)) OR
 					(reg_q1443 AND symb_decoder(16#29#)) OR
 					(reg_q1443 AND symb_decoder(16#9a#)) OR
 					(reg_q1443 AND symb_decoder(16#bb#)) OR
 					(reg_q1443 AND symb_decoder(16#af#)) OR
 					(reg_q1443 AND symb_decoder(16#e2#)) OR
 					(reg_q1443 AND symb_decoder(16#00#)) OR
 					(reg_q1443 AND symb_decoder(16#19#)) OR
 					(reg_q1443 AND symb_decoder(16#89#)) OR
 					(reg_q1443 AND symb_decoder(16#01#)) OR
 					(reg_q1443 AND symb_decoder(16#77#)) OR
 					(reg_q1443 AND symb_decoder(16#c2#)) OR
 					(reg_q1443 AND symb_decoder(16#9b#)) OR
 					(reg_q1443 AND symb_decoder(16#f3#)) OR
 					(reg_q1443 AND symb_decoder(16#db#)) OR
 					(reg_q1443 AND symb_decoder(16#17#)) OR
 					(reg_q1443 AND symb_decoder(16#46#)) OR
 					(reg_q1443 AND symb_decoder(16#1d#)) OR
 					(reg_q1443 AND symb_decoder(16#34#)) OR
 					(reg_q1443 AND symb_decoder(16#a3#)) OR
 					(reg_q1443 AND symb_decoder(16#82#)) OR
 					(reg_q1443 AND symb_decoder(16#e1#)) OR
 					(reg_q1443 AND symb_decoder(16#d5#)) OR
 					(reg_q1443 AND symb_decoder(16#1a#)) OR
 					(reg_q1443 AND symb_decoder(16#d8#)) OR
 					(reg_q1443 AND symb_decoder(16#be#)) OR
 					(reg_q1443 AND symb_decoder(16#fa#)) OR
 					(reg_q1443 AND symb_decoder(16#53#)) OR
 					(reg_q1443 AND symb_decoder(16#2b#)) OR
 					(reg_q1443 AND symb_decoder(16#57#)) OR
 					(reg_q1443 AND symb_decoder(16#8c#)) OR
 					(reg_q1443 AND symb_decoder(16#b8#)) OR
 					(reg_q1443 AND symb_decoder(16#0e#)) OR
 					(reg_q1443 AND symb_decoder(16#99#)) OR
 					(reg_q1443 AND symb_decoder(16#20#)) OR
 					(reg_q1443 AND symb_decoder(16#68#)) OR
 					(reg_q1443 AND symb_decoder(16#3a#)) OR
 					(reg_q1443 AND symb_decoder(16#dc#)) OR
 					(reg_q1443 AND symb_decoder(16#73#)) OR
 					(reg_q1443 AND symb_decoder(16#18#)) OR
 					(reg_q1443 AND symb_decoder(16#32#)) OR
 					(reg_q1443 AND symb_decoder(16#da#)) OR
 					(reg_q1443 AND symb_decoder(16#8d#)) OR
 					(reg_q1443 AND symb_decoder(16#b4#)) OR
 					(reg_q1443 AND symb_decoder(16#88#)) OR
 					(reg_q1443 AND symb_decoder(16#9f#)) OR
 					(reg_q1443 AND symb_decoder(16#94#)) OR
 					(reg_q1443 AND symb_decoder(16#7a#)) OR
 					(reg_q1443 AND symb_decoder(16#35#)) OR
 					(reg_q1443 AND symb_decoder(16#40#)) OR
 					(reg_q1443 AND symb_decoder(16#44#)) OR
 					(reg_q1443 AND symb_decoder(16#74#)) OR
 					(reg_q1443 AND symb_decoder(16#fd#)) OR
 					(reg_q1443 AND symb_decoder(16#63#)) OR
 					(reg_q1443 AND symb_decoder(16#37#)) OR
 					(reg_q1443 AND symb_decoder(16#c1#)) OR
 					(reg_q1443 AND symb_decoder(16#47#)) OR
 					(reg_q1443 AND symb_decoder(16#cd#)) OR
 					(reg_q1443 AND symb_decoder(16#f5#)) OR
 					(reg_q1443 AND symb_decoder(16#3b#)) OR
 					(reg_q1443 AND symb_decoder(16#d0#)) OR
 					(reg_q1443 AND symb_decoder(16#07#)) OR
 					(reg_q1443 AND symb_decoder(16#70#)) OR
 					(reg_q1443 AND symb_decoder(16#cc#)) OR
 					(reg_q1443 AND symb_decoder(16#43#)) OR
 					(reg_q1443 AND symb_decoder(16#f8#)) OR
 					(reg_q1443 AND symb_decoder(16#31#)) OR
 					(reg_q1443 AND symb_decoder(16#10#)) OR
 					(reg_q1443 AND symb_decoder(16#7c#)) OR
 					(reg_q1443 AND symb_decoder(16#30#)) OR
 					(reg_q1443 AND symb_decoder(16#b7#)) OR
 					(reg_q1443 AND symb_decoder(16#f0#)) OR
 					(reg_q1443 AND symb_decoder(16#c6#)) OR
 					(reg_q1443 AND symb_decoder(16#2c#)) OR
 					(reg_q1443 AND symb_decoder(16#33#)) OR
 					(reg_q1443 AND symb_decoder(16#03#)) OR
 					(reg_q1443 AND symb_decoder(16#78#)) OR
 					(reg_q1443 AND symb_decoder(16#ab#)) OR
 					(reg_q1443 AND symb_decoder(16#69#)) OR
 					(reg_q1443 AND symb_decoder(16#5f#)) OR
 					(reg_q1443 AND symb_decoder(16#87#)) OR
 					(reg_q1443 AND symb_decoder(16#a9#)) OR
 					(reg_q1443 AND symb_decoder(16#d7#)) OR
 					(reg_q1443 AND symb_decoder(16#6e#)) OR
 					(reg_q1443 AND symb_decoder(16#5d#)) OR
 					(reg_q1443 AND symb_decoder(16#96#)) OR
 					(reg_q1443 AND symb_decoder(16#ac#)) OR
 					(reg_q1443 AND symb_decoder(16#b9#)) OR
 					(reg_q1443 AND symb_decoder(16#2e#)) OR
 					(reg_q1443 AND symb_decoder(16#9c#)) OR
 					(reg_q1443 AND symb_decoder(16#f1#)) OR
 					(reg_q1443 AND symb_decoder(16#4e#)) OR
 					(reg_q1443 AND symb_decoder(16#b5#)) OR
 					(reg_q1443 AND symb_decoder(16#a2#)) OR
 					(reg_q1443 AND symb_decoder(16#22#)) OR
 					(reg_q1443 AND symb_decoder(16#13#)) OR
 					(reg_q1443 AND symb_decoder(16#93#)) OR
 					(reg_q1443 AND symb_decoder(16#d2#)) OR
 					(reg_q1443 AND symb_decoder(16#0a#)) OR
 					(reg_q1443 AND symb_decoder(16#24#)) OR
 					(reg_q1443 AND symb_decoder(16#95#)) OR
 					(reg_q1443 AND symb_decoder(16#ea#)) OR
 					(reg_q1443 AND symb_decoder(16#21#)) OR
 					(reg_q1443 AND symb_decoder(16#7e#)) OR
 					(reg_q1443 AND symb_decoder(16#3d#)) OR
 					(reg_q1443 AND symb_decoder(16#60#)) OR
 					(reg_q1443 AND symb_decoder(16#55#)) OR
 					(reg_q1443 AND symb_decoder(16#97#)) OR
 					(reg_q1443 AND symb_decoder(16#e6#)) OR
 					(reg_q1443 AND symb_decoder(16#ed#)) OR
 					(reg_q1443 AND symb_decoder(16#11#)) OR
 					(reg_q1443 AND symb_decoder(16#25#)) OR
 					(reg_q1443 AND symb_decoder(16#50#)) OR
 					(reg_q1443 AND symb_decoder(16#6c#)) OR
 					(reg_q1443 AND symb_decoder(16#62#)) OR
 					(reg_q1443 AND symb_decoder(16#76#)) OR
 					(reg_q1443 AND symb_decoder(16#51#)) OR
 					(reg_q1443 AND symb_decoder(16#90#)) OR
 					(reg_q1443 AND symb_decoder(16#cb#)) OR
 					(reg_q1443 AND symb_decoder(16#3e#)) OR
 					(reg_q1443 AND symb_decoder(16#ee#)) OR
 					(reg_q1443 AND symb_decoder(16#e0#)) OR
 					(reg_q1443 AND symb_decoder(16#54#)) OR
 					(reg_q1443 AND symb_decoder(16#02#)) OR
 					(reg_q1443 AND symb_decoder(16#66#)) OR
 					(reg_q1443 AND symb_decoder(16#d1#)) OR
 					(reg_q1443 AND symb_decoder(16#d4#)) OR
 					(reg_q1443 AND symb_decoder(16#4a#)) OR
 					(reg_q1443 AND symb_decoder(16#65#)) OR
 					(reg_q1443 AND symb_decoder(16#e4#)) OR
 					(reg_q1443 AND symb_decoder(16#d3#)) OR
 					(reg_q1443 AND symb_decoder(16#bd#)) OR
 					(reg_q1443 AND symb_decoder(16#e8#)) OR
 					(reg_q1443 AND symb_decoder(16#b1#)) OR
 					(reg_q1443 AND symb_decoder(16#85#)) OR
 					(reg_q1443 AND symb_decoder(16#8e#)) OR
 					(reg_q1443 AND symb_decoder(16#86#)) OR
 					(reg_q1443 AND symb_decoder(16#5e#)) OR
 					(reg_q1443 AND symb_decoder(16#80#)) OR
 					(reg_q1443 AND symb_decoder(16#dd#)) OR
 					(reg_q1443 AND symb_decoder(16#4b#)) OR
 					(reg_q1443 AND symb_decoder(16#ca#)) OR
 					(reg_q1443 AND symb_decoder(16#75#)) OR
 					(reg_q1443 AND symb_decoder(16#2a#)) OR
 					(reg_q1443 AND symb_decoder(16#7b#)) OR
 					(reg_q1443 AND symb_decoder(16#9e#)) OR
 					(reg_q1443 AND symb_decoder(16#c3#)) OR
 					(reg_q1443 AND symb_decoder(16#4d#)) OR
 					(reg_q1443 AND symb_decoder(16#f7#)) OR
 					(reg_q1443 AND symb_decoder(16#3f#)) OR
 					(reg_q1443 AND symb_decoder(16#79#)) OR
 					(reg_q1443 AND symb_decoder(16#fe#)) OR
 					(reg_q1443 AND symb_decoder(16#27#)) OR
 					(reg_q1443 AND symb_decoder(16#aa#)) OR
 					(reg_q1443 AND symb_decoder(16#6b#)) OR
 					(reg_q1443 AND symb_decoder(16#61#)) OR
 					(reg_q1443 AND symb_decoder(16#3c#)) OR
 					(reg_q1443 AND symb_decoder(16#a8#)) OR
 					(reg_q1443 AND symb_decoder(16#15#)) OR
 					(reg_q1443 AND symb_decoder(16#ef#)) OR
 					(reg_q1443 AND symb_decoder(16#59#)) OR
 					(reg_q1443 AND symb_decoder(16#42#)) OR
 					(reg_q1443 AND symb_decoder(16#1e#)) OR
 					(reg_q1443 AND symb_decoder(16#08#)) OR
 					(reg_q1443 AND symb_decoder(16#92#)) OR
 					(reg_q1443 AND symb_decoder(16#06#)) OR
 					(reg_q1443 AND symb_decoder(16#64#)) OR
 					(reg_q1443 AND symb_decoder(16#de#)) OR
 					(reg_q1443 AND symb_decoder(16#16#)) OR
 					(reg_q1443 AND symb_decoder(16#b2#)) OR
 					(reg_q1443 AND symb_decoder(16#0f#)) OR
 					(reg_q1443 AND symb_decoder(16#c0#)) OR
 					(reg_q1443 AND symb_decoder(16#49#)) OR
 					(reg_q1443 AND symb_decoder(16#2f#)) OR
 					(reg_q1443 AND symb_decoder(16#bf#)) OR
 					(reg_q1443 AND symb_decoder(16#91#)) OR
 					(reg_q1443 AND symb_decoder(16#26#)) OR
 					(reg_q1443 AND symb_decoder(16#12#)) OR
 					(reg_q1443 AND symb_decoder(16#7d#)) OR
 					(reg_q1443 AND symb_decoder(16#a4#)) OR
 					(reg_q1443 AND symb_decoder(16#c4#)) OR
 					(reg_q1443 AND symb_decoder(16#67#)) OR
 					(reg_q1443 AND symb_decoder(16#f2#)) OR
 					(reg_q1443 AND symb_decoder(16#6f#)) OR
 					(reg_q1443 AND symb_decoder(16#28#)) OR
 					(reg_q1443 AND symb_decoder(16#23#)) OR
 					(reg_q1443 AND symb_decoder(16#45#)) OR
 					(reg_q1443 AND symb_decoder(16#b0#)) OR
 					(reg_q1443 AND symb_decoder(16#9d#)) OR
 					(reg_q1443 AND symb_decoder(16#58#)) OR
 					(reg_q1443 AND symb_decoder(16#c8#)) OR
 					(reg_q1443 AND symb_decoder(16#7f#)) OR
 					(reg_q1443 AND symb_decoder(16#2d#)) OR
 					(reg_q1443 AND symb_decoder(16#56#)) OR
 					(reg_q1443 AND symb_decoder(16#1f#)) OR
 					(reg_q1443 AND symb_decoder(16#f4#)) OR
 					(reg_q1443 AND symb_decoder(16#c9#)) OR
 					(reg_q1443 AND symb_decoder(16#c7#)) OR
 					(reg_q1443 AND symb_decoder(16#0d#)) OR
 					(reg_q1443 AND symb_decoder(16#36#)) OR
 					(reg_q1443 AND symb_decoder(16#48#)) OR
 					(reg_q1443 AND symb_decoder(16#bc#)) OR
 					(reg_q1443 AND symb_decoder(16#4c#)) OR
 					(reg_q1443 AND symb_decoder(16#72#)) OR
 					(reg_q1443 AND symb_decoder(16#fc#)) OR
 					(reg_q1443 AND symb_decoder(16#1b#)) OR
 					(reg_q1443 AND symb_decoder(16#a1#)) OR
 					(reg_q1443 AND symb_decoder(16#ff#)) OR
 					(reg_q1443 AND symb_decoder(16#ae#)) OR
 					(reg_q1443 AND symb_decoder(16#0b#)) OR
 					(reg_q1443 AND symb_decoder(16#c5#)) OR
 					(reg_q1443 AND symb_decoder(16#a0#)) OR
 					(reg_q1443 AND symb_decoder(16#0c#)) OR
 					(reg_q1443 AND symb_decoder(16#84#)) OR
 					(reg_q1443 AND symb_decoder(16#cf#)) OR
 					(reg_q1443 AND symb_decoder(16#05#)) OR
 					(reg_q1443 AND symb_decoder(16#14#)) OR
 					(reg_q1443 AND symb_decoder(16#98#)) OR
 					(reg_q1443 AND symb_decoder(16#1c#)) OR
 					(reg_q1443 AND symb_decoder(16#e3#)) OR
 					(reg_q1443 AND symb_decoder(16#b6#)) OR
 					(reg_q1443 AND symb_decoder(16#ba#)) OR
 					(reg_q1443 AND symb_decoder(16#f9#));
reg_q1479_init <= '0' ;
	p_reg_q1479: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1479 <= reg_q1479_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1479 <= reg_q1479_init;
        else
          reg_q1479 <= reg_q1479_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2583_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q2583 AND symb_decoder(16#9c#)) OR
 					(reg_q2583 AND symb_decoder(16#2c#)) OR
 					(reg_q2583 AND symb_decoder(16#90#)) OR
 					(reg_q2583 AND symb_decoder(16#2a#)) OR
 					(reg_q2583 AND symb_decoder(16#54#)) OR
 					(reg_q2583 AND symb_decoder(16#2b#)) OR
 					(reg_q2583 AND symb_decoder(16#0b#)) OR
 					(reg_q2583 AND symb_decoder(16#75#)) OR
 					(reg_q2583 AND symb_decoder(16#dd#)) OR
 					(reg_q2583 AND symb_decoder(16#23#)) OR
 					(reg_q2583 AND symb_decoder(16#05#)) OR
 					(reg_q2583 AND symb_decoder(16#11#)) OR
 					(reg_q2583 AND symb_decoder(16#69#)) OR
 					(reg_q2583 AND symb_decoder(16#70#)) OR
 					(reg_q2583 AND symb_decoder(16#96#)) OR
 					(reg_q2583 AND symb_decoder(16#44#)) OR
 					(reg_q2583 AND symb_decoder(16#47#)) OR
 					(reg_q2583 AND symb_decoder(16#a1#)) OR
 					(reg_q2583 AND symb_decoder(16#e9#)) OR
 					(reg_q2583 AND symb_decoder(16#62#)) OR
 					(reg_q2583 AND symb_decoder(16#d8#)) OR
 					(reg_q2583 AND symb_decoder(16#bb#)) OR
 					(reg_q2583 AND symb_decoder(16#87#)) OR
 					(reg_q2583 AND symb_decoder(16#24#)) OR
 					(reg_q2583 AND symb_decoder(16#ab#)) OR
 					(reg_q2583 AND symb_decoder(16#9b#)) OR
 					(reg_q2583 AND symb_decoder(16#fb#)) OR
 					(reg_q2583 AND symb_decoder(16#83#)) OR
 					(reg_q2583 AND symb_decoder(16#ce#)) OR
 					(reg_q2583 AND symb_decoder(16#99#)) OR
 					(reg_q2583 AND symb_decoder(16#6f#)) OR
 					(reg_q2583 AND symb_decoder(16#91#)) OR
 					(reg_q2583 AND symb_decoder(16#98#)) OR
 					(reg_q2583 AND symb_decoder(16#19#)) OR
 					(reg_q2583 AND symb_decoder(16#16#)) OR
 					(reg_q2583 AND symb_decoder(16#73#)) OR
 					(reg_q2583 AND symb_decoder(16#6e#)) OR
 					(reg_q2583 AND symb_decoder(16#da#)) OR
 					(reg_q2583 AND symb_decoder(16#7f#)) OR
 					(reg_q2583 AND symb_decoder(16#bd#)) OR
 					(reg_q2583 AND symb_decoder(16#b9#)) OR
 					(reg_q2583 AND symb_decoder(16#88#)) OR
 					(reg_q2583 AND symb_decoder(16#93#)) OR
 					(reg_q2583 AND symb_decoder(16#36#)) OR
 					(reg_q2583 AND symb_decoder(16#08#)) OR
 					(reg_q2583 AND symb_decoder(16#2e#)) OR
 					(reg_q2583 AND symb_decoder(16#ed#)) OR
 					(reg_q2583 AND symb_decoder(16#32#)) OR
 					(reg_q2583 AND symb_decoder(16#17#)) OR
 					(reg_q2583 AND symb_decoder(16#49#)) OR
 					(reg_q2583 AND symb_decoder(16#1f#)) OR
 					(reg_q2583 AND symb_decoder(16#f9#)) OR
 					(reg_q2583 AND symb_decoder(16#1e#)) OR
 					(reg_q2583 AND symb_decoder(16#74#)) OR
 					(reg_q2583 AND symb_decoder(16#31#)) OR
 					(reg_q2583 AND symb_decoder(16#cd#)) OR
 					(reg_q2583 AND symb_decoder(16#aa#)) OR
 					(reg_q2583 AND symb_decoder(16#fc#)) OR
 					(reg_q2583 AND symb_decoder(16#56#)) OR
 					(reg_q2583 AND symb_decoder(16#58#)) OR
 					(reg_q2583 AND symb_decoder(16#a9#)) OR
 					(reg_q2583 AND symb_decoder(16#3c#)) OR
 					(reg_q2583 AND symb_decoder(16#42#)) OR
 					(reg_q2583 AND symb_decoder(16#d7#)) OR
 					(reg_q2583 AND symb_decoder(16#46#)) OR
 					(reg_q2583 AND symb_decoder(16#97#)) OR
 					(reg_q2583 AND symb_decoder(16#5e#)) OR
 					(reg_q2583 AND symb_decoder(16#b7#)) OR
 					(reg_q2583 AND symb_decoder(16#d4#)) OR
 					(reg_q2583 AND symb_decoder(16#ff#)) OR
 					(reg_q2583 AND symb_decoder(16#db#)) OR
 					(reg_q2583 AND symb_decoder(16#c2#)) OR
 					(reg_q2583 AND symb_decoder(16#79#)) OR
 					(reg_q2583 AND symb_decoder(16#f7#)) OR
 					(reg_q2583 AND symb_decoder(16#f8#)) OR
 					(reg_q2583 AND symb_decoder(16#78#)) OR
 					(reg_q2583 AND symb_decoder(16#d0#)) OR
 					(reg_q2583 AND symb_decoder(16#82#)) OR
 					(reg_q2583 AND symb_decoder(16#50#)) OR
 					(reg_q2583 AND symb_decoder(16#43#)) OR
 					(reg_q2583 AND symb_decoder(16#12#)) OR
 					(reg_q2583 AND symb_decoder(16#5b#)) OR
 					(reg_q2583 AND symb_decoder(16#b1#)) OR
 					(reg_q2583 AND symb_decoder(16#4e#)) OR
 					(reg_q2583 AND symb_decoder(16#40#)) OR
 					(reg_q2583 AND symb_decoder(16#de#)) OR
 					(reg_q2583 AND symb_decoder(16#37#)) OR
 					(reg_q2583 AND symb_decoder(16#4f#)) OR
 					(reg_q2583 AND symb_decoder(16#af#)) OR
 					(reg_q2583 AND symb_decoder(16#38#)) OR
 					(reg_q2583 AND symb_decoder(16#c4#)) OR
 					(reg_q2583 AND symb_decoder(16#59#)) OR
 					(reg_q2583 AND symb_decoder(16#57#)) OR
 					(reg_q2583 AND symb_decoder(16#ac#)) OR
 					(reg_q2583 AND symb_decoder(16#25#)) OR
 					(reg_q2583 AND symb_decoder(16#ef#)) OR
 					(reg_q2583 AND symb_decoder(16#60#)) OR
 					(reg_q2583 AND symb_decoder(16#45#)) OR
 					(reg_q2583 AND symb_decoder(16#fd#)) OR
 					(reg_q2583 AND symb_decoder(16#b0#)) OR
 					(reg_q2583 AND symb_decoder(16#48#)) OR
 					(reg_q2583 AND symb_decoder(16#03#)) OR
 					(reg_q2583 AND symb_decoder(16#04#)) OR
 					(reg_q2583 AND symb_decoder(16#be#)) OR
 					(reg_q2583 AND symb_decoder(16#7d#)) OR
 					(reg_q2583 AND symb_decoder(16#f3#)) OR
 					(reg_q2583 AND symb_decoder(16#3a#)) OR
 					(reg_q2583 AND symb_decoder(16#c5#)) OR
 					(reg_q2583 AND symb_decoder(16#e2#)) OR
 					(reg_q2583 AND symb_decoder(16#c7#)) OR
 					(reg_q2583 AND symb_decoder(16#15#)) OR
 					(reg_q2583 AND symb_decoder(16#c9#)) OR
 					(reg_q2583 AND symb_decoder(16#f1#)) OR
 					(reg_q2583 AND symb_decoder(16#6d#)) OR
 					(reg_q2583 AND symb_decoder(16#e6#)) OR
 					(reg_q2583 AND symb_decoder(16#06#)) OR
 					(reg_q2583 AND symb_decoder(16#10#)) OR
 					(reg_q2583 AND symb_decoder(16#7e#)) OR
 					(reg_q2583 AND symb_decoder(16#30#)) OR
 					(reg_q2583 AND symb_decoder(16#e8#)) OR
 					(reg_q2583 AND symb_decoder(16#fa#)) OR
 					(reg_q2583 AND symb_decoder(16#1a#)) OR
 					(reg_q2583 AND symb_decoder(16#21#)) OR
 					(reg_q2583 AND symb_decoder(16#4c#)) OR
 					(reg_q2583 AND symb_decoder(16#4a#)) OR
 					(reg_q2583 AND symb_decoder(16#8a#)) OR
 					(reg_q2583 AND symb_decoder(16#72#)) OR
 					(reg_q2583 AND symb_decoder(16#9a#)) OR
 					(reg_q2583 AND symb_decoder(16#77#)) OR
 					(reg_q2583 AND symb_decoder(16#d5#)) OR
 					(reg_q2583 AND symb_decoder(16#00#)) OR
 					(reg_q2583 AND symb_decoder(16#cb#)) OR
 					(reg_q2583 AND symb_decoder(16#64#)) OR
 					(reg_q2583 AND symb_decoder(16#ba#)) OR
 					(reg_q2583 AND symb_decoder(16#ea#)) OR
 					(reg_q2583 AND symb_decoder(16#b8#)) OR
 					(reg_q2583 AND symb_decoder(16#e0#)) OR
 					(reg_q2583 AND symb_decoder(16#9d#)) OR
 					(reg_q2583 AND symb_decoder(16#b4#)) OR
 					(reg_q2583 AND symb_decoder(16#14#)) OR
 					(reg_q2583 AND symb_decoder(16#fe#)) OR
 					(reg_q2583 AND symb_decoder(16#28#)) OR
 					(reg_q2583 AND symb_decoder(16#07#)) OR
 					(reg_q2583 AND symb_decoder(16#02#)) OR
 					(reg_q2583 AND symb_decoder(16#29#)) OR
 					(reg_q2583 AND symb_decoder(16#13#)) OR
 					(reg_q2583 AND symb_decoder(16#8f#)) OR
 					(reg_q2583 AND symb_decoder(16#d6#)) OR
 					(reg_q2583 AND symb_decoder(16#dc#)) OR
 					(reg_q2583 AND symb_decoder(16#c0#)) OR
 					(reg_q2583 AND symb_decoder(16#61#)) OR
 					(reg_q2583 AND symb_decoder(16#f6#)) OR
 					(reg_q2583 AND symb_decoder(16#01#)) OR
 					(reg_q2583 AND symb_decoder(16#c8#)) OR
 					(reg_q2583 AND symb_decoder(16#6c#)) OR
 					(reg_q2583 AND symb_decoder(16#55#)) OR
 					(reg_q2583 AND symb_decoder(16#b6#)) OR
 					(reg_q2583 AND symb_decoder(16#63#)) OR
 					(reg_q2583 AND symb_decoder(16#a7#)) OR
 					(reg_q2583 AND symb_decoder(16#22#)) OR
 					(reg_q2583 AND symb_decoder(16#d3#)) OR
 					(reg_q2583 AND symb_decoder(16#71#)) OR
 					(reg_q2583 AND symb_decoder(16#65#)) OR
 					(reg_q2583 AND symb_decoder(16#a8#)) OR
 					(reg_q2583 AND symb_decoder(16#20#)) OR
 					(reg_q2583 AND symb_decoder(16#c1#)) OR
 					(reg_q2583 AND symb_decoder(16#e5#)) OR
 					(reg_q2583 AND symb_decoder(16#b3#)) OR
 					(reg_q2583 AND symb_decoder(16#33#)) OR
 					(reg_q2583 AND symb_decoder(16#35#)) OR
 					(reg_q2583 AND symb_decoder(16#6b#)) OR
 					(reg_q2583 AND symb_decoder(16#80#)) OR
 					(reg_q2583 AND symb_decoder(16#f5#)) OR
 					(reg_q2583 AND symb_decoder(16#3d#)) OR
 					(reg_q2583 AND symb_decoder(16#2f#)) OR
 					(reg_q2583 AND symb_decoder(16#bf#)) OR
 					(reg_q2583 AND symb_decoder(16#e4#)) OR
 					(reg_q2583 AND symb_decoder(16#ee#)) OR
 					(reg_q2583 AND symb_decoder(16#0a#)) OR
 					(reg_q2583 AND symb_decoder(16#d1#)) OR
 					(reg_q2583 AND symb_decoder(16#1c#)) OR
 					(reg_q2583 AND symb_decoder(16#1d#)) OR
 					(reg_q2583 AND symb_decoder(16#89#)) OR
 					(reg_q2583 AND symb_decoder(16#8d#)) OR
 					(reg_q2583 AND symb_decoder(16#41#)) OR
 					(reg_q2583 AND symb_decoder(16#bc#)) OR
 					(reg_q2583 AND symb_decoder(16#e3#)) OR
 					(reg_q2583 AND symb_decoder(16#3b#)) OR
 					(reg_q2583 AND symb_decoder(16#85#)) OR
 					(reg_q2583 AND symb_decoder(16#d9#)) OR
 					(reg_q2583 AND symb_decoder(16#66#)) OR
 					(reg_q2583 AND symb_decoder(16#76#)) OR
 					(reg_q2583 AND symb_decoder(16#a3#)) OR
 					(reg_q2583 AND symb_decoder(16#5d#)) OR
 					(reg_q2583 AND symb_decoder(16#18#)) OR
 					(reg_q2583 AND symb_decoder(16#ec#)) OR
 					(reg_q2583 AND symb_decoder(16#5a#)) OR
 					(reg_q2583 AND symb_decoder(16#d2#)) OR
 					(reg_q2583 AND symb_decoder(16#5f#)) OR
 					(reg_q2583 AND symb_decoder(16#8b#)) OR
 					(reg_q2583 AND symb_decoder(16#51#)) OR
 					(reg_q2583 AND symb_decoder(16#81#)) OR
 					(reg_q2583 AND symb_decoder(16#09#)) OR
 					(reg_q2583 AND symb_decoder(16#ca#)) OR
 					(reg_q2583 AND symb_decoder(16#92#)) OR
 					(reg_q2583 AND symb_decoder(16#9f#)) OR
 					(reg_q2583 AND symb_decoder(16#2d#)) OR
 					(reg_q2583 AND symb_decoder(16#53#)) OR
 					(reg_q2583 AND symb_decoder(16#ad#)) OR
 					(reg_q2583 AND symb_decoder(16#cc#)) OR
 					(reg_q2583 AND symb_decoder(16#ae#)) OR
 					(reg_q2583 AND symb_decoder(16#3f#)) OR
 					(reg_q2583 AND symb_decoder(16#5c#)) OR
 					(reg_q2583 AND symb_decoder(16#f2#)) OR
 					(reg_q2583 AND symb_decoder(16#67#)) OR
 					(reg_q2583 AND symb_decoder(16#0e#)) OR
 					(reg_q2583 AND symb_decoder(16#34#)) OR
 					(reg_q2583 AND symb_decoder(16#4b#)) OR
 					(reg_q2583 AND symb_decoder(16#cf#)) OR
 					(reg_q2583 AND symb_decoder(16#26#)) OR
 					(reg_q2583 AND symb_decoder(16#1b#)) OR
 					(reg_q2583 AND symb_decoder(16#e1#)) OR
 					(reg_q2583 AND symb_decoder(16#f0#)) OR
 					(reg_q2583 AND symb_decoder(16#8c#)) OR
 					(reg_q2583 AND symb_decoder(16#4d#)) OR
 					(reg_q2583 AND symb_decoder(16#86#)) OR
 					(reg_q2583 AND symb_decoder(16#a6#)) OR
 					(reg_q2583 AND symb_decoder(16#0d#)) OR
 					(reg_q2583 AND symb_decoder(16#9e#)) OR
 					(reg_q2583 AND symb_decoder(16#3e#)) OR
 					(reg_q2583 AND symb_decoder(16#b2#)) OR
 					(reg_q2583 AND symb_decoder(16#52#)) OR
 					(reg_q2583 AND symb_decoder(16#c3#)) OR
 					(reg_q2583 AND symb_decoder(16#e7#)) OR
 					(reg_q2583 AND symb_decoder(16#7c#)) OR
 					(reg_q2583 AND symb_decoder(16#8e#)) OR
 					(reg_q2583 AND symb_decoder(16#27#)) OR
 					(reg_q2583 AND symb_decoder(16#f4#)) OR
 					(reg_q2583 AND symb_decoder(16#39#)) OR
 					(reg_q2583 AND symb_decoder(16#84#)) OR
 					(reg_q2583 AND symb_decoder(16#7a#)) OR
 					(reg_q2583 AND symb_decoder(16#eb#)) OR
 					(reg_q2583 AND symb_decoder(16#6a#)) OR
 					(reg_q2583 AND symb_decoder(16#95#)) OR
 					(reg_q2583 AND symb_decoder(16#68#)) OR
 					(reg_q2583 AND symb_decoder(16#df#)) OR
 					(reg_q2583 AND symb_decoder(16#a0#)) OR
 					(reg_q2583 AND symb_decoder(16#a2#)) OR
 					(reg_q2583 AND symb_decoder(16#94#)) OR
 					(reg_q2583 AND symb_decoder(16#0c#)) OR
 					(reg_q2583 AND symb_decoder(16#b5#)) OR
 					(reg_q2583 AND symb_decoder(16#0f#)) OR
 					(reg_q2583 AND symb_decoder(16#a4#)) OR
 					(reg_q2583 AND symb_decoder(16#a5#)) OR
 					(reg_q2583 AND symb_decoder(16#c6#)) OR
 					(reg_q2583 AND symb_decoder(16#7b#));
reg_q2583_init <= '0' ;
	p_reg_q2583: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2583 <= reg_q2583_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2583 <= reg_q2583_init;
        else
          reg_q2583 <= reg_q2583_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph20

reg_q393_in <= (reg_q377 AND symb_decoder(16#29#)) OR
 					(reg_q377 AND symb_decoder(16#05#)) OR
 					(reg_q377 AND symb_decoder(16#6e#)) OR
 					(reg_q377 AND symb_decoder(16#d3#)) OR
 					(reg_q377 AND symb_decoder(16#dd#)) OR
 					(reg_q377 AND symb_decoder(16#14#)) OR
 					(reg_q377 AND symb_decoder(16#f0#)) OR
 					(reg_q377 AND symb_decoder(16#ea#)) OR
 					(reg_q377 AND symb_decoder(16#83#)) OR
 					(reg_q377 AND symb_decoder(16#52#)) OR
 					(reg_q377 AND symb_decoder(16#7f#)) OR
 					(reg_q377 AND symb_decoder(16#a5#)) OR
 					(reg_q377 AND symb_decoder(16#df#)) OR
 					(reg_q377 AND symb_decoder(16#8d#)) OR
 					(reg_q377 AND symb_decoder(16#d5#)) OR
 					(reg_q377 AND symb_decoder(16#e1#)) OR
 					(reg_q377 AND symb_decoder(16#e3#)) OR
 					(reg_q377 AND symb_decoder(16#02#)) OR
 					(reg_q377 AND symb_decoder(16#64#)) OR
 					(reg_q377 AND symb_decoder(16#bd#)) OR
 					(reg_q377 AND symb_decoder(16#d9#)) OR
 					(reg_q377 AND symb_decoder(16#ee#)) OR
 					(reg_q377 AND symb_decoder(16#b1#)) OR
 					(reg_q377 AND symb_decoder(16#a1#)) OR
 					(reg_q377 AND symb_decoder(16#6d#)) OR
 					(reg_q377 AND symb_decoder(16#32#)) OR
 					(reg_q377 AND symb_decoder(16#c1#)) OR
 					(reg_q377 AND symb_decoder(16#69#)) OR
 					(reg_q377 AND symb_decoder(16#f8#)) OR
 					(reg_q377 AND symb_decoder(16#c9#)) OR
 					(reg_q377 AND symb_decoder(16#2a#)) OR
 					(reg_q377 AND symb_decoder(16#30#)) OR
 					(reg_q377 AND symb_decoder(16#16#)) OR
 					(reg_q377 AND symb_decoder(16#36#)) OR
 					(reg_q377 AND symb_decoder(16#12#)) OR
 					(reg_q377 AND symb_decoder(16#bc#)) OR
 					(reg_q377 AND symb_decoder(16#4b#)) OR
 					(reg_q377 AND symb_decoder(16#1b#)) OR
 					(reg_q377 AND symb_decoder(16#43#)) OR
 					(reg_q377 AND symb_decoder(16#03#)) OR
 					(reg_q377 AND symb_decoder(16#cd#)) OR
 					(reg_q377 AND symb_decoder(16#ff#)) OR
 					(reg_q377 AND symb_decoder(16#d2#)) OR
 					(reg_q377 AND symb_decoder(16#8f#)) OR
 					(reg_q377 AND symb_decoder(16#68#)) OR
 					(reg_q377 AND symb_decoder(16#7c#)) OR
 					(reg_q377 AND symb_decoder(16#9c#)) OR
 					(reg_q377 AND symb_decoder(16#61#)) OR
 					(reg_q377 AND symb_decoder(16#31#)) OR
 					(reg_q377 AND symb_decoder(16#63#)) OR
 					(reg_q377 AND symb_decoder(16#37#)) OR
 					(reg_q377 AND symb_decoder(16#0e#)) OR
 					(reg_q377 AND symb_decoder(16#e7#)) OR
 					(reg_q377 AND symb_decoder(16#89#)) OR
 					(reg_q377 AND symb_decoder(16#f7#)) OR
 					(reg_q377 AND symb_decoder(16#d1#)) OR
 					(reg_q377 AND symb_decoder(16#35#)) OR
 					(reg_q377 AND symb_decoder(16#dc#)) OR
 					(reg_q377 AND symb_decoder(16#73#)) OR
 					(reg_q377 AND symb_decoder(16#c0#)) OR
 					(reg_q377 AND symb_decoder(16#8a#)) OR
 					(reg_q377 AND symb_decoder(16#d7#)) OR
 					(reg_q377 AND symb_decoder(16#f4#)) OR
 					(reg_q377 AND symb_decoder(16#3a#)) OR
 					(reg_q377 AND symb_decoder(16#0b#)) OR
 					(reg_q377 AND symb_decoder(16#42#)) OR
 					(reg_q377 AND symb_decoder(16#01#)) OR
 					(reg_q377 AND symb_decoder(16#ef#)) OR
 					(reg_q377 AND symb_decoder(16#b3#)) OR
 					(reg_q377 AND symb_decoder(16#25#)) OR
 					(reg_q377 AND symb_decoder(16#b2#)) OR
 					(reg_q377 AND symb_decoder(16#3c#)) OR
 					(reg_q377 AND symb_decoder(16#7a#)) OR
 					(reg_q377 AND symb_decoder(16#00#)) OR
 					(reg_q377 AND symb_decoder(16#93#)) OR
 					(reg_q377 AND symb_decoder(16#53#)) OR
 					(reg_q377 AND symb_decoder(16#98#)) OR
 					(reg_q377 AND symb_decoder(16#b4#)) OR
 					(reg_q377 AND symb_decoder(16#c5#)) OR
 					(reg_q377 AND symb_decoder(16#79#)) OR
 					(reg_q377 AND symb_decoder(16#4f#)) OR
 					(reg_q377 AND symb_decoder(16#74#)) OR
 					(reg_q377 AND symb_decoder(16#17#)) OR
 					(reg_q377 AND symb_decoder(16#d4#)) OR
 					(reg_q377 AND symb_decoder(16#4a#)) OR
 					(reg_q377 AND symb_decoder(16#4c#)) OR
 					(reg_q377 AND symb_decoder(16#ae#)) OR
 					(reg_q377 AND symb_decoder(16#d8#)) OR
 					(reg_q377 AND symb_decoder(16#7b#)) OR
 					(reg_q377 AND symb_decoder(16#07#)) OR
 					(reg_q377 AND symb_decoder(16#2c#)) OR
 					(reg_q377 AND symb_decoder(16#b5#)) OR
 					(reg_q377 AND symb_decoder(16#a8#)) OR
 					(reg_q377 AND symb_decoder(16#cf#)) OR
 					(reg_q377 AND symb_decoder(16#82#)) OR
 					(reg_q377 AND symb_decoder(16#d6#)) OR
 					(reg_q377 AND symb_decoder(16#80#)) OR
 					(reg_q377 AND symb_decoder(16#eb#)) OR
 					(reg_q377 AND symb_decoder(16#9a#)) OR
 					(reg_q377 AND symb_decoder(16#40#)) OR
 					(reg_q377 AND symb_decoder(16#95#)) OR
 					(reg_q377 AND symb_decoder(16#e9#)) OR
 					(reg_q377 AND symb_decoder(16#a3#)) OR
 					(reg_q377 AND symb_decoder(16#e4#)) OR
 					(reg_q377 AND symb_decoder(16#11#)) OR
 					(reg_q377 AND symb_decoder(16#2e#)) OR
 					(reg_q377 AND symb_decoder(16#fc#)) OR
 					(reg_q377 AND symb_decoder(16#0c#)) OR
 					(reg_q377 AND symb_decoder(16#27#)) OR
 					(reg_q377 AND symb_decoder(16#67#)) OR
 					(reg_q377 AND symb_decoder(16#7d#)) OR
 					(reg_q377 AND symb_decoder(16#6f#)) OR
 					(reg_q377 AND symb_decoder(16#1f#)) OR
 					(reg_q377 AND symb_decoder(16#8e#)) OR
 					(reg_q377 AND symb_decoder(16#f3#)) OR
 					(reg_q377 AND symb_decoder(16#db#)) OR
 					(reg_q377 AND symb_decoder(16#fa#)) OR
 					(reg_q377 AND symb_decoder(16#21#)) OR
 					(reg_q377 AND symb_decoder(16#48#)) OR
 					(reg_q377 AND symb_decoder(16#1c#)) OR
 					(reg_q377 AND symb_decoder(16#66#)) OR
 					(reg_q377 AND symb_decoder(16#b0#)) OR
 					(reg_q377 AND symb_decoder(16#75#)) OR
 					(reg_q377 AND symb_decoder(16#23#)) OR
 					(reg_q377 AND symb_decoder(16#be#)) OR
 					(reg_q377 AND symb_decoder(16#81#)) OR
 					(reg_q377 AND symb_decoder(16#94#)) OR
 					(reg_q377 AND symb_decoder(16#13#)) OR
 					(reg_q377 AND symb_decoder(16#e2#)) OR
 					(reg_q377 AND symb_decoder(16#1a#)) OR
 					(reg_q377 AND symb_decoder(16#8c#)) OR
 					(reg_q377 AND symb_decoder(16#0f#)) OR
 					(reg_q377 AND symb_decoder(16#78#)) OR
 					(reg_q377 AND symb_decoder(16#4e#)) OR
 					(reg_q377 AND symb_decoder(16#88#)) OR
 					(reg_q377 AND symb_decoder(16#6b#)) OR
 					(reg_q377 AND symb_decoder(16#2f#)) OR
 					(reg_q377 AND symb_decoder(16#e0#)) OR
 					(reg_q377 AND symb_decoder(16#f5#)) OR
 					(reg_q377 AND symb_decoder(16#d0#)) OR
 					(reg_q377 AND symb_decoder(16#24#)) OR
 					(reg_q377 AND symb_decoder(16#09#)) OR
 					(reg_q377 AND symb_decoder(16#bb#)) OR
 					(reg_q377 AND symb_decoder(16#59#)) OR
 					(reg_q377 AND symb_decoder(16#c3#)) OR
 					(reg_q377 AND symb_decoder(16#e5#)) OR
 					(reg_q377 AND symb_decoder(16#de#)) OR
 					(reg_q377 AND symb_decoder(16#19#)) OR
 					(reg_q377 AND symb_decoder(16#fd#)) OR
 					(reg_q377 AND symb_decoder(16#47#)) OR
 					(reg_q377 AND symb_decoder(16#b6#)) OR
 					(reg_q377 AND symb_decoder(16#e6#)) OR
 					(reg_q377 AND symb_decoder(16#65#)) OR
 					(reg_q377 AND symb_decoder(16#ba#)) OR
 					(reg_q377 AND symb_decoder(16#38#)) OR
 					(reg_q377 AND symb_decoder(16#84#)) OR
 					(reg_q377 AND symb_decoder(16#96#)) OR
 					(reg_q377 AND symb_decoder(16#c4#)) OR
 					(reg_q377 AND symb_decoder(16#26#)) OR
 					(reg_q377 AND symb_decoder(16#b9#)) OR
 					(reg_q377 AND symb_decoder(16#a7#)) OR
 					(reg_q377 AND symb_decoder(16#3f#)) OR
 					(reg_q377 AND symb_decoder(16#55#)) OR
 					(reg_q377 AND symb_decoder(16#f6#)) OR
 					(reg_q377 AND symb_decoder(16#6c#)) OR
 					(reg_q377 AND symb_decoder(16#57#)) OR
 					(reg_q377 AND symb_decoder(16#22#)) OR
 					(reg_q377 AND symb_decoder(16#f1#)) OR
 					(reg_q377 AND symb_decoder(16#5e#)) OR
 					(reg_q377 AND symb_decoder(16#da#)) OR
 					(reg_q377 AND symb_decoder(16#08#)) OR
 					(reg_q377 AND symb_decoder(16#a0#)) OR
 					(reg_q377 AND symb_decoder(16#90#)) OR
 					(reg_q377 AND symb_decoder(16#9f#)) OR
 					(reg_q377 AND symb_decoder(16#72#)) OR
 					(reg_q377 AND symb_decoder(16#77#)) OR
 					(reg_q377 AND symb_decoder(16#2d#)) OR
 					(reg_q377 AND symb_decoder(16#51#)) OR
 					(reg_q377 AND symb_decoder(16#34#)) OR
 					(reg_q377 AND symb_decoder(16#ed#)) OR
 					(reg_q377 AND symb_decoder(16#cb#)) OR
 					(reg_q377 AND symb_decoder(16#92#)) OR
 					(reg_q377 AND symb_decoder(16#33#)) OR
 					(reg_q377 AND symb_decoder(16#e8#)) OR
 					(reg_q377 AND symb_decoder(16#1d#)) OR
 					(reg_q377 AND symb_decoder(16#41#)) OR
 					(reg_q377 AND symb_decoder(16#5d#)) OR
 					(reg_q377 AND symb_decoder(16#6a#)) OR
 					(reg_q377 AND symb_decoder(16#91#)) OR
 					(reg_q377 AND symb_decoder(16#4d#)) OR
 					(reg_q377 AND symb_decoder(16#2b#)) OR
 					(reg_q377 AND symb_decoder(16#70#)) OR
 					(reg_q377 AND symb_decoder(16#5c#)) OR
 					(reg_q377 AND symb_decoder(16#ca#)) OR
 					(reg_q377 AND symb_decoder(16#04#)) OR
 					(reg_q377 AND symb_decoder(16#15#)) OR
 					(reg_q377 AND symb_decoder(16#cc#)) OR
 					(reg_q377 AND symb_decoder(16#97#)) OR
 					(reg_q377 AND symb_decoder(16#ac#)) OR
 					(reg_q377 AND symb_decoder(16#b8#)) OR
 					(reg_q377 AND symb_decoder(16#7e#)) OR
 					(reg_q377 AND symb_decoder(16#bf#)) OR
 					(reg_q377 AND symb_decoder(16#50#)) OR
 					(reg_q377 AND symb_decoder(16#45#)) OR
 					(reg_q377 AND symb_decoder(16#f2#)) OR
 					(reg_q377 AND symb_decoder(16#87#)) OR
 					(reg_q377 AND symb_decoder(16#60#)) OR
 					(reg_q377 AND symb_decoder(16#18#)) OR
 					(reg_q377 AND symb_decoder(16#a2#)) OR
 					(reg_q377 AND symb_decoder(16#54#)) OR
 					(reg_q377 AND symb_decoder(16#3b#)) OR
 					(reg_q377 AND symb_decoder(16#06#)) OR
 					(reg_q377 AND symb_decoder(16#5b#)) OR
 					(reg_q377 AND symb_decoder(16#20#)) OR
 					(reg_q377 AND symb_decoder(16#44#)) OR
 					(reg_q377 AND symb_decoder(16#99#)) OR
 					(reg_q377 AND symb_decoder(16#ab#)) OR
 					(reg_q377 AND symb_decoder(16#b7#)) OR
 					(reg_q377 AND symb_decoder(16#8b#)) OR
 					(reg_q377 AND symb_decoder(16#56#)) OR
 					(reg_q377 AND symb_decoder(16#5f#)) OR
 					(reg_q377 AND symb_decoder(16#39#)) OR
 					(reg_q377 AND symb_decoder(16#af#)) OR
 					(reg_q377 AND symb_decoder(16#1e#)) OR
 					(reg_q377 AND symb_decoder(16#c6#)) OR
 					(reg_q377 AND symb_decoder(16#3d#)) OR
 					(reg_q377 AND symb_decoder(16#a4#)) OR
 					(reg_q377 AND symb_decoder(16#10#)) OR
 					(reg_q377 AND symb_decoder(16#58#)) OR
 					(reg_q377 AND symb_decoder(16#c2#)) OR
 					(reg_q377 AND symb_decoder(16#46#)) OR
 					(reg_q377 AND symb_decoder(16#c7#)) OR
 					(reg_q377 AND symb_decoder(16#28#)) OR
 					(reg_q377 AND symb_decoder(16#a6#)) OR
 					(reg_q377 AND symb_decoder(16#76#)) OR
 					(reg_q377 AND symb_decoder(16#f9#)) OR
 					(reg_q377 AND symb_decoder(16#c8#)) OR
 					(reg_q377 AND symb_decoder(16#ad#)) OR
 					(reg_q377 AND symb_decoder(16#86#)) OR
 					(reg_q377 AND symb_decoder(16#49#)) OR
 					(reg_q377 AND symb_decoder(16#fe#)) OR
 					(reg_q377 AND symb_decoder(16#ce#)) OR
 					(reg_q377 AND symb_decoder(16#9e#)) OR
 					(reg_q377 AND symb_decoder(16#85#)) OR
 					(reg_q377 AND symb_decoder(16#9d#)) OR
 					(reg_q377 AND symb_decoder(16#9b#)) OR
 					(reg_q377 AND symb_decoder(16#a9#)) OR
 					(reg_q377 AND symb_decoder(16#3e#)) OR
 					(reg_q377 AND symb_decoder(16#62#)) OR
 					(reg_q377 AND symb_decoder(16#ec#)) OR
 					(reg_q377 AND symb_decoder(16#fb#)) OR
 					(reg_q377 AND symb_decoder(16#5a#)) OR
 					(reg_q377 AND symb_decoder(16#aa#)) OR
 					(reg_q377 AND symb_decoder(16#71#)) OR
 					(reg_q393 AND symb_decoder(16#e2#)) OR
 					(reg_q393 AND symb_decoder(16#ba#)) OR
 					(reg_q393 AND symb_decoder(16#c7#)) OR
 					(reg_q393 AND symb_decoder(16#8a#)) OR
 					(reg_q393 AND symb_decoder(16#e9#)) OR
 					(reg_q393 AND symb_decoder(16#a3#)) OR
 					(reg_q393 AND symb_decoder(16#9d#)) OR
 					(reg_q393 AND symb_decoder(16#38#)) OR
 					(reg_q393 AND symb_decoder(16#ff#)) OR
 					(reg_q393 AND symb_decoder(16#08#)) OR
 					(reg_q393 AND symb_decoder(16#cd#)) OR
 					(reg_q393 AND symb_decoder(16#36#)) OR
 					(reg_q393 AND symb_decoder(16#49#)) OR
 					(reg_q393 AND symb_decoder(16#14#)) OR
 					(reg_q393 AND symb_decoder(16#d1#)) OR
 					(reg_q393 AND symb_decoder(16#77#)) OR
 					(reg_q393 AND symb_decoder(16#b4#)) OR
 					(reg_q393 AND symb_decoder(16#70#)) OR
 					(reg_q393 AND symb_decoder(16#8b#)) OR
 					(reg_q393 AND symb_decoder(16#c9#)) OR
 					(reg_q393 AND symb_decoder(16#97#)) OR
 					(reg_q393 AND symb_decoder(16#8c#)) OR
 					(reg_q393 AND symb_decoder(16#a9#)) OR
 					(reg_q393 AND symb_decoder(16#75#)) OR
 					(reg_q393 AND symb_decoder(16#eb#)) OR
 					(reg_q393 AND symb_decoder(16#1f#)) OR
 					(reg_q393 AND symb_decoder(16#e6#)) OR
 					(reg_q393 AND symb_decoder(16#23#)) OR
 					(reg_q393 AND symb_decoder(16#47#)) OR
 					(reg_q393 AND symb_decoder(16#74#)) OR
 					(reg_q393 AND symb_decoder(16#6a#)) OR
 					(reg_q393 AND symb_decoder(16#a4#)) OR
 					(reg_q393 AND symb_decoder(16#12#)) OR
 					(reg_q393 AND symb_decoder(16#e3#)) OR
 					(reg_q393 AND symb_decoder(16#13#)) OR
 					(reg_q393 AND symb_decoder(16#42#)) OR
 					(reg_q393 AND symb_decoder(16#55#)) OR
 					(reg_q393 AND symb_decoder(16#c6#)) OR
 					(reg_q393 AND symb_decoder(16#9e#)) OR
 					(reg_q393 AND symb_decoder(16#96#)) OR
 					(reg_q393 AND symb_decoder(16#39#)) OR
 					(reg_q393 AND symb_decoder(16#7e#)) OR
 					(reg_q393 AND symb_decoder(16#22#)) OR
 					(reg_q393 AND symb_decoder(16#fb#)) OR
 					(reg_q393 AND symb_decoder(16#09#)) OR
 					(reg_q393 AND symb_decoder(16#5a#)) OR
 					(reg_q393 AND symb_decoder(16#82#)) OR
 					(reg_q393 AND symb_decoder(16#3a#)) OR
 					(reg_q393 AND symb_decoder(16#cf#)) OR
 					(reg_q393 AND symb_decoder(16#c5#)) OR
 					(reg_q393 AND symb_decoder(16#26#)) OR
 					(reg_q393 AND symb_decoder(16#24#)) OR
 					(reg_q393 AND symb_decoder(16#17#)) OR
 					(reg_q393 AND symb_decoder(16#34#)) OR
 					(reg_q393 AND symb_decoder(16#48#)) OR
 					(reg_q393 AND symb_decoder(16#ec#)) OR
 					(reg_q393 AND symb_decoder(16#02#)) OR
 					(reg_q393 AND symb_decoder(16#8e#)) OR
 					(reg_q393 AND symb_decoder(16#be#)) OR
 					(reg_q393 AND symb_decoder(16#7c#)) OR
 					(reg_q393 AND symb_decoder(16#6b#)) OR
 					(reg_q393 AND symb_decoder(16#f8#)) OR
 					(reg_q393 AND symb_decoder(16#19#)) OR
 					(reg_q393 AND symb_decoder(16#fd#)) OR
 					(reg_q393 AND symb_decoder(16#4a#)) OR
 					(reg_q393 AND symb_decoder(16#da#)) OR
 					(reg_q393 AND symb_decoder(16#f0#)) OR
 					(reg_q393 AND symb_decoder(16#2d#)) OR
 					(reg_q393 AND symb_decoder(16#3b#)) OR
 					(reg_q393 AND symb_decoder(16#07#)) OR
 					(reg_q393 AND symb_decoder(16#41#)) OR
 					(reg_q393 AND symb_decoder(16#a2#)) OR
 					(reg_q393 AND symb_decoder(16#16#)) OR
 					(reg_q393 AND symb_decoder(16#35#)) OR
 					(reg_q393 AND symb_decoder(16#e4#)) OR
 					(reg_q393 AND symb_decoder(16#69#)) OR
 					(reg_q393 AND symb_decoder(16#37#)) OR
 					(reg_q393 AND symb_decoder(16#29#)) OR
 					(reg_q393 AND symb_decoder(16#01#)) OR
 					(reg_q393 AND symb_decoder(16#7b#)) OR
 					(reg_q393 AND symb_decoder(16#db#)) OR
 					(reg_q393 AND symb_decoder(16#f7#)) OR
 					(reg_q393 AND symb_decoder(16#df#)) OR
 					(reg_q393 AND symb_decoder(16#dd#)) OR
 					(reg_q393 AND symb_decoder(16#53#)) OR
 					(reg_q393 AND symb_decoder(16#f2#)) OR
 					(reg_q393 AND symb_decoder(16#d6#)) OR
 					(reg_q393 AND symb_decoder(16#89#)) OR
 					(reg_q393 AND symb_decoder(16#f4#)) OR
 					(reg_q393 AND symb_decoder(16#63#)) OR
 					(reg_q393 AND symb_decoder(16#bf#)) OR
 					(reg_q393 AND symb_decoder(16#72#)) OR
 					(reg_q393 AND symb_decoder(16#06#)) OR
 					(reg_q393 AND symb_decoder(16#af#)) OR
 					(reg_q393 AND symb_decoder(16#a0#)) OR
 					(reg_q393 AND symb_decoder(16#84#)) OR
 					(reg_q393 AND symb_decoder(16#76#)) OR
 					(reg_q393 AND symb_decoder(16#d2#)) OR
 					(reg_q393 AND symb_decoder(16#d3#)) OR
 					(reg_q393 AND symb_decoder(16#4e#)) OR
 					(reg_q393 AND symb_decoder(16#25#)) OR
 					(reg_q393 AND symb_decoder(16#30#)) OR
 					(reg_q393 AND symb_decoder(16#ef#)) OR
 					(reg_q393 AND symb_decoder(16#b7#)) OR
 					(reg_q393 AND symb_decoder(16#66#)) OR
 					(reg_q393 AND symb_decoder(16#5e#)) OR
 					(reg_q393 AND symb_decoder(16#e8#)) OR
 					(reg_q393 AND symb_decoder(16#78#)) OR
 					(reg_q393 AND symb_decoder(16#73#)) OR
 					(reg_q393 AND symb_decoder(16#e0#)) OR
 					(reg_q393 AND symb_decoder(16#94#)) OR
 					(reg_q393 AND symb_decoder(16#04#)) OR
 					(reg_q393 AND symb_decoder(16#d0#)) OR
 					(reg_q393 AND symb_decoder(16#1e#)) OR
 					(reg_q393 AND symb_decoder(16#68#)) OR
 					(reg_q393 AND symb_decoder(16#d7#)) OR
 					(reg_q393 AND symb_decoder(16#6d#)) OR
 					(reg_q393 AND symb_decoder(16#5c#)) OR
 					(reg_q393 AND symb_decoder(16#e7#)) OR
 					(reg_q393 AND symb_decoder(16#10#)) OR
 					(reg_q393 AND symb_decoder(16#a6#)) OR
 					(reg_q393 AND symb_decoder(16#9b#)) OR
 					(reg_q393 AND symb_decoder(16#9c#)) OR
 					(reg_q393 AND symb_decoder(16#54#)) OR
 					(reg_q393 AND symb_decoder(16#b2#)) OR
 					(reg_q393 AND symb_decoder(16#88#)) OR
 					(reg_q393 AND symb_decoder(16#21#)) OR
 					(reg_q393 AND symb_decoder(16#9a#)) OR
 					(reg_q393 AND symb_decoder(16#9f#)) OR
 					(reg_q393 AND symb_decoder(16#a7#)) OR
 					(reg_q393 AND symb_decoder(16#65#)) OR
 					(reg_q393 AND symb_decoder(16#1c#)) OR
 					(reg_q393 AND symb_decoder(16#4d#)) OR
 					(reg_q393 AND symb_decoder(16#b5#)) OR
 					(reg_q393 AND symb_decoder(16#7f#)) OR
 					(reg_q393 AND symb_decoder(16#b9#)) OR
 					(reg_q393 AND symb_decoder(16#85#)) OR
 					(reg_q393 AND symb_decoder(16#90#)) OR
 					(reg_q393 AND symb_decoder(16#7a#)) OR
 					(reg_q393 AND symb_decoder(16#4c#)) OR
 					(reg_q393 AND symb_decoder(16#80#)) OR
 					(reg_q393 AND symb_decoder(16#79#)) OR
 					(reg_q393 AND symb_decoder(16#58#)) OR
 					(reg_q393 AND symb_decoder(16#1b#)) OR
 					(reg_q393 AND symb_decoder(16#64#)) OR
 					(reg_q393 AND symb_decoder(16#15#)) OR
 					(reg_q393 AND symb_decoder(16#32#)) OR
 					(reg_q393 AND symb_decoder(16#ee#)) OR
 					(reg_q393 AND symb_decoder(16#cb#)) OR
 					(reg_q393 AND symb_decoder(16#ac#)) OR
 					(reg_q393 AND symb_decoder(16#60#)) OR
 					(reg_q393 AND symb_decoder(16#2c#)) OR
 					(reg_q393 AND symb_decoder(16#a1#)) OR
 					(reg_q393 AND symb_decoder(16#d5#)) OR
 					(reg_q393 AND symb_decoder(16#27#)) OR
 					(reg_q393 AND symb_decoder(16#33#)) OR
 					(reg_q393 AND symb_decoder(16#c0#)) OR
 					(reg_q393 AND symb_decoder(16#c1#)) OR
 					(reg_q393 AND symb_decoder(16#6c#)) OR
 					(reg_q393 AND symb_decoder(16#95#)) OR
 					(reg_q393 AND symb_decoder(16#71#)) OR
 					(reg_q393 AND symb_decoder(16#56#)) OR
 					(reg_q393 AND symb_decoder(16#c2#)) OR
 					(reg_q393 AND symb_decoder(16#a5#)) OR
 					(reg_q393 AND symb_decoder(16#98#)) OR
 					(reg_q393 AND symb_decoder(16#31#)) OR
 					(reg_q393 AND symb_decoder(16#ab#)) OR
 					(reg_q393 AND symb_decoder(16#b0#)) OR
 					(reg_q393 AND symb_decoder(16#bb#)) OR
 					(reg_q393 AND symb_decoder(16#0e#)) OR
 					(reg_q393 AND symb_decoder(16#ed#)) OR
 					(reg_q393 AND symb_decoder(16#fc#)) OR
 					(reg_q393 AND symb_decoder(16#d8#)) OR
 					(reg_q393 AND symb_decoder(16#7d#)) OR
 					(reg_q393 AND symb_decoder(16#bc#)) OR
 					(reg_q393 AND symb_decoder(16#c3#)) OR
 					(reg_q393 AND symb_decoder(16#fe#)) OR
 					(reg_q393 AND symb_decoder(16#b8#)) OR
 					(reg_q393 AND symb_decoder(16#57#)) OR
 					(reg_q393 AND symb_decoder(16#03#)) OR
 					(reg_q393 AND symb_decoder(16#93#)) OR
 					(reg_q393 AND symb_decoder(16#fa#)) OR
 					(reg_q393 AND symb_decoder(16#c4#)) OR
 					(reg_q393 AND symb_decoder(16#44#)) OR
 					(reg_q393 AND symb_decoder(16#f3#)) OR
 					(reg_q393 AND symb_decoder(16#f9#)) OR
 					(reg_q393 AND symb_decoder(16#8f#)) OR
 					(reg_q393 AND symb_decoder(16#43#)) OR
 					(reg_q393 AND symb_decoder(16#45#)) OR
 					(reg_q393 AND symb_decoder(16#91#)) OR
 					(reg_q393 AND symb_decoder(16#5f#)) OR
 					(reg_q393 AND symb_decoder(16#20#)) OR
 					(reg_q393 AND symb_decoder(16#ad#)) OR
 					(reg_q393 AND symb_decoder(16#ae#)) OR
 					(reg_q393 AND symb_decoder(16#52#)) OR
 					(reg_q393 AND symb_decoder(16#59#)) OR
 					(reg_q393 AND symb_decoder(16#1d#)) OR
 					(reg_q393 AND symb_decoder(16#d9#)) OR
 					(reg_q393 AND symb_decoder(16#1a#)) OR
 					(reg_q393 AND symb_decoder(16#b6#)) OR
 					(reg_q393 AND symb_decoder(16#40#)) OR
 					(reg_q393 AND symb_decoder(16#92#)) OR
 					(reg_q393 AND symb_decoder(16#87#)) OR
 					(reg_q393 AND symb_decoder(16#6f#)) OR
 					(reg_q393 AND symb_decoder(16#f6#)) OR
 					(reg_q393 AND symb_decoder(16#f5#)) OR
 					(reg_q393 AND symb_decoder(16#6e#)) OR
 					(reg_q393 AND symb_decoder(16#4f#)) OR
 					(reg_q393 AND symb_decoder(16#5d#)) OR
 					(reg_q393 AND symb_decoder(16#e5#)) OR
 					(reg_q393 AND symb_decoder(16#46#)) OR
 					(reg_q393 AND symb_decoder(16#e1#)) OR
 					(reg_q393 AND symb_decoder(16#d4#)) OR
 					(reg_q393 AND symb_decoder(16#50#)) OR
 					(reg_q393 AND symb_decoder(16#b3#)) OR
 					(reg_q393 AND symb_decoder(16#05#)) OR
 					(reg_q393 AND symb_decoder(16#3c#)) OR
 					(reg_q393 AND symb_decoder(16#cc#)) OR
 					(reg_q393 AND symb_decoder(16#2a#)) OR
 					(reg_q393 AND symb_decoder(16#2f#)) OR
 					(reg_q393 AND symb_decoder(16#de#)) OR
 					(reg_q393 AND symb_decoder(16#2b#)) OR
 					(reg_q393 AND symb_decoder(16#4b#)) OR
 					(reg_q393 AND symb_decoder(16#00#)) OR
 					(reg_q393 AND symb_decoder(16#51#)) OR
 					(reg_q393 AND symb_decoder(16#99#)) OR
 					(reg_q393 AND symb_decoder(16#0f#)) OR
 					(reg_q393 AND symb_decoder(16#3f#)) OR
 					(reg_q393 AND symb_decoder(16#28#)) OR
 					(reg_q393 AND symb_decoder(16#5b#)) OR
 					(reg_q393 AND symb_decoder(16#b1#)) OR
 					(reg_q393 AND symb_decoder(16#aa#)) OR
 					(reg_q393 AND symb_decoder(16#0c#)) OR
 					(reg_q393 AND symb_decoder(16#ea#)) OR
 					(reg_q393 AND symb_decoder(16#2e#)) OR
 					(reg_q393 AND symb_decoder(16#0b#)) OR
 					(reg_q393 AND symb_decoder(16#ca#)) OR
 					(reg_q393 AND symb_decoder(16#81#)) OR
 					(reg_q393 AND symb_decoder(16#18#)) OR
 					(reg_q393 AND symb_decoder(16#8d#)) OR
 					(reg_q393 AND symb_decoder(16#dc#)) OR
 					(reg_q393 AND symb_decoder(16#86#)) OR
 					(reg_q393 AND symb_decoder(16#67#)) OR
 					(reg_q393 AND symb_decoder(16#62#)) OR
 					(reg_q393 AND symb_decoder(16#c8#)) OR
 					(reg_q393 AND symb_decoder(16#a8#)) OR
 					(reg_q393 AND symb_decoder(16#f1#)) OR
 					(reg_q393 AND symb_decoder(16#61#)) OR
 					(reg_q393 AND symb_decoder(16#83#)) OR
 					(reg_q393 AND symb_decoder(16#bd#)) OR
 					(reg_q393 AND symb_decoder(16#ce#)) OR
 					(reg_q393 AND symb_decoder(16#3e#)) OR
 					(reg_q393 AND symb_decoder(16#11#)) OR
 					(reg_q393 AND symb_decoder(16#3d#));
reg_q542_in <= (reg_q522 AND symb_decoder(16#da#)) OR
 					(reg_q522 AND symb_decoder(16#5a#)) OR
 					(reg_q522 AND symb_decoder(16#60#)) OR
 					(reg_q522 AND symb_decoder(16#ab#)) OR
 					(reg_q522 AND symb_decoder(16#68#)) OR
 					(reg_q522 AND symb_decoder(16#52#)) OR
 					(reg_q522 AND symb_decoder(16#01#)) OR
 					(reg_q522 AND symb_decoder(16#e4#)) OR
 					(reg_q522 AND symb_decoder(16#ef#)) OR
 					(reg_q522 AND symb_decoder(16#ed#)) OR
 					(reg_q522 AND symb_decoder(16#3e#)) OR
 					(reg_q522 AND symb_decoder(16#34#)) OR
 					(reg_q522 AND symb_decoder(16#cc#)) OR
 					(reg_q522 AND symb_decoder(16#70#)) OR
 					(reg_q522 AND symb_decoder(16#79#)) OR
 					(reg_q522 AND symb_decoder(16#ff#)) OR
 					(reg_q522 AND symb_decoder(16#6f#)) OR
 					(reg_q522 AND symb_decoder(16#64#)) OR
 					(reg_q522 AND symb_decoder(16#8e#)) OR
 					(reg_q522 AND symb_decoder(16#e6#)) OR
 					(reg_q522 AND symb_decoder(16#47#)) OR
 					(reg_q522 AND symb_decoder(16#d0#)) OR
 					(reg_q522 AND symb_decoder(16#10#)) OR
 					(reg_q522 AND symb_decoder(16#bf#)) OR
 					(reg_q522 AND symb_decoder(16#22#)) OR
 					(reg_q522 AND symb_decoder(16#41#)) OR
 					(reg_q522 AND symb_decoder(16#2d#)) OR
 					(reg_q522 AND symb_decoder(16#11#)) OR
 					(reg_q522 AND symb_decoder(16#e7#)) OR
 					(reg_q522 AND symb_decoder(16#1e#)) OR
 					(reg_q522 AND symb_decoder(16#0e#)) OR
 					(reg_q522 AND symb_decoder(16#a5#)) OR
 					(reg_q522 AND symb_decoder(16#2a#)) OR
 					(reg_q522 AND symb_decoder(16#42#)) OR
 					(reg_q522 AND symb_decoder(16#e3#)) OR
 					(reg_q522 AND symb_decoder(16#7d#)) OR
 					(reg_q522 AND symb_decoder(16#9c#)) OR
 					(reg_q522 AND symb_decoder(16#fc#)) OR
 					(reg_q522 AND symb_decoder(16#5e#)) OR
 					(reg_q522 AND symb_decoder(16#f7#)) OR
 					(reg_q522 AND symb_decoder(16#f8#)) OR
 					(reg_q522 AND symb_decoder(16#e8#)) OR
 					(reg_q522 AND symb_decoder(16#c8#)) OR
 					(reg_q522 AND symb_decoder(16#49#)) OR
 					(reg_q522 AND symb_decoder(16#92#)) OR
 					(reg_q522 AND symb_decoder(16#98#)) OR
 					(reg_q522 AND symb_decoder(16#6e#)) OR
 					(reg_q522 AND symb_decoder(16#5f#)) OR
 					(reg_q522 AND symb_decoder(16#9e#)) OR
 					(reg_q522 AND symb_decoder(16#40#)) OR
 					(reg_q522 AND symb_decoder(16#1a#)) OR
 					(reg_q522 AND symb_decoder(16#78#)) OR
 					(reg_q522 AND symb_decoder(16#35#)) OR
 					(reg_q522 AND symb_decoder(16#83#)) OR
 					(reg_q522 AND symb_decoder(16#a2#)) OR
 					(reg_q522 AND symb_decoder(16#90#)) OR
 					(reg_q522 AND symb_decoder(16#36#)) OR
 					(reg_q522 AND symb_decoder(16#a8#)) OR
 					(reg_q522 AND symb_decoder(16#24#)) OR
 					(reg_q522 AND symb_decoder(16#17#)) OR
 					(reg_q522 AND symb_decoder(16#5c#)) OR
 					(reg_q522 AND symb_decoder(16#69#)) OR
 					(reg_q522 AND symb_decoder(16#0b#)) OR
 					(reg_q522 AND symb_decoder(16#85#)) OR
 					(reg_q522 AND symb_decoder(16#51#)) OR
 					(reg_q522 AND symb_decoder(16#16#)) OR
 					(reg_q522 AND symb_decoder(16#95#)) OR
 					(reg_q522 AND symb_decoder(16#13#)) OR
 					(reg_q522 AND symb_decoder(16#50#)) OR
 					(reg_q522 AND symb_decoder(16#58#)) OR
 					(reg_q522 AND symb_decoder(16#f6#)) OR
 					(reg_q522 AND symb_decoder(16#94#)) OR
 					(reg_q522 AND symb_decoder(16#4a#)) OR
 					(reg_q522 AND symb_decoder(16#dd#)) OR
 					(reg_q522 AND symb_decoder(16#dc#)) OR
 					(reg_q522 AND symb_decoder(16#de#)) OR
 					(reg_q522 AND symb_decoder(16#ec#)) OR
 					(reg_q522 AND symb_decoder(16#86#)) OR
 					(reg_q522 AND symb_decoder(16#81#)) OR
 					(reg_q522 AND symb_decoder(16#9a#)) OR
 					(reg_q522 AND symb_decoder(16#d5#)) OR
 					(reg_q522 AND symb_decoder(16#cf#)) OR
 					(reg_q522 AND symb_decoder(16#18#)) OR
 					(reg_q522 AND symb_decoder(16#31#)) OR
 					(reg_q522 AND symb_decoder(16#04#)) OR
 					(reg_q522 AND symb_decoder(16#d8#)) OR
 					(reg_q522 AND symb_decoder(16#8d#)) OR
 					(reg_q522 AND symb_decoder(16#15#)) OR
 					(reg_q522 AND symb_decoder(16#bc#)) OR
 					(reg_q522 AND symb_decoder(16#fa#)) OR
 					(reg_q522 AND symb_decoder(16#66#)) OR
 					(reg_q522 AND symb_decoder(16#2f#)) OR
 					(reg_q522 AND symb_decoder(16#e9#)) OR
 					(reg_q522 AND symb_decoder(16#7c#)) OR
 					(reg_q522 AND symb_decoder(16#d7#)) OR
 					(reg_q522 AND symb_decoder(16#07#)) OR
 					(reg_q522 AND symb_decoder(16#fb#)) OR
 					(reg_q522 AND symb_decoder(16#6b#)) OR
 					(reg_q522 AND symb_decoder(16#a9#)) OR
 					(reg_q522 AND symb_decoder(16#30#)) OR
 					(reg_q522 AND symb_decoder(16#14#)) OR
 					(reg_q522 AND symb_decoder(16#6d#)) OR
 					(reg_q522 AND symb_decoder(16#6a#)) OR
 					(reg_q522 AND symb_decoder(16#b1#)) OR
 					(reg_q522 AND symb_decoder(16#4b#)) OR
 					(reg_q522 AND symb_decoder(16#4d#)) OR
 					(reg_q522 AND symb_decoder(16#27#)) OR
 					(reg_q522 AND symb_decoder(16#c1#)) OR
 					(reg_q522 AND symb_decoder(16#be#)) OR
 					(reg_q522 AND symb_decoder(16#99#)) OR
 					(reg_q522 AND symb_decoder(16#77#)) OR
 					(reg_q522 AND symb_decoder(16#cd#)) OR
 					(reg_q522 AND symb_decoder(16#1c#)) OR
 					(reg_q522 AND symb_decoder(16#f5#)) OR
 					(reg_q522 AND symb_decoder(16#9d#)) OR
 					(reg_q522 AND symb_decoder(16#eb#)) OR
 					(reg_q522 AND symb_decoder(16#93#)) OR
 					(reg_q522 AND symb_decoder(16#d3#)) OR
 					(reg_q522 AND symb_decoder(16#8b#)) OR
 					(reg_q522 AND symb_decoder(16#a1#)) OR
 					(reg_q522 AND symb_decoder(16#db#)) OR
 					(reg_q522 AND symb_decoder(16#c9#)) OR
 					(reg_q522 AND symb_decoder(16#73#)) OR
 					(reg_q522 AND symb_decoder(16#5d#)) OR
 					(reg_q522 AND symb_decoder(16#0f#)) OR
 					(reg_q522 AND symb_decoder(16#3d#)) OR
 					(reg_q522 AND symb_decoder(16#ae#)) OR
 					(reg_q522 AND symb_decoder(16#2b#)) OR
 					(reg_q522 AND symb_decoder(16#8a#)) OR
 					(reg_q522 AND symb_decoder(16#c3#)) OR
 					(reg_q522 AND symb_decoder(16#28#)) OR
 					(reg_q522 AND symb_decoder(16#26#)) OR
 					(reg_q522 AND symb_decoder(16#91#)) OR
 					(reg_q522 AND symb_decoder(16#29#)) OR
 					(reg_q522 AND symb_decoder(16#bb#)) OR
 					(reg_q522 AND symb_decoder(16#9b#)) OR
 					(reg_q522 AND symb_decoder(16#b6#)) OR
 					(reg_q522 AND symb_decoder(16#b5#)) OR
 					(reg_q522 AND symb_decoder(16#1d#)) OR
 					(reg_q522 AND symb_decoder(16#0c#)) OR
 					(reg_q522 AND symb_decoder(16#b7#)) OR
 					(reg_q522 AND symb_decoder(16#e0#)) OR
 					(reg_q522 AND symb_decoder(16#f1#)) OR
 					(reg_q522 AND symb_decoder(16#a4#)) OR
 					(reg_q522 AND symb_decoder(16#fe#)) OR
 					(reg_q522 AND symb_decoder(16#3c#)) OR
 					(reg_q522 AND symb_decoder(16#e5#)) OR
 					(reg_q522 AND symb_decoder(16#d1#)) OR
 					(reg_q522 AND symb_decoder(16#ad#)) OR
 					(reg_q522 AND symb_decoder(16#df#)) OR
 					(reg_q522 AND symb_decoder(16#f2#)) OR
 					(reg_q522 AND symb_decoder(16#c7#)) OR
 					(reg_q522 AND symb_decoder(16#06#)) OR
 					(reg_q522 AND symb_decoder(16#00#)) OR
 					(reg_q522 AND symb_decoder(16#b4#)) OR
 					(reg_q522 AND symb_decoder(16#20#)) OR
 					(reg_q522 AND symb_decoder(16#f3#)) OR
 					(reg_q522 AND symb_decoder(16#62#)) OR
 					(reg_q522 AND symb_decoder(16#5b#)) OR
 					(reg_q522 AND symb_decoder(16#3b#)) OR
 					(reg_q522 AND symb_decoder(16#57#)) OR
 					(reg_q522 AND symb_decoder(16#59#)) OR
 					(reg_q522 AND symb_decoder(16#bd#)) OR
 					(reg_q522 AND symb_decoder(16#80#)) OR
 					(reg_q522 AND symb_decoder(16#4f#)) OR
 					(reg_q522 AND symb_decoder(16#d4#)) OR
 					(reg_q522 AND symb_decoder(16#f9#)) OR
 					(reg_q522 AND symb_decoder(16#7e#)) OR
 					(reg_q522 AND symb_decoder(16#ee#)) OR
 					(reg_q522 AND symb_decoder(16#76#)) OR
 					(reg_q522 AND symb_decoder(16#61#)) OR
 					(reg_q522 AND symb_decoder(16#7f#)) OR
 					(reg_q522 AND symb_decoder(16#c0#)) OR
 					(reg_q522 AND symb_decoder(16#b8#)) OR
 					(reg_q522 AND symb_decoder(16#56#)) OR
 					(reg_q522 AND symb_decoder(16#7a#)) OR
 					(reg_q522 AND symb_decoder(16#89#)) OR
 					(reg_q522 AND symb_decoder(16#a0#)) OR
 					(reg_q522 AND symb_decoder(16#45#)) OR
 					(reg_q522 AND symb_decoder(16#8f#)) OR
 					(reg_q522 AND symb_decoder(16#c2#)) OR
 					(reg_q522 AND symb_decoder(16#43#)) OR
 					(reg_q522 AND symb_decoder(16#46#)) OR
 					(reg_q522 AND symb_decoder(16#09#)) OR
 					(reg_q522 AND symb_decoder(16#05#)) OR
 					(reg_q522 AND symb_decoder(16#3f#)) OR
 					(reg_q522 AND symb_decoder(16#7b#)) OR
 					(reg_q522 AND symb_decoder(16#1b#)) OR
 					(reg_q522 AND symb_decoder(16#d2#)) OR
 					(reg_q522 AND symb_decoder(16#71#)) OR
 					(reg_q522 AND symb_decoder(16#84#)) OR
 					(reg_q522 AND symb_decoder(16#c4#)) OR
 					(reg_q522 AND symb_decoder(16#8c#)) OR
 					(reg_q522 AND symb_decoder(16#65#)) OR
 					(reg_q522 AND symb_decoder(16#b0#)) OR
 					(reg_q522 AND symb_decoder(16#a3#)) OR
 					(reg_q522 AND symb_decoder(16#63#)) OR
 					(reg_q522 AND symb_decoder(16#3a#)) OR
 					(reg_q522 AND symb_decoder(16#55#)) OR
 					(reg_q522 AND symb_decoder(16#b3#)) OR
 					(reg_q522 AND symb_decoder(16#b9#)) OR
 					(reg_q522 AND symb_decoder(16#02#)) OR
 					(reg_q522 AND symb_decoder(16#a7#)) OR
 					(reg_q522 AND symb_decoder(16#ac#)) OR
 					(reg_q522 AND symb_decoder(16#c5#)) OR
 					(reg_q522 AND symb_decoder(16#25#)) OR
 					(reg_q522 AND symb_decoder(16#33#)) OR
 					(reg_q522 AND symb_decoder(16#e1#)) OR
 					(reg_q522 AND symb_decoder(16#ca#)) OR
 					(reg_q522 AND symb_decoder(16#67#)) OR
 					(reg_q522 AND symb_decoder(16#38#)) OR
 					(reg_q522 AND symb_decoder(16#39#)) OR
 					(reg_q522 AND symb_decoder(16#af#)) OR
 					(reg_q522 AND symb_decoder(16#54#)) OR
 					(reg_q522 AND symb_decoder(16#12#)) OR
 					(reg_q522 AND symb_decoder(16#44#)) OR
 					(reg_q522 AND symb_decoder(16#37#)) OR
 					(reg_q522 AND symb_decoder(16#2c#)) OR
 					(reg_q522 AND symb_decoder(16#ba#)) OR
 					(reg_q522 AND symb_decoder(16#08#)) OR
 					(reg_q522 AND symb_decoder(16#e2#)) OR
 					(reg_q522 AND symb_decoder(16#97#)) OR
 					(reg_q522 AND symb_decoder(16#88#)) OR
 					(reg_q522 AND symb_decoder(16#ea#)) OR
 					(reg_q522 AND symb_decoder(16#21#)) OR
 					(reg_q522 AND symb_decoder(16#2e#)) OR
 					(reg_q522 AND symb_decoder(16#ce#)) OR
 					(reg_q522 AND symb_decoder(16#72#)) OR
 					(reg_q522 AND symb_decoder(16#82#)) OR
 					(reg_q522 AND symb_decoder(16#19#)) OR
 					(reg_q522 AND symb_decoder(16#53#)) OR
 					(reg_q522 AND symb_decoder(16#f0#)) OR
 					(reg_q522 AND symb_decoder(16#96#)) OR
 					(reg_q522 AND symb_decoder(16#c6#)) OR
 					(reg_q522 AND symb_decoder(16#4e#)) OR
 					(reg_q522 AND symb_decoder(16#4c#)) OR
 					(reg_q522 AND symb_decoder(16#1f#)) OR
 					(reg_q522 AND symb_decoder(16#d9#)) OR
 					(reg_q522 AND symb_decoder(16#87#)) OR
 					(reg_q522 AND symb_decoder(16#fd#)) OR
 					(reg_q522 AND symb_decoder(16#23#)) OR
 					(reg_q522 AND symb_decoder(16#03#)) OR
 					(reg_q522 AND symb_decoder(16#aa#)) OR
 					(reg_q522 AND symb_decoder(16#75#)) OR
 					(reg_q522 AND symb_decoder(16#d6#)) OR
 					(reg_q522 AND symb_decoder(16#9f#)) OR
 					(reg_q522 AND symb_decoder(16#a6#)) OR
 					(reg_q522 AND symb_decoder(16#b2#)) OR
 					(reg_q522 AND symb_decoder(16#74#)) OR
 					(reg_q522 AND symb_decoder(16#48#)) OR
 					(reg_q522 AND symb_decoder(16#f4#)) OR
 					(reg_q522 AND symb_decoder(16#32#)) OR
 					(reg_q522 AND symb_decoder(16#cb#)) OR
 					(reg_q522 AND symb_decoder(16#6c#)) OR
 					(reg_q542 AND symb_decoder(16#14#)) OR
 					(reg_q542 AND symb_decoder(16#03#)) OR
 					(reg_q542 AND symb_decoder(16#89#)) OR
 					(reg_q542 AND symb_decoder(16#58#)) OR
 					(reg_q542 AND symb_decoder(16#95#)) OR
 					(reg_q542 AND symb_decoder(16#0f#)) OR
 					(reg_q542 AND symb_decoder(16#45#)) OR
 					(reg_q542 AND symb_decoder(16#8a#)) OR
 					(reg_q542 AND symb_decoder(16#f0#)) OR
 					(reg_q542 AND symb_decoder(16#d5#)) OR
 					(reg_q542 AND symb_decoder(16#75#)) OR
 					(reg_q542 AND symb_decoder(16#91#)) OR
 					(reg_q542 AND symb_decoder(16#1b#)) OR
 					(reg_q542 AND symb_decoder(16#d8#)) OR
 					(reg_q542 AND symb_decoder(16#5e#)) OR
 					(reg_q542 AND symb_decoder(16#cd#)) OR
 					(reg_q542 AND symb_decoder(16#27#)) OR
 					(reg_q542 AND symb_decoder(16#10#)) OR
 					(reg_q542 AND symb_decoder(16#dd#)) OR
 					(reg_q542 AND symb_decoder(16#b2#)) OR
 					(reg_q542 AND symb_decoder(16#1f#)) OR
 					(reg_q542 AND symb_decoder(16#4c#)) OR
 					(reg_q542 AND symb_decoder(16#c2#)) OR
 					(reg_q542 AND symb_decoder(16#2a#)) OR
 					(reg_q542 AND symb_decoder(16#07#)) OR
 					(reg_q542 AND symb_decoder(16#39#)) OR
 					(reg_q542 AND symb_decoder(16#f4#)) OR
 					(reg_q542 AND symb_decoder(16#8e#)) OR
 					(reg_q542 AND symb_decoder(16#46#)) OR
 					(reg_q542 AND symb_decoder(16#61#)) OR
 					(reg_q542 AND symb_decoder(16#3b#)) OR
 					(reg_q542 AND symb_decoder(16#7f#)) OR
 					(reg_q542 AND symb_decoder(16#4d#)) OR
 					(reg_q542 AND symb_decoder(16#bc#)) OR
 					(reg_q542 AND symb_decoder(16#b7#)) OR
 					(reg_q542 AND symb_decoder(16#5b#)) OR
 					(reg_q542 AND symb_decoder(16#86#)) OR
 					(reg_q542 AND symb_decoder(16#da#)) OR
 					(reg_q542 AND symb_decoder(16#25#)) OR
 					(reg_q542 AND symb_decoder(16#ad#)) OR
 					(reg_q542 AND symb_decoder(16#fe#)) OR
 					(reg_q542 AND symb_decoder(16#9b#)) OR
 					(reg_q542 AND symb_decoder(16#21#)) OR
 					(reg_q542 AND symb_decoder(16#5c#)) OR
 					(reg_q542 AND symb_decoder(16#8b#)) OR
 					(reg_q542 AND symb_decoder(16#b1#)) OR
 					(reg_q542 AND symb_decoder(16#34#)) OR
 					(reg_q542 AND symb_decoder(16#4b#)) OR
 					(reg_q542 AND symb_decoder(16#55#)) OR
 					(reg_q542 AND symb_decoder(16#24#)) OR
 					(reg_q542 AND symb_decoder(16#70#)) OR
 					(reg_q542 AND symb_decoder(16#ec#)) OR
 					(reg_q542 AND symb_decoder(16#82#)) OR
 					(reg_q542 AND symb_decoder(16#17#)) OR
 					(reg_q542 AND symb_decoder(16#ed#)) OR
 					(reg_q542 AND symb_decoder(16#c9#)) OR
 					(reg_q542 AND symb_decoder(16#19#)) OR
 					(reg_q542 AND symb_decoder(16#59#)) OR
 					(reg_q542 AND symb_decoder(16#d2#)) OR
 					(reg_q542 AND symb_decoder(16#2b#)) OR
 					(reg_q542 AND symb_decoder(16#5d#)) OR
 					(reg_q542 AND symb_decoder(16#13#)) OR
 					(reg_q542 AND symb_decoder(16#5f#)) OR
 					(reg_q542 AND symb_decoder(16#08#)) OR
 					(reg_q542 AND symb_decoder(16#7d#)) OR
 					(reg_q542 AND symb_decoder(16#3d#)) OR
 					(reg_q542 AND symb_decoder(16#64#)) OR
 					(reg_q542 AND symb_decoder(16#a1#)) OR
 					(reg_q542 AND symb_decoder(16#e7#)) OR
 					(reg_q542 AND symb_decoder(16#bf#)) OR
 					(reg_q542 AND symb_decoder(16#69#)) OR
 					(reg_q542 AND symb_decoder(16#dc#)) OR
 					(reg_q542 AND symb_decoder(16#0c#)) OR
 					(reg_q542 AND symb_decoder(16#e6#)) OR
 					(reg_q542 AND symb_decoder(16#33#)) OR
 					(reg_q542 AND symb_decoder(16#35#)) OR
 					(reg_q542 AND symb_decoder(16#e0#)) OR
 					(reg_q542 AND symb_decoder(16#f1#)) OR
 					(reg_q542 AND symb_decoder(16#88#)) OR
 					(reg_q542 AND symb_decoder(16#b0#)) OR
 					(reg_q542 AND symb_decoder(16#2f#)) OR
 					(reg_q542 AND symb_decoder(16#9f#)) OR
 					(reg_q542 AND symb_decoder(16#62#)) OR
 					(reg_q542 AND symb_decoder(16#81#)) OR
 					(reg_q542 AND symb_decoder(16#52#)) OR
 					(reg_q542 AND symb_decoder(16#1c#)) OR
 					(reg_q542 AND symb_decoder(16#6e#)) OR
 					(reg_q542 AND symb_decoder(16#a7#)) OR
 					(reg_q542 AND symb_decoder(16#3f#)) OR
 					(reg_q542 AND symb_decoder(16#47#)) OR
 					(reg_q542 AND symb_decoder(16#e8#)) OR
 					(reg_q542 AND symb_decoder(16#6a#)) OR
 					(reg_q542 AND symb_decoder(16#22#)) OR
 					(reg_q542 AND symb_decoder(16#2e#)) OR
 					(reg_q542 AND symb_decoder(16#6c#)) OR
 					(reg_q542 AND symb_decoder(16#cb#)) OR
 					(reg_q542 AND symb_decoder(16#f6#)) OR
 					(reg_q542 AND symb_decoder(16#15#)) OR
 					(reg_q542 AND symb_decoder(16#74#)) OR
 					(reg_q542 AND symb_decoder(16#eb#)) OR
 					(reg_q542 AND symb_decoder(16#31#)) OR
 					(reg_q542 AND symb_decoder(16#d9#)) OR
 					(reg_q542 AND symb_decoder(16#01#)) OR
 					(reg_q542 AND symb_decoder(16#66#)) OR
 					(reg_q542 AND symb_decoder(16#40#)) OR
 					(reg_q542 AND symb_decoder(16#f2#)) OR
 					(reg_q542 AND symb_decoder(16#98#)) OR
 					(reg_q542 AND symb_decoder(16#c5#)) OR
 					(reg_q542 AND symb_decoder(16#be#)) OR
 					(reg_q542 AND symb_decoder(16#50#)) OR
 					(reg_q542 AND symb_decoder(16#cc#)) OR
 					(reg_q542 AND symb_decoder(16#cf#)) OR
 					(reg_q542 AND symb_decoder(16#a4#)) OR
 					(reg_q542 AND symb_decoder(16#3c#)) OR
 					(reg_q542 AND symb_decoder(16#b9#)) OR
 					(reg_q542 AND symb_decoder(16#73#)) OR
 					(reg_q542 AND symb_decoder(16#a5#)) OR
 					(reg_q542 AND symb_decoder(16#ab#)) OR
 					(reg_q542 AND symb_decoder(16#2c#)) OR
 					(reg_q542 AND symb_decoder(16#e2#)) OR
 					(reg_q542 AND symb_decoder(16#ba#)) OR
 					(reg_q542 AND symb_decoder(16#8d#)) OR
 					(reg_q542 AND symb_decoder(16#8f#)) OR
 					(reg_q542 AND symb_decoder(16#d7#)) OR
 					(reg_q542 AND symb_decoder(16#1e#)) OR
 					(reg_q542 AND symb_decoder(16#00#)) OR
 					(reg_q542 AND symb_decoder(16#f9#)) OR
 					(reg_q542 AND symb_decoder(16#4e#)) OR
 					(reg_q542 AND symb_decoder(16#68#)) OR
 					(reg_q542 AND symb_decoder(16#80#)) OR
 					(reg_q542 AND symb_decoder(16#6b#)) OR
 					(reg_q542 AND symb_decoder(16#2d#)) OR
 					(reg_q542 AND symb_decoder(16#ef#)) OR
 					(reg_q542 AND symb_decoder(16#aa#)) OR
 					(reg_q542 AND symb_decoder(16#30#)) OR
 					(reg_q542 AND symb_decoder(16#48#)) OR
 					(reg_q542 AND symb_decoder(16#e5#)) OR
 					(reg_q542 AND symb_decoder(16#78#)) OR
 					(reg_q542 AND symb_decoder(16#b3#)) OR
 					(reg_q542 AND symb_decoder(16#ce#)) OR
 					(reg_q542 AND symb_decoder(16#d3#)) OR
 					(reg_q542 AND symb_decoder(16#ae#)) OR
 					(reg_q542 AND symb_decoder(16#76#)) OR
 					(reg_q542 AND symb_decoder(16#85#)) OR
 					(reg_q542 AND symb_decoder(16#23#)) OR
 					(reg_q542 AND symb_decoder(16#0e#)) OR
 					(reg_q542 AND symb_decoder(16#60#)) OR
 					(reg_q542 AND symb_decoder(16#e1#)) OR
 					(reg_q542 AND symb_decoder(16#1d#)) OR
 					(reg_q542 AND symb_decoder(16#a8#)) OR
 					(reg_q542 AND symb_decoder(16#3a#)) OR
 					(reg_q542 AND symb_decoder(16#9c#)) OR
 					(reg_q542 AND symb_decoder(16#fc#)) OR
 					(reg_q542 AND symb_decoder(16#a9#)) OR
 					(reg_q542 AND symb_decoder(16#51#)) OR
 					(reg_q542 AND symb_decoder(16#ff#)) OR
 					(reg_q542 AND symb_decoder(16#9a#)) OR
 					(reg_q542 AND symb_decoder(16#57#)) OR
 					(reg_q542 AND symb_decoder(16#49#)) OR
 					(reg_q542 AND symb_decoder(16#c7#)) OR
 					(reg_q542 AND symb_decoder(16#11#)) OR
 					(reg_q542 AND symb_decoder(16#f5#)) OR
 					(reg_q542 AND symb_decoder(16#d4#)) OR
 					(reg_q542 AND symb_decoder(16#f8#)) OR
 					(reg_q542 AND symb_decoder(16#5a#)) OR
 					(reg_q542 AND symb_decoder(16#bb#)) OR
 					(reg_q542 AND symb_decoder(16#20#)) OR
 					(reg_q542 AND symb_decoder(16#32#)) OR
 					(reg_q542 AND symb_decoder(16#8c#)) OR
 					(reg_q542 AND symb_decoder(16#97#)) OR
 					(reg_q542 AND symb_decoder(16#67#)) OR
 					(reg_q542 AND symb_decoder(16#de#)) OR
 					(reg_q542 AND symb_decoder(16#d6#)) OR
 					(reg_q542 AND symb_decoder(16#94#)) OR
 					(reg_q542 AND symb_decoder(16#29#)) OR
 					(reg_q542 AND symb_decoder(16#a6#)) OR
 					(reg_q542 AND symb_decoder(16#a2#)) OR
 					(reg_q542 AND symb_decoder(16#9e#)) OR
 					(reg_q542 AND symb_decoder(16#b6#)) OR
 					(reg_q542 AND symb_decoder(16#65#)) OR
 					(reg_q542 AND symb_decoder(16#b8#)) OR
 					(reg_q542 AND symb_decoder(16#b5#)) OR
 					(reg_q542 AND symb_decoder(16#f3#)) OR
 					(reg_q542 AND symb_decoder(16#ea#)) OR
 					(reg_q542 AND symb_decoder(16#d0#)) OR
 					(reg_q542 AND symb_decoder(16#c6#)) OR
 					(reg_q542 AND symb_decoder(16#fd#)) OR
 					(reg_q542 AND symb_decoder(16#3e#)) OR
 					(reg_q542 AND symb_decoder(16#a3#)) OR
 					(reg_q542 AND symb_decoder(16#6f#)) OR
 					(reg_q542 AND symb_decoder(16#c1#)) OR
 					(reg_q542 AND symb_decoder(16#79#)) OR
 					(reg_q542 AND symb_decoder(16#84#)) OR
 					(reg_q542 AND symb_decoder(16#54#)) OR
 					(reg_q542 AND symb_decoder(16#6d#)) OR
 					(reg_q542 AND symb_decoder(16#77#)) OR
 					(reg_q542 AND symb_decoder(16#72#)) OR
 					(reg_q542 AND symb_decoder(16#37#)) OR
 					(reg_q542 AND symb_decoder(16#c0#)) OR
 					(reg_q542 AND symb_decoder(16#28#)) OR
 					(reg_q542 AND symb_decoder(16#38#)) OR
 					(reg_q542 AND symb_decoder(16#fb#)) OR
 					(reg_q542 AND symb_decoder(16#56#)) OR
 					(reg_q542 AND symb_decoder(16#ee#)) OR
 					(reg_q542 AND symb_decoder(16#c3#)) OR
 					(reg_q542 AND symb_decoder(16#63#)) OR
 					(reg_q542 AND symb_decoder(16#05#)) OR
 					(reg_q542 AND symb_decoder(16#83#)) OR
 					(reg_q542 AND symb_decoder(16#87#)) OR
 					(reg_q542 AND symb_decoder(16#bd#)) OR
 					(reg_q542 AND symb_decoder(16#ac#)) OR
 					(reg_q542 AND symb_decoder(16#09#)) OR
 					(reg_q542 AND symb_decoder(16#7e#)) OR
 					(reg_q542 AND symb_decoder(16#06#)) OR
 					(reg_q542 AND symb_decoder(16#92#)) OR
 					(reg_q542 AND symb_decoder(16#ca#)) OR
 					(reg_q542 AND symb_decoder(16#26#)) OR
 					(reg_q542 AND symb_decoder(16#41#)) OR
 					(reg_q542 AND symb_decoder(16#42#)) OR
 					(reg_q542 AND symb_decoder(16#e4#)) OR
 					(reg_q542 AND symb_decoder(16#a0#)) OR
 					(reg_q542 AND symb_decoder(16#c4#)) OR
 					(reg_q542 AND symb_decoder(16#18#)) OR
 					(reg_q542 AND symb_decoder(16#e3#)) OR
 					(reg_q542 AND symb_decoder(16#e9#)) OR
 					(reg_q542 AND symb_decoder(16#7b#)) OR
 					(reg_q542 AND symb_decoder(16#99#)) OR
 					(reg_q542 AND symb_decoder(16#53#)) OR
 					(reg_q542 AND symb_decoder(16#db#)) OR
 					(reg_q542 AND symb_decoder(16#93#)) OR
 					(reg_q542 AND symb_decoder(16#0b#)) OR
 					(reg_q542 AND symb_decoder(16#df#)) OR
 					(reg_q542 AND symb_decoder(16#43#)) OR
 					(reg_q542 AND symb_decoder(16#44#)) OR
 					(reg_q542 AND symb_decoder(16#b4#)) OR
 					(reg_q542 AND symb_decoder(16#f7#)) OR
 					(reg_q542 AND symb_decoder(16#fa#)) OR
 					(reg_q542 AND symb_decoder(16#c8#)) OR
 					(reg_q542 AND symb_decoder(16#4a#)) OR
 					(reg_q542 AND symb_decoder(16#16#)) OR
 					(reg_q542 AND symb_decoder(16#9d#)) OR
 					(reg_q542 AND symb_decoder(16#1a#)) OR
 					(reg_q542 AND symb_decoder(16#d1#)) OR
 					(reg_q542 AND symb_decoder(16#12#)) OR
 					(reg_q542 AND symb_decoder(16#4f#)) OR
 					(reg_q542 AND symb_decoder(16#04#)) OR
 					(reg_q542 AND symb_decoder(16#96#)) OR
 					(reg_q542 AND symb_decoder(16#7c#)) OR
 					(reg_q542 AND symb_decoder(16#7a#)) OR
 					(reg_q542 AND symb_decoder(16#af#)) OR
 					(reg_q542 AND symb_decoder(16#90#)) OR
 					(reg_q542 AND symb_decoder(16#02#)) OR
 					(reg_q542 AND symb_decoder(16#36#)) OR
 					(reg_q542 AND symb_decoder(16#71#));
reg_q857_in <= (reg_q819 AND symb_decoder(16#17#)) OR
 					(reg_q819 AND symb_decoder(16#98#)) OR
 					(reg_q819 AND symb_decoder(16#7f#)) OR
 					(reg_q819 AND symb_decoder(16#93#)) OR
 					(reg_q819 AND symb_decoder(16#b4#)) OR
 					(reg_q819 AND symb_decoder(16#ca#)) OR
 					(reg_q819 AND symb_decoder(16#6c#)) OR
 					(reg_q819 AND symb_decoder(16#43#)) OR
 					(reg_q819 AND symb_decoder(16#31#)) OR
 					(reg_q819 AND symb_decoder(16#72#)) OR
 					(reg_q819 AND symb_decoder(16#e6#)) OR
 					(reg_q819 AND symb_decoder(16#8e#)) OR
 					(reg_q819 AND symb_decoder(16#68#)) OR
 					(reg_q819 AND symb_decoder(16#40#)) OR
 					(reg_q819 AND symb_decoder(16#ff#)) OR
 					(reg_q819 AND symb_decoder(16#1f#)) OR
 					(reg_q819 AND symb_decoder(16#3c#)) OR
 					(reg_q819 AND symb_decoder(16#df#)) OR
 					(reg_q819 AND symb_decoder(16#ef#)) OR
 					(reg_q819 AND symb_decoder(16#b7#)) OR
 					(reg_q819 AND symb_decoder(16#9d#)) OR
 					(reg_q819 AND symb_decoder(16#0f#)) OR
 					(reg_q819 AND symb_decoder(16#29#)) OR
 					(reg_q819 AND symb_decoder(16#c6#)) OR
 					(reg_q819 AND symb_decoder(16#7a#)) OR
 					(reg_q819 AND symb_decoder(16#22#)) OR
 					(reg_q819 AND symb_decoder(16#ab#)) OR
 					(reg_q819 AND symb_decoder(16#44#)) OR
 					(reg_q819 AND symb_decoder(16#8a#)) OR
 					(reg_q819 AND symb_decoder(16#0e#)) OR
 					(reg_q819 AND symb_decoder(16#e4#)) OR
 					(reg_q819 AND symb_decoder(16#42#)) OR
 					(reg_q819 AND symb_decoder(16#ac#)) OR
 					(reg_q819 AND symb_decoder(16#73#)) OR
 					(reg_q819 AND symb_decoder(16#c5#)) OR
 					(reg_q819 AND symb_decoder(16#5b#)) OR
 					(reg_q819 AND symb_decoder(16#1a#)) OR
 					(reg_q819 AND symb_decoder(16#c8#)) OR
 					(reg_q819 AND symb_decoder(16#57#)) OR
 					(reg_q819 AND symb_decoder(16#fa#)) OR
 					(reg_q819 AND symb_decoder(16#67#)) OR
 					(reg_q819 AND symb_decoder(16#6d#)) OR
 					(reg_q819 AND symb_decoder(16#7b#)) OR
 					(reg_q819 AND symb_decoder(16#81#)) OR
 					(reg_q819 AND symb_decoder(16#10#)) OR
 					(reg_q819 AND symb_decoder(16#6f#)) OR
 					(reg_q819 AND symb_decoder(16#ec#)) OR
 					(reg_q819 AND symb_decoder(16#00#)) OR
 					(reg_q819 AND symb_decoder(16#85#)) OR
 					(reg_q819 AND symb_decoder(16#48#)) OR
 					(reg_q819 AND symb_decoder(16#90#)) OR
 					(reg_q819 AND symb_decoder(16#e3#)) OR
 					(reg_q819 AND symb_decoder(16#59#)) OR
 					(reg_q819 AND symb_decoder(16#08#)) OR
 					(reg_q819 AND symb_decoder(16#ed#)) OR
 					(reg_q819 AND symb_decoder(16#dd#)) OR
 					(reg_q819 AND symb_decoder(16#09#)) OR
 					(reg_q819 AND symb_decoder(16#88#)) OR
 					(reg_q819 AND symb_decoder(16#d8#)) OR
 					(reg_q819 AND symb_decoder(16#02#)) OR
 					(reg_q819 AND symb_decoder(16#30#)) OR
 					(reg_q819 AND symb_decoder(16#f1#)) OR
 					(reg_q819 AND symb_decoder(16#f7#)) OR
 					(reg_q819 AND symb_decoder(16#5d#)) OR
 					(reg_q819 AND symb_decoder(16#db#)) OR
 					(reg_q819 AND symb_decoder(16#58#)) OR
 					(reg_q819 AND symb_decoder(16#3b#)) OR
 					(reg_q819 AND symb_decoder(16#28#)) OR
 					(reg_q819 AND symb_decoder(16#fe#)) OR
 					(reg_q819 AND symb_decoder(16#d0#)) OR
 					(reg_q819 AND symb_decoder(16#69#)) OR
 					(reg_q819 AND symb_decoder(16#24#)) OR
 					(reg_q819 AND symb_decoder(16#2a#)) OR
 					(reg_q819 AND symb_decoder(16#f3#)) OR
 					(reg_q819 AND symb_decoder(16#a1#)) OR
 					(reg_q819 AND symb_decoder(16#60#)) OR
 					(reg_q819 AND symb_decoder(16#49#)) OR
 					(reg_q819 AND symb_decoder(16#ea#)) OR
 					(reg_q819 AND symb_decoder(16#1d#)) OR
 					(reg_q819 AND symb_decoder(16#91#)) OR
 					(reg_q819 AND symb_decoder(16#11#)) OR
 					(reg_q819 AND symb_decoder(16#18#)) OR
 					(reg_q819 AND symb_decoder(16#2b#)) OR
 					(reg_q819 AND symb_decoder(16#7d#)) OR
 					(reg_q819 AND symb_decoder(16#76#)) OR
 					(reg_q819 AND symb_decoder(16#bb#)) OR
 					(reg_q819 AND symb_decoder(16#c0#)) OR
 					(reg_q819 AND symb_decoder(16#b2#)) OR
 					(reg_q819 AND symb_decoder(16#92#)) OR
 					(reg_q819 AND symb_decoder(16#b6#)) OR
 					(reg_q819 AND symb_decoder(16#c4#)) OR
 					(reg_q819 AND symb_decoder(16#53#)) OR
 					(reg_q819 AND symb_decoder(16#d4#)) OR
 					(reg_q819 AND symb_decoder(16#e1#)) OR
 					(reg_q819 AND symb_decoder(16#a5#)) OR
 					(reg_q819 AND symb_decoder(16#ce#)) OR
 					(reg_q819 AND symb_decoder(16#ae#)) OR
 					(reg_q819 AND symb_decoder(16#2e#)) OR
 					(reg_q819 AND symb_decoder(16#a7#)) OR
 					(reg_q819 AND symb_decoder(16#a9#)) OR
 					(reg_q819 AND symb_decoder(16#47#)) OR
 					(reg_q819 AND symb_decoder(16#1b#)) OR
 					(reg_q819 AND symb_decoder(16#5a#)) OR
 					(reg_q819 AND symb_decoder(16#63#)) OR
 					(reg_q819 AND symb_decoder(16#a0#)) OR
 					(reg_q819 AND symb_decoder(16#4f#)) OR
 					(reg_q819 AND symb_decoder(16#de#)) OR
 					(reg_q819 AND symb_decoder(16#0c#)) OR
 					(reg_q819 AND symb_decoder(16#46#)) OR
 					(reg_q819 AND symb_decoder(16#3a#)) OR
 					(reg_q819 AND symb_decoder(16#97#)) OR
 					(reg_q819 AND symb_decoder(16#da#)) OR
 					(reg_q819 AND symb_decoder(16#eb#)) OR
 					(reg_q819 AND symb_decoder(16#5e#)) OR
 					(reg_q819 AND symb_decoder(16#33#)) OR
 					(reg_q819 AND symb_decoder(16#64#)) OR
 					(reg_q819 AND symb_decoder(16#50#)) OR
 					(reg_q819 AND symb_decoder(16#e0#)) OR
 					(reg_q819 AND symb_decoder(16#c1#)) OR
 					(reg_q819 AND symb_decoder(16#75#)) OR
 					(reg_q819 AND symb_decoder(16#ee#)) OR
 					(reg_q819 AND symb_decoder(16#12#)) OR
 					(reg_q819 AND symb_decoder(16#d3#)) OR
 					(reg_q819 AND symb_decoder(16#b0#)) OR
 					(reg_q819 AND symb_decoder(16#b5#)) OR
 					(reg_q819 AND symb_decoder(16#04#)) OR
 					(reg_q819 AND symb_decoder(16#77#)) OR
 					(reg_q819 AND symb_decoder(16#52#)) OR
 					(reg_q819 AND symb_decoder(16#86#)) OR
 					(reg_q819 AND symb_decoder(16#14#)) OR
 					(reg_q819 AND symb_decoder(16#d1#)) OR
 					(reg_q819 AND symb_decoder(16#d2#)) OR
 					(reg_q819 AND symb_decoder(16#38#)) OR
 					(reg_q819 AND symb_decoder(16#ba#)) OR
 					(reg_q819 AND symb_decoder(16#45#)) OR
 					(reg_q819 AND symb_decoder(16#70#)) OR
 					(reg_q819 AND symb_decoder(16#3e#)) OR
 					(reg_q819 AND symb_decoder(16#55#)) OR
 					(reg_q819 AND symb_decoder(16#20#)) OR
 					(reg_q819 AND symb_decoder(16#82#)) OR
 					(reg_q819 AND symb_decoder(16#e2#)) OR
 					(reg_q819 AND symb_decoder(16#4a#)) OR
 					(reg_q819 AND symb_decoder(16#26#)) OR
 					(reg_q819 AND symb_decoder(16#84#)) OR
 					(reg_q819 AND symb_decoder(16#ad#)) OR
 					(reg_q819 AND symb_decoder(16#af#)) OR
 					(reg_q819 AND symb_decoder(16#87#)) OR
 					(reg_q819 AND symb_decoder(16#f6#)) OR
 					(reg_q819 AND symb_decoder(16#54#)) OR
 					(reg_q819 AND symb_decoder(16#be#)) OR
 					(reg_q819 AND symb_decoder(16#83#)) OR
 					(reg_q819 AND symb_decoder(16#41#)) OR
 					(reg_q819 AND symb_decoder(16#9a#)) OR
 					(reg_q819 AND symb_decoder(16#39#)) OR
 					(reg_q819 AND symb_decoder(16#96#)) OR
 					(reg_q819 AND symb_decoder(16#78#)) OR
 					(reg_q819 AND symb_decoder(16#b9#)) OR
 					(reg_q819 AND symb_decoder(16#9b#)) OR
 					(reg_q819 AND symb_decoder(16#4b#)) OR
 					(reg_q819 AND symb_decoder(16#6b#)) OR
 					(reg_q819 AND symb_decoder(16#9c#)) OR
 					(reg_q819 AND symb_decoder(16#f4#)) OR
 					(reg_q819 AND symb_decoder(16#06#)) OR
 					(reg_q819 AND symb_decoder(16#2d#)) OR
 					(reg_q819 AND symb_decoder(16#36#)) OR
 					(reg_q819 AND symb_decoder(16#d5#)) OR
 					(reg_q819 AND symb_decoder(16#fc#)) OR
 					(reg_q819 AND symb_decoder(16#cc#)) OR
 					(reg_q819 AND symb_decoder(16#c3#)) OR
 					(reg_q819 AND symb_decoder(16#89#)) OR
 					(reg_q819 AND symb_decoder(16#25#)) OR
 					(reg_q819 AND symb_decoder(16#07#)) OR
 					(reg_q819 AND symb_decoder(16#c7#)) OR
 					(reg_q819 AND symb_decoder(16#80#)) OR
 					(reg_q819 AND symb_decoder(16#f9#)) OR
 					(reg_q819 AND symb_decoder(16#51#)) OR
 					(reg_q819 AND symb_decoder(16#5c#)) OR
 					(reg_q819 AND symb_decoder(16#9f#)) OR
 					(reg_q819 AND symb_decoder(16#cb#)) OR
 					(reg_q819 AND symb_decoder(16#95#)) OR
 					(reg_q819 AND symb_decoder(16#c9#)) OR
 					(reg_q819 AND symb_decoder(16#e9#)) OR
 					(reg_q819 AND symb_decoder(16#0b#)) OR
 					(reg_q819 AND symb_decoder(16#c2#)) OR
 					(reg_q819 AND symb_decoder(16#4c#)) OR
 					(reg_q819 AND symb_decoder(16#61#)) OR
 					(reg_q819 AND symb_decoder(16#15#)) OR
 					(reg_q819 AND symb_decoder(16#3d#)) OR
 					(reg_q819 AND symb_decoder(16#16#)) OR
 					(reg_q819 AND symb_decoder(16#37#)) OR
 					(reg_q819 AND symb_decoder(16#79#)) OR
 					(reg_q819 AND symb_decoder(16#e7#)) OR
 					(reg_q819 AND symb_decoder(16#66#)) OR
 					(reg_q819 AND symb_decoder(16#05#)) OR
 					(reg_q819 AND symb_decoder(16#21#)) OR
 					(reg_q819 AND symb_decoder(16#a6#)) OR
 					(reg_q819 AND symb_decoder(16#6e#)) OR
 					(reg_q819 AND symb_decoder(16#6a#)) OR
 					(reg_q819 AND symb_decoder(16#b3#)) OR
 					(reg_q819 AND symb_decoder(16#8c#)) OR
 					(reg_q819 AND symb_decoder(16#7c#)) OR
 					(reg_q819 AND symb_decoder(16#13#)) OR
 					(reg_q819 AND symb_decoder(16#a8#)) OR
 					(reg_q819 AND symb_decoder(16#2f#)) OR
 					(reg_q819 AND symb_decoder(16#99#)) OR
 					(reg_q819 AND symb_decoder(16#bc#)) OR
 					(reg_q819 AND symb_decoder(16#71#)) OR
 					(reg_q819 AND symb_decoder(16#56#)) OR
 					(reg_q819 AND symb_decoder(16#b8#)) OR
 					(reg_q819 AND symb_decoder(16#2c#)) OR
 					(reg_q819 AND symb_decoder(16#7e#)) OR
 					(reg_q819 AND symb_decoder(16#dc#)) OR
 					(reg_q819 AND symb_decoder(16#f5#)) OR
 					(reg_q819 AND symb_decoder(16#fd#)) OR
 					(reg_q819 AND symb_decoder(16#f2#)) OR
 					(reg_q819 AND symb_decoder(16#65#)) OR
 					(reg_q819 AND symb_decoder(16#5f#)) OR
 					(reg_q819 AND symb_decoder(16#e8#)) OR
 					(reg_q819 AND symb_decoder(16#fb#)) OR
 					(reg_q819 AND symb_decoder(16#b1#)) OR
 					(reg_q819 AND symb_decoder(16#19#)) OR
 					(reg_q819 AND symb_decoder(16#4e#)) OR
 					(reg_q819 AND symb_decoder(16#1c#)) OR
 					(reg_q819 AND symb_decoder(16#01#)) OR
 					(reg_q819 AND symb_decoder(16#cf#)) OR
 					(reg_q819 AND symb_decoder(16#a4#)) OR
 					(reg_q819 AND symb_decoder(16#8b#)) OR
 					(reg_q819 AND symb_decoder(16#3f#)) OR
 					(reg_q819 AND symb_decoder(16#f0#)) OR
 					(reg_q819 AND symb_decoder(16#9e#)) OR
 					(reg_q819 AND symb_decoder(16#35#)) OR
 					(reg_q819 AND symb_decoder(16#f8#)) OR
 					(reg_q819 AND symb_decoder(16#a2#)) OR
 					(reg_q819 AND symb_decoder(16#aa#)) OR
 					(reg_q819 AND symb_decoder(16#e5#)) OR
 					(reg_q819 AND symb_decoder(16#bf#)) OR
 					(reg_q819 AND symb_decoder(16#23#)) OR
 					(reg_q819 AND symb_decoder(16#34#)) OR
 					(reg_q819 AND symb_decoder(16#62#)) OR
 					(reg_q819 AND symb_decoder(16#27#)) OR
 					(reg_q819 AND symb_decoder(16#bd#)) OR
 					(reg_q819 AND symb_decoder(16#a3#)) OR
 					(reg_q819 AND symb_decoder(16#8d#)) OR
 					(reg_q819 AND symb_decoder(16#74#)) OR
 					(reg_q819 AND symb_decoder(16#d7#)) OR
 					(reg_q819 AND symb_decoder(16#32#)) OR
 					(reg_q819 AND symb_decoder(16#03#)) OR
 					(reg_q819 AND symb_decoder(16#d9#)) OR
 					(reg_q819 AND symb_decoder(16#1e#)) OR
 					(reg_q819 AND symb_decoder(16#8f#)) OR
 					(reg_q819 AND symb_decoder(16#94#)) OR
 					(reg_q819 AND symb_decoder(16#d6#)) OR
 					(reg_q819 AND symb_decoder(16#cd#)) OR
 					(reg_q819 AND symb_decoder(16#4d#)) OR
 					(reg_q857 AND symb_decoder(16#56#)) OR
 					(reg_q857 AND symb_decoder(16#ac#)) OR
 					(reg_q857 AND symb_decoder(16#50#)) OR
 					(reg_q857 AND symb_decoder(16#6d#)) OR
 					(reg_q857 AND symb_decoder(16#6f#)) OR
 					(reg_q857 AND symb_decoder(16#d6#)) OR
 					(reg_q857 AND symb_decoder(16#84#)) OR
 					(reg_q857 AND symb_decoder(16#d7#)) OR
 					(reg_q857 AND symb_decoder(16#d1#)) OR
 					(reg_q857 AND symb_decoder(16#69#)) OR
 					(reg_q857 AND symb_decoder(16#89#)) OR
 					(reg_q857 AND symb_decoder(16#c3#)) OR
 					(reg_q857 AND symb_decoder(16#44#)) OR
 					(reg_q857 AND symb_decoder(16#c6#)) OR
 					(reg_q857 AND symb_decoder(16#1e#)) OR
 					(reg_q857 AND symb_decoder(16#59#)) OR
 					(reg_q857 AND symb_decoder(16#ba#)) OR
 					(reg_q857 AND symb_decoder(16#b5#)) OR
 					(reg_q857 AND symb_decoder(16#f8#)) OR
 					(reg_q857 AND symb_decoder(16#31#)) OR
 					(reg_q857 AND symb_decoder(16#0f#)) OR
 					(reg_q857 AND symb_decoder(16#bb#)) OR
 					(reg_q857 AND symb_decoder(16#b8#)) OR
 					(reg_q857 AND symb_decoder(16#1f#)) OR
 					(reg_q857 AND symb_decoder(16#d0#)) OR
 					(reg_q857 AND symb_decoder(16#ab#)) OR
 					(reg_q857 AND symb_decoder(16#20#)) OR
 					(reg_q857 AND symb_decoder(16#1c#)) OR
 					(reg_q857 AND symb_decoder(16#ce#)) OR
 					(reg_q857 AND symb_decoder(16#58#)) OR
 					(reg_q857 AND symb_decoder(16#a5#)) OR
 					(reg_q857 AND symb_decoder(16#49#)) OR
 					(reg_q857 AND symb_decoder(16#23#)) OR
 					(reg_q857 AND symb_decoder(16#9d#)) OR
 					(reg_q857 AND symb_decoder(16#a2#)) OR
 					(reg_q857 AND symb_decoder(16#38#)) OR
 					(reg_q857 AND symb_decoder(16#21#)) OR
 					(reg_q857 AND symb_decoder(16#14#)) OR
 					(reg_q857 AND symb_decoder(16#cb#)) OR
 					(reg_q857 AND symb_decoder(16#b7#)) OR
 					(reg_q857 AND symb_decoder(16#f0#)) OR
 					(reg_q857 AND symb_decoder(16#94#)) OR
 					(reg_q857 AND symb_decoder(16#e1#)) OR
 					(reg_q857 AND symb_decoder(16#66#)) OR
 					(reg_q857 AND symb_decoder(16#52#)) OR
 					(reg_q857 AND symb_decoder(16#a7#)) OR
 					(reg_q857 AND symb_decoder(16#22#)) OR
 					(reg_q857 AND symb_decoder(16#87#)) OR
 					(reg_q857 AND symb_decoder(16#8b#)) OR
 					(reg_q857 AND symb_decoder(16#5a#)) OR
 					(reg_q857 AND symb_decoder(16#16#)) OR
 					(reg_q857 AND symb_decoder(16#ff#)) OR
 					(reg_q857 AND symb_decoder(16#8a#)) OR
 					(reg_q857 AND symb_decoder(16#78#)) OR
 					(reg_q857 AND symb_decoder(16#8f#)) OR
 					(reg_q857 AND symb_decoder(16#b3#)) OR
 					(reg_q857 AND symb_decoder(16#ae#)) OR
 					(reg_q857 AND symb_decoder(16#db#)) OR
 					(reg_q857 AND symb_decoder(16#70#)) OR
 					(reg_q857 AND symb_decoder(16#af#)) OR
 					(reg_q857 AND symb_decoder(16#a8#)) OR
 					(reg_q857 AND symb_decoder(16#47#)) OR
 					(reg_q857 AND symb_decoder(16#26#)) OR
 					(reg_q857 AND symb_decoder(16#e4#)) OR
 					(reg_q857 AND symb_decoder(16#43#)) OR
 					(reg_q857 AND symb_decoder(16#8e#)) OR
 					(reg_q857 AND symb_decoder(16#f5#)) OR
 					(reg_q857 AND symb_decoder(16#30#)) OR
 					(reg_q857 AND symb_decoder(16#fa#)) OR
 					(reg_q857 AND symb_decoder(16#5b#)) OR
 					(reg_q857 AND symb_decoder(16#32#)) OR
 					(reg_q857 AND symb_decoder(16#df#)) OR
 					(reg_q857 AND symb_decoder(16#24#)) OR
 					(reg_q857 AND symb_decoder(16#9b#)) OR
 					(reg_q857 AND symb_decoder(16#08#)) OR
 					(reg_q857 AND symb_decoder(16#06#)) OR
 					(reg_q857 AND symb_decoder(16#a4#)) OR
 					(reg_q857 AND symb_decoder(16#c8#)) OR
 					(reg_q857 AND symb_decoder(16#09#)) OR
 					(reg_q857 AND symb_decoder(16#1b#)) OR
 					(reg_q857 AND symb_decoder(16#05#)) OR
 					(reg_q857 AND symb_decoder(16#0b#)) OR
 					(reg_q857 AND symb_decoder(16#9f#)) OR
 					(reg_q857 AND symb_decoder(16#e5#)) OR
 					(reg_q857 AND symb_decoder(16#02#)) OR
 					(reg_q857 AND symb_decoder(16#51#)) OR
 					(reg_q857 AND symb_decoder(16#2a#)) OR
 					(reg_q857 AND symb_decoder(16#f2#)) OR
 					(reg_q857 AND symb_decoder(16#71#)) OR
 					(reg_q857 AND symb_decoder(16#ee#)) OR
 					(reg_q857 AND symb_decoder(16#93#)) OR
 					(reg_q857 AND symb_decoder(16#da#)) OR
 					(reg_q857 AND symb_decoder(16#63#)) OR
 					(reg_q857 AND symb_decoder(16#64#)) OR
 					(reg_q857 AND symb_decoder(16#b9#)) OR
 					(reg_q857 AND symb_decoder(16#a3#)) OR
 					(reg_q857 AND symb_decoder(16#2f#)) OR
 					(reg_q857 AND symb_decoder(16#42#)) OR
 					(reg_q857 AND symb_decoder(16#4f#)) OR
 					(reg_q857 AND symb_decoder(16#eb#)) OR
 					(reg_q857 AND symb_decoder(16#79#)) OR
 					(reg_q857 AND symb_decoder(16#85#)) OR
 					(reg_q857 AND symb_decoder(16#5f#)) OR
 					(reg_q857 AND symb_decoder(16#f6#)) OR
 					(reg_q857 AND symb_decoder(16#76#)) OR
 					(reg_q857 AND symb_decoder(16#9e#)) OR
 					(reg_q857 AND symb_decoder(16#46#)) OR
 					(reg_q857 AND symb_decoder(16#e8#)) OR
 					(reg_q857 AND symb_decoder(16#e0#)) OR
 					(reg_q857 AND symb_decoder(16#6e#)) OR
 					(reg_q857 AND symb_decoder(16#5e#)) OR
 					(reg_q857 AND symb_decoder(16#d4#)) OR
 					(reg_q857 AND symb_decoder(16#c7#)) OR
 					(reg_q857 AND symb_decoder(16#10#)) OR
 					(reg_q857 AND symb_decoder(16#e3#)) OR
 					(reg_q857 AND symb_decoder(16#f4#)) OR
 					(reg_q857 AND symb_decoder(16#61#)) OR
 					(reg_q857 AND symb_decoder(16#17#)) OR
 					(reg_q857 AND symb_decoder(16#ef#)) OR
 					(reg_q857 AND symb_decoder(16#48#)) OR
 					(reg_q857 AND symb_decoder(16#7e#)) OR
 					(reg_q857 AND symb_decoder(16#3f#)) OR
 					(reg_q857 AND symb_decoder(16#25#)) OR
 					(reg_q857 AND symb_decoder(16#91#)) OR
 					(reg_q857 AND symb_decoder(16#fb#)) OR
 					(reg_q857 AND symb_decoder(16#4a#)) OR
 					(reg_q857 AND symb_decoder(16#3d#)) OR
 					(reg_q857 AND symb_decoder(16#53#)) OR
 					(reg_q857 AND symb_decoder(16#c1#)) OR
 					(reg_q857 AND symb_decoder(16#96#)) OR
 					(reg_q857 AND symb_decoder(16#74#)) OR
 					(reg_q857 AND symb_decoder(16#e9#)) OR
 					(reg_q857 AND symb_decoder(16#a0#)) OR
 					(reg_q857 AND symb_decoder(16#95#)) OR
 					(reg_q857 AND symb_decoder(16#73#)) OR
 					(reg_q857 AND symb_decoder(16#7d#)) OR
 					(reg_q857 AND symb_decoder(16#57#)) OR
 					(reg_q857 AND symb_decoder(16#12#)) OR
 					(reg_q857 AND symb_decoder(16#3a#)) OR
 					(reg_q857 AND symb_decoder(16#3e#)) OR
 					(reg_q857 AND symb_decoder(16#b4#)) OR
 					(reg_q857 AND symb_decoder(16#aa#)) OR
 					(reg_q857 AND symb_decoder(16#98#)) OR
 					(reg_q857 AND symb_decoder(16#40#)) OR
 					(reg_q857 AND symb_decoder(16#de#)) OR
 					(reg_q857 AND symb_decoder(16#13#)) OR
 					(reg_q857 AND symb_decoder(16#cf#)) OR
 					(reg_q857 AND symb_decoder(16#2e#)) OR
 					(reg_q857 AND symb_decoder(16#83#)) OR
 					(reg_q857 AND symb_decoder(16#d3#)) OR
 					(reg_q857 AND symb_decoder(16#82#)) OR
 					(reg_q857 AND symb_decoder(16#7a#)) OR
 					(reg_q857 AND symb_decoder(16#68#)) OR
 					(reg_q857 AND symb_decoder(16#7c#)) OR
 					(reg_q857 AND symb_decoder(16#d2#)) OR
 					(reg_q857 AND symb_decoder(16#e7#)) OR
 					(reg_q857 AND symb_decoder(16#c2#)) OR
 					(reg_q857 AND symb_decoder(16#72#)) OR
 					(reg_q857 AND symb_decoder(16#b0#)) OR
 					(reg_q857 AND symb_decoder(16#15#)) OR
 					(reg_q857 AND symb_decoder(16#a6#)) OR
 					(reg_q857 AND symb_decoder(16#54#)) OR
 					(reg_q857 AND symb_decoder(16#7b#)) OR
 					(reg_q857 AND symb_decoder(16#d5#)) OR
 					(reg_q857 AND symb_decoder(16#cc#)) OR
 					(reg_q857 AND symb_decoder(16#ea#)) OR
 					(reg_q857 AND symb_decoder(16#99#)) OR
 					(reg_q857 AND symb_decoder(16#bf#)) OR
 					(reg_q857 AND symb_decoder(16#65#)) OR
 					(reg_q857 AND symb_decoder(16#dc#)) OR
 					(reg_q857 AND symb_decoder(16#90#)) OR
 					(reg_q857 AND symb_decoder(16#62#)) OR
 					(reg_q857 AND symb_decoder(16#a1#)) OR
 					(reg_q857 AND symb_decoder(16#80#)) OR
 					(reg_q857 AND symb_decoder(16#0c#)) OR
 					(reg_q857 AND symb_decoder(16#36#)) OR
 					(reg_q857 AND symb_decoder(16#8c#)) OR
 					(reg_q857 AND symb_decoder(16#88#)) OR
 					(reg_q857 AND symb_decoder(16#39#)) OR
 					(reg_q857 AND symb_decoder(16#b6#)) OR
 					(reg_q857 AND symb_decoder(16#f3#)) OR
 					(reg_q857 AND symb_decoder(16#2d#)) OR
 					(reg_q857 AND symb_decoder(16#f7#)) OR
 					(reg_q857 AND symb_decoder(16#86#)) OR
 					(reg_q857 AND symb_decoder(16#d9#)) OR
 					(reg_q857 AND symb_decoder(16#04#)) OR
 					(reg_q857 AND symb_decoder(16#6b#)) OR
 					(reg_q857 AND symb_decoder(16#c9#)) OR
 					(reg_q857 AND symb_decoder(16#fd#)) OR
 					(reg_q857 AND symb_decoder(16#cd#)) OR
 					(reg_q857 AND symb_decoder(16#18#)) OR
 					(reg_q857 AND symb_decoder(16#37#)) OR
 					(reg_q857 AND symb_decoder(16#4e#)) OR
 					(reg_q857 AND symb_decoder(16#2c#)) OR
 					(reg_q857 AND symb_decoder(16#41#)) OR
 					(reg_q857 AND symb_decoder(16#6a#)) OR
 					(reg_q857 AND symb_decoder(16#d8#)) OR
 					(reg_q857 AND symb_decoder(16#c0#)) OR
 					(reg_q857 AND symb_decoder(16#45#)) OR
 					(reg_q857 AND symb_decoder(16#4b#)) OR
 					(reg_q857 AND symb_decoder(16#dd#)) OR
 					(reg_q857 AND symb_decoder(16#0e#)) OR
 					(reg_q857 AND symb_decoder(16#fc#)) OR
 					(reg_q857 AND symb_decoder(16#34#)) OR
 					(reg_q857 AND symb_decoder(16#4d#)) OR
 					(reg_q857 AND symb_decoder(16#60#)) OR
 					(reg_q857 AND symb_decoder(16#29#)) OR
 					(reg_q857 AND symb_decoder(16#07#)) OR
 					(reg_q857 AND symb_decoder(16#e6#)) OR
 					(reg_q857 AND symb_decoder(16#a9#)) OR
 					(reg_q857 AND symb_decoder(16#f1#)) OR
 					(reg_q857 AND symb_decoder(16#3b#)) OR
 					(reg_q857 AND symb_decoder(16#fe#)) OR
 					(reg_q857 AND symb_decoder(16#3c#)) OR
 					(reg_q857 AND symb_decoder(16#be#)) OR
 					(reg_q857 AND symb_decoder(16#55#)) OR
 					(reg_q857 AND symb_decoder(16#ec#)) OR
 					(reg_q857 AND symb_decoder(16#27#)) OR
 					(reg_q857 AND symb_decoder(16#ed#)) OR
 					(reg_q857 AND symb_decoder(16#03#)) OR
 					(reg_q857 AND symb_decoder(16#33#)) OR
 					(reg_q857 AND symb_decoder(16#ad#)) OR
 					(reg_q857 AND symb_decoder(16#1a#)) OR
 					(reg_q857 AND symb_decoder(16#1d#)) OR
 					(reg_q857 AND symb_decoder(16#97#)) OR
 					(reg_q857 AND symb_decoder(16#2b#)) OR
 					(reg_q857 AND symb_decoder(16#c4#)) OR
 					(reg_q857 AND symb_decoder(16#8d#)) OR
 					(reg_q857 AND symb_decoder(16#81#)) OR
 					(reg_q857 AND symb_decoder(16#7f#)) OR
 					(reg_q857 AND symb_decoder(16#ca#)) OR
 					(reg_q857 AND symb_decoder(16#4c#)) OR
 					(reg_q857 AND symb_decoder(16#c5#)) OR
 					(reg_q857 AND symb_decoder(16#f9#)) OR
 					(reg_q857 AND symb_decoder(16#9c#)) OR
 					(reg_q857 AND symb_decoder(16#b2#)) OR
 					(reg_q857 AND symb_decoder(16#00#)) OR
 					(reg_q857 AND symb_decoder(16#9a#)) OR
 					(reg_q857 AND symb_decoder(16#11#)) OR
 					(reg_q857 AND symb_decoder(16#75#)) OR
 					(reg_q857 AND symb_decoder(16#67#)) OR
 					(reg_q857 AND symb_decoder(16#19#)) OR
 					(reg_q857 AND symb_decoder(16#5d#)) OR
 					(reg_q857 AND symb_decoder(16#b1#)) OR
 					(reg_q857 AND symb_decoder(16#6c#)) OR
 					(reg_q857 AND symb_decoder(16#5c#)) OR
 					(reg_q857 AND symb_decoder(16#bd#)) OR
 					(reg_q857 AND symb_decoder(16#77#)) OR
 					(reg_q857 AND symb_decoder(16#01#)) OR
 					(reg_q857 AND symb_decoder(16#e2#)) OR
 					(reg_q857 AND symb_decoder(16#92#)) OR
 					(reg_q857 AND symb_decoder(16#bc#)) OR
 					(reg_q857 AND symb_decoder(16#35#)) OR
 					(reg_q857 AND symb_decoder(16#28#));
reg_q2629_in <= (reg_q2627 AND symb_decoder(16#dd#)) OR
 					(reg_q2627 AND symb_decoder(16#b6#)) OR
 					(reg_q2627 AND symb_decoder(16#b4#)) OR
 					(reg_q2627 AND symb_decoder(16#2f#)) OR
 					(reg_q2627 AND symb_decoder(16#03#)) OR
 					(reg_q2627 AND symb_decoder(16#00#)) OR
 					(reg_q2627 AND symb_decoder(16#2c#)) OR
 					(reg_q2627 AND symb_decoder(16#d3#)) OR
 					(reg_q2627 AND symb_decoder(16#8f#)) OR
 					(reg_q2627 AND symb_decoder(16#f1#)) OR
 					(reg_q2627 AND symb_decoder(16#2e#)) OR
 					(reg_q2627 AND symb_decoder(16#65#)) OR
 					(reg_q2627 AND symb_decoder(16#02#)) OR
 					(reg_q2627 AND symb_decoder(16#07#)) OR
 					(reg_q2627 AND symb_decoder(16#be#)) OR
 					(reg_q2627 AND symb_decoder(16#fe#)) OR
 					(reg_q2627 AND symb_decoder(16#ef#)) OR
 					(reg_q2627 AND symb_decoder(16#0e#)) OR
 					(reg_q2627 AND symb_decoder(16#ea#)) OR
 					(reg_q2627 AND symb_decoder(16#cc#)) OR
 					(reg_q2627 AND symb_decoder(16#9a#)) OR
 					(reg_q2627 AND symb_decoder(16#ca#)) OR
 					(reg_q2627 AND symb_decoder(16#86#)) OR
 					(reg_q2627 AND symb_decoder(16#fc#)) OR
 					(reg_q2627 AND symb_decoder(16#5b#)) OR
 					(reg_q2627 AND symb_decoder(16#5a#)) OR
 					(reg_q2627 AND symb_decoder(16#37#)) OR
 					(reg_q2627 AND symb_decoder(16#44#)) OR
 					(reg_q2627 AND symb_decoder(16#c3#)) OR
 					(reg_q2627 AND symb_decoder(16#92#)) OR
 					(reg_q2627 AND symb_decoder(16#72#)) OR
 					(reg_q2627 AND symb_decoder(16#e6#)) OR
 					(reg_q2627 AND symb_decoder(16#f8#)) OR
 					(reg_q2627 AND symb_decoder(16#f0#)) OR
 					(reg_q2627 AND symb_decoder(16#a6#)) OR
 					(reg_q2627 AND symb_decoder(16#25#)) OR
 					(reg_q2627 AND symb_decoder(16#b7#)) OR
 					(reg_q2627 AND symb_decoder(16#78#)) OR
 					(reg_q2627 AND symb_decoder(16#2a#)) OR
 					(reg_q2627 AND symb_decoder(16#5f#)) OR
 					(reg_q2627 AND symb_decoder(16#c7#)) OR
 					(reg_q2627 AND symb_decoder(16#50#)) OR
 					(reg_q2627 AND symb_decoder(16#9f#)) OR
 					(reg_q2627 AND symb_decoder(16#1e#)) OR
 					(reg_q2627 AND symb_decoder(16#08#)) OR
 					(reg_q2627 AND symb_decoder(16#a4#)) OR
 					(reg_q2627 AND symb_decoder(16#a8#)) OR
 					(reg_q2627 AND symb_decoder(16#b0#)) OR
 					(reg_q2627 AND symb_decoder(16#a2#)) OR
 					(reg_q2627 AND symb_decoder(16#d4#)) OR
 					(reg_q2627 AND symb_decoder(16#96#)) OR
 					(reg_q2627 AND symb_decoder(16#7b#)) OR
 					(reg_q2627 AND symb_decoder(16#cd#)) OR
 					(reg_q2627 AND symb_decoder(16#39#)) OR
 					(reg_q2627 AND symb_decoder(16#f4#)) OR
 					(reg_q2627 AND symb_decoder(16#34#)) OR
 					(reg_q2627 AND symb_decoder(16#ae#)) OR
 					(reg_q2627 AND symb_decoder(16#a5#)) OR
 					(reg_q2627 AND symb_decoder(16#4d#)) OR
 					(reg_q2627 AND symb_decoder(16#e0#)) OR
 					(reg_q2627 AND symb_decoder(16#fb#)) OR
 					(reg_q2627 AND symb_decoder(16#85#)) OR
 					(reg_q2627 AND symb_decoder(16#51#)) OR
 					(reg_q2627 AND symb_decoder(16#67#)) OR
 					(reg_q2627 AND symb_decoder(16#33#)) OR
 					(reg_q2627 AND symb_decoder(16#52#)) OR
 					(reg_q2627 AND symb_decoder(16#a1#)) OR
 					(reg_q2627 AND symb_decoder(16#e3#)) OR
 					(reg_q2627 AND symb_decoder(16#24#)) OR
 					(reg_q2627 AND symb_decoder(16#90#)) OR
 					(reg_q2627 AND symb_decoder(16#32#)) OR
 					(reg_q2627 AND symb_decoder(16#30#)) OR
 					(reg_q2627 AND symb_decoder(16#b2#)) OR
 					(reg_q2627 AND symb_decoder(16#13#)) OR
 					(reg_q2627 AND symb_decoder(16#99#)) OR
 					(reg_q2627 AND symb_decoder(16#19#)) OR
 					(reg_q2627 AND symb_decoder(16#22#)) OR
 					(reg_q2627 AND symb_decoder(16#71#)) OR
 					(reg_q2627 AND symb_decoder(16#26#)) OR
 					(reg_q2627 AND symb_decoder(16#ee#)) OR
 					(reg_q2627 AND symb_decoder(16#4f#)) OR
 					(reg_q2627 AND symb_decoder(16#9e#)) OR
 					(reg_q2627 AND symb_decoder(16#66#)) OR
 					(reg_q2627 AND symb_decoder(16#b8#)) OR
 					(reg_q2627 AND symb_decoder(16#b5#)) OR
 					(reg_q2627 AND symb_decoder(16#2b#)) OR
 					(reg_q2627 AND symb_decoder(16#81#)) OR
 					(reg_q2627 AND symb_decoder(16#09#)) OR
 					(reg_q2627 AND symb_decoder(16#2d#)) OR
 					(reg_q2627 AND symb_decoder(16#fa#)) OR
 					(reg_q2627 AND symb_decoder(16#0c#)) OR
 					(reg_q2627 AND symb_decoder(16#70#)) OR
 					(reg_q2627 AND symb_decoder(16#6f#)) OR
 					(reg_q2627 AND symb_decoder(16#d8#)) OR
 					(reg_q2627 AND symb_decoder(16#e8#)) OR
 					(reg_q2627 AND symb_decoder(16#c1#)) OR
 					(reg_q2627 AND symb_decoder(16#7a#)) OR
 					(reg_q2627 AND symb_decoder(16#63#)) OR
 					(reg_q2627 AND symb_decoder(16#98#)) OR
 					(reg_q2627 AND symb_decoder(16#68#)) OR
 					(reg_q2627 AND symb_decoder(16#d5#)) OR
 					(reg_q2627 AND symb_decoder(16#40#)) OR
 					(reg_q2627 AND symb_decoder(16#80#)) OR
 					(reg_q2627 AND symb_decoder(16#11#)) OR
 					(reg_q2627 AND symb_decoder(16#ac#)) OR
 					(reg_q2627 AND symb_decoder(16#dc#)) OR
 					(reg_q2627 AND symb_decoder(16#05#)) OR
 					(reg_q2627 AND symb_decoder(16#4a#)) OR
 					(reg_q2627 AND symb_decoder(16#3e#)) OR
 					(reg_q2627 AND symb_decoder(16#c9#)) OR
 					(reg_q2627 AND symb_decoder(16#9c#)) OR
 					(reg_q2627 AND symb_decoder(16#e7#)) OR
 					(reg_q2627 AND symb_decoder(16#69#)) OR
 					(reg_q2627 AND symb_decoder(16#12#)) OR
 					(reg_q2627 AND symb_decoder(16#5d#)) OR
 					(reg_q2627 AND symb_decoder(16#75#)) OR
 					(reg_q2627 AND symb_decoder(16#0f#)) OR
 					(reg_q2627 AND symb_decoder(16#7e#)) OR
 					(reg_q2627 AND symb_decoder(16#7f#)) OR
 					(reg_q2627 AND symb_decoder(16#e1#)) OR
 					(reg_q2627 AND symb_decoder(16#f7#)) OR
 					(reg_q2627 AND symb_decoder(16#89#)) OR
 					(reg_q2627 AND symb_decoder(16#35#)) OR
 					(reg_q2627 AND symb_decoder(16#b9#)) OR
 					(reg_q2627 AND symb_decoder(16#36#)) OR
 					(reg_q2627 AND symb_decoder(16#17#)) OR
 					(reg_q2627 AND symb_decoder(16#cb#)) OR
 					(reg_q2627 AND symb_decoder(16#ad#)) OR
 					(reg_q2627 AND symb_decoder(16#8d#)) OR
 					(reg_q2627 AND symb_decoder(16#aa#)) OR
 					(reg_q2627 AND symb_decoder(16#27#)) OR
 					(reg_q2627 AND symb_decoder(16#45#)) OR
 					(reg_q2627 AND symb_decoder(16#fd#)) OR
 					(reg_q2627 AND symb_decoder(16#d9#)) OR
 					(reg_q2627 AND symb_decoder(16#eb#)) OR
 					(reg_q2627 AND symb_decoder(16#0a#)) OR
 					(reg_q2627 AND symb_decoder(16#8e#)) OR
 					(reg_q2627 AND symb_decoder(16#c0#)) OR
 					(reg_q2627 AND symb_decoder(16#91#)) OR
 					(reg_q2627 AND symb_decoder(16#77#)) OR
 					(reg_q2627 AND symb_decoder(16#c2#)) OR
 					(reg_q2627 AND symb_decoder(16#20#)) OR
 					(reg_q2627 AND symb_decoder(16#31#)) OR
 					(reg_q2627 AND symb_decoder(16#4e#)) OR
 					(reg_q2627 AND symb_decoder(16#9b#)) OR
 					(reg_q2627 AND symb_decoder(16#79#)) OR
 					(reg_q2627 AND symb_decoder(16#8a#)) OR
 					(reg_q2627 AND symb_decoder(16#db#)) OR
 					(reg_q2627 AND symb_decoder(16#42#)) OR
 					(reg_q2627 AND symb_decoder(16#da#)) OR
 					(reg_q2627 AND symb_decoder(16#3f#)) OR
 					(reg_q2627 AND symb_decoder(16#9d#)) OR
 					(reg_q2627 AND symb_decoder(16#6b#)) OR
 					(reg_q2627 AND symb_decoder(16#d7#)) OR
 					(reg_q2627 AND symb_decoder(16#5c#)) OR
 					(reg_q2627 AND symb_decoder(16#46#)) OR
 					(reg_q2627 AND symb_decoder(16#1d#)) OR
 					(reg_q2627 AND symb_decoder(16#de#)) OR
 					(reg_q2627 AND symb_decoder(16#84#)) OR
 					(reg_q2627 AND symb_decoder(16#06#)) OR
 					(reg_q2627 AND symb_decoder(16#0d#)) OR
 					(reg_q2627 AND symb_decoder(16#64#)) OR
 					(reg_q2627 AND symb_decoder(16#6a#)) OR
 					(reg_q2627 AND symb_decoder(16#b1#)) OR
 					(reg_q2627 AND symb_decoder(16#48#)) OR
 					(reg_q2627 AND symb_decoder(16#5e#)) OR
 					(reg_q2627 AND symb_decoder(16#8c#)) OR
 					(reg_q2627 AND symb_decoder(16#ed#)) OR
 					(reg_q2627 AND symb_decoder(16#04#)) OR
 					(reg_q2627 AND symb_decoder(16#83#)) OR
 					(reg_q2627 AND symb_decoder(16#bd#)) OR
 					(reg_q2627 AND symb_decoder(16#c5#)) OR
 					(reg_q2627 AND symb_decoder(16#c4#)) OR
 					(reg_q2627 AND symb_decoder(16#47#)) OR
 					(reg_q2627 AND symb_decoder(16#16#)) OR
 					(reg_q2627 AND symb_decoder(16#bc#)) OR
 					(reg_q2627 AND symb_decoder(16#41#)) OR
 					(reg_q2627 AND symb_decoder(16#28#)) OR
 					(reg_q2627 AND symb_decoder(16#3c#)) OR
 					(reg_q2627 AND symb_decoder(16#01#)) OR
 					(reg_q2627 AND symb_decoder(16#1c#)) OR
 					(reg_q2627 AND symb_decoder(16#61#)) OR
 					(reg_q2627 AND symb_decoder(16#d6#)) OR
 					(reg_q2627 AND symb_decoder(16#ba#)) OR
 					(reg_q2627 AND symb_decoder(16#a3#)) OR
 					(reg_q2627 AND symb_decoder(16#bb#)) OR
 					(reg_q2627 AND symb_decoder(16#d0#)) OR
 					(reg_q2627 AND symb_decoder(16#94#)) OR
 					(reg_q2627 AND symb_decoder(16#af#)) OR
 					(reg_q2627 AND symb_decoder(16#4b#)) OR
 					(reg_q2627 AND symb_decoder(16#ab#)) OR
 					(reg_q2627 AND symb_decoder(16#f6#)) OR
 					(reg_q2627 AND symb_decoder(16#74#)) OR
 					(reg_q2627 AND symb_decoder(16#a0#)) OR
 					(reg_q2627 AND symb_decoder(16#4c#)) OR
 					(reg_q2627 AND symb_decoder(16#a9#)) OR
 					(reg_q2627 AND symb_decoder(16#38#)) OR
 					(reg_q2627 AND symb_decoder(16#6e#)) OR
 					(reg_q2627 AND symb_decoder(16#0b#)) OR
 					(reg_q2627 AND symb_decoder(16#df#)) OR
 					(reg_q2627 AND symb_decoder(16#43#)) OR
 					(reg_q2627 AND symb_decoder(16#29#)) OR
 					(reg_q2627 AND symb_decoder(16#7d#)) OR
 					(reg_q2627 AND symb_decoder(16#93#)) OR
 					(reg_q2627 AND symb_decoder(16#87#)) OR
 					(reg_q2627 AND symb_decoder(16#1f#)) OR
 					(reg_q2627 AND symb_decoder(16#7c#)) OR
 					(reg_q2627 AND symb_decoder(16#c6#)) OR
 					(reg_q2627 AND symb_decoder(16#ec#)) OR
 					(reg_q2627 AND symb_decoder(16#60#)) OR
 					(reg_q2627 AND symb_decoder(16#c8#)) OR
 					(reg_q2627 AND symb_decoder(16#10#)) OR
 					(reg_q2627 AND symb_decoder(16#f2#)) OR
 					(reg_q2627 AND symb_decoder(16#f9#)) OR
 					(reg_q2627 AND symb_decoder(16#49#)) OR
 					(reg_q2627 AND symb_decoder(16#62#)) OR
 					(reg_q2627 AND symb_decoder(16#cf#)) OR
 					(reg_q2627 AND symb_decoder(16#a7#)) OR
 					(reg_q2627 AND symb_decoder(16#ff#)) OR
 					(reg_q2627 AND symb_decoder(16#f3#)) OR
 					(reg_q2627 AND symb_decoder(16#6c#)) OR
 					(reg_q2627 AND symb_decoder(16#55#)) OR
 					(reg_q2627 AND symb_decoder(16#3a#)) OR
 					(reg_q2627 AND symb_decoder(16#3d#)) OR
 					(reg_q2627 AND symb_decoder(16#f5#)) OR
 					(reg_q2627 AND symb_decoder(16#54#)) OR
 					(reg_q2627 AND symb_decoder(16#14#)) OR
 					(reg_q2627 AND symb_decoder(16#58#)) OR
 					(reg_q2627 AND symb_decoder(16#88#)) OR
 					(reg_q2627 AND symb_decoder(16#d1#)) OR
 					(reg_q2627 AND symb_decoder(16#21#)) OR
 					(reg_q2627 AND symb_decoder(16#59#)) OR
 					(reg_q2627 AND symb_decoder(16#3b#)) OR
 					(reg_q2627 AND symb_decoder(16#8b#)) OR
 					(reg_q2627 AND symb_decoder(16#73#)) OR
 					(reg_q2627 AND symb_decoder(16#e2#)) OR
 					(reg_q2627 AND symb_decoder(16#76#)) OR
 					(reg_q2627 AND symb_decoder(16#e9#)) OR
 					(reg_q2627 AND symb_decoder(16#6d#)) OR
 					(reg_q2627 AND symb_decoder(16#23#)) OR
 					(reg_q2627 AND symb_decoder(16#82#)) OR
 					(reg_q2627 AND symb_decoder(16#b3#)) OR
 					(reg_q2627 AND symb_decoder(16#1a#)) OR
 					(reg_q2627 AND symb_decoder(16#53#)) OR
 					(reg_q2627 AND symb_decoder(16#bf#)) OR
 					(reg_q2627 AND symb_decoder(16#e5#)) OR
 					(reg_q2627 AND symb_decoder(16#e4#)) OR
 					(reg_q2627 AND symb_decoder(16#57#)) OR
 					(reg_q2627 AND symb_decoder(16#ce#)) OR
 					(reg_q2627 AND symb_decoder(16#95#)) OR
 					(reg_q2627 AND symb_decoder(16#15#)) OR
 					(reg_q2627 AND symb_decoder(16#56#)) OR
 					(reg_q2627 AND symb_decoder(16#d2#)) OR
 					(reg_q2627 AND symb_decoder(16#18#)) OR
 					(reg_q2627 AND symb_decoder(16#97#)) OR
 					(reg_q2627 AND symb_decoder(16#1b#));
reg_q569_in <= (reg_q565 AND symb_decoder(16#23#)) OR
 					(reg_q587 AND symb_decoder(16#23#));
reg_q571_in <= (reg_q569 AND symb_decoder(16#36#)) OR
 					(reg_q569 AND symb_decoder(16#33#)) OR
 					(reg_q569 AND symb_decoder(16#38#)) OR
 					(reg_q569 AND symb_decoder(16#34#)) OR
 					(reg_q569 AND symb_decoder(16#35#)) OR
 					(reg_q569 AND symb_decoder(16#30#)) OR
 					(reg_q569 AND symb_decoder(16#39#)) OR
 					(reg_q569 AND symb_decoder(16#31#)) OR
 					(reg_q569 AND symb_decoder(16#32#)) OR
 					(reg_q569 AND symb_decoder(16#37#)) OR
 					(reg_q571 AND symb_decoder(16#39#)) OR
 					(reg_q571 AND symb_decoder(16#34#)) OR
 					(reg_q571 AND symb_decoder(16#35#)) OR
 					(reg_q571 AND symb_decoder(16#38#)) OR
 					(reg_q571 AND symb_decoder(16#31#)) OR
 					(reg_q571 AND symb_decoder(16#32#)) OR
 					(reg_q571 AND symb_decoder(16#33#)) OR
 					(reg_q571 AND symb_decoder(16#37#)) OR
 					(reg_q571 AND symb_decoder(16#36#)) OR
 					(reg_q571 AND symb_decoder(16#30#));
reg_q696_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q695 AND symb_decoder(16#73#)) OR
 					(reg_q695 AND symb_decoder(16#53#));
reg_q177_in <= (reg_q185 AND symb_decoder(16#52#)) OR
 					(reg_q185 AND symb_decoder(16#72#)) OR
 					(reg_q173 AND symb_decoder(16#52#)) OR
 					(reg_q173 AND symb_decoder(16#72#));
reg_q665_in <= (reg_q663 AND symb_decoder(16#0a#)) OR
 					(reg_q663 AND symb_decoder(16#20#)) OR
 					(reg_q663 AND symb_decoder(16#0c#)) OR
 					(reg_q663 AND symb_decoder(16#0d#)) OR
 					(reg_q663 AND symb_decoder(16#09#));
reg_q948_in <= (reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q946 AND symb_decoder(16#57#));
reg_q135_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q134 AND symb_decoder(16#52#)) OR
 					(reg_q134 AND symb_decoder(16#72#));
reg_fullgraph20_init <= "0000";

reg_fullgraph20_sel <= "00000" & reg_q135_in & reg_q948_in & reg_q665_in & reg_q177_in & reg_q696_in & reg_q571_in & reg_q569_in & reg_q2629_in & reg_q857_in & reg_q542_in & reg_q393_in;

	--coder fullgraph20
with reg_fullgraph20_sel select
reg_fullgraph20_in <=
	"0001" when "0000000000000001",
	"0010" when "0000000000000010",
	"0011" when "0000000000000100",
	"0100" when "0000000000001000",
	"0101" when "0000000000010000",
	"0110" when "0000000000100000",
	"0111" when "0000000001000000",
	"1000" when "0000000010000000",
	"1001" when "0000000100000000",
	"1010" when "0000001000000000",
	"1011" when "0000010000000000",
	"0000" when others;
 --end coder

	p_reg_fullgraph20: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph20 <= reg_fullgraph20_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph20 <= reg_fullgraph20_init;
        else
          reg_fullgraph20 <= reg_fullgraph20_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph20

		reg_q393 <= '1' when reg_fullgraph20 = "0001" else '0'; 
		reg_q542 <= '1' when reg_fullgraph20 = "0010" else '0'; 
		reg_q857 <= '1' when reg_fullgraph20 = "0011" else '0'; 
		reg_q2629 <= '1' when reg_fullgraph20 = "0100" else '0'; 
		reg_q569 <= '1' when reg_fullgraph20 = "0101" else '0'; 
		reg_q571 <= '1' when reg_fullgraph20 = "0110" else '0'; 
		reg_q696 <= '1' when reg_fullgraph20 = "0111" else '0'; 
		reg_q177 <= '1' when reg_fullgraph20 = "1000" else '0'; 
		reg_q665 <= '1' when reg_fullgraph20 = "1001" else '0'; 
		reg_q948 <= '1' when reg_fullgraph20 = "1010" else '0'; 
		reg_q135 <= '1' when reg_fullgraph20 = "1011" else '0'; 
--end decoder 

reg_q2520_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q2520 AND symb_decoder(16#d0#)) OR
 					(reg_q2520 AND symb_decoder(16#46#)) OR
 					(reg_q2520 AND symb_decoder(16#31#)) OR
 					(reg_q2520 AND symb_decoder(16#4d#)) OR
 					(reg_q2520 AND symb_decoder(16#32#)) OR
 					(reg_q2520 AND symb_decoder(16#fb#)) OR
 					(reg_q2520 AND symb_decoder(16#12#)) OR
 					(reg_q2520 AND symb_decoder(16#f5#)) OR
 					(reg_q2520 AND symb_decoder(16#50#)) OR
 					(reg_q2520 AND symb_decoder(16#57#)) OR
 					(reg_q2520 AND symb_decoder(16#c8#)) OR
 					(reg_q2520 AND symb_decoder(16#dc#)) OR
 					(reg_q2520 AND symb_decoder(16#4a#)) OR
 					(reg_q2520 AND symb_decoder(16#b4#)) OR
 					(reg_q2520 AND symb_decoder(16#77#)) OR
 					(reg_q2520 AND symb_decoder(16#2c#)) OR
 					(reg_q2520 AND symb_decoder(16#9b#)) OR
 					(reg_q2520 AND symb_decoder(16#a9#)) OR
 					(reg_q2520 AND symb_decoder(16#20#)) OR
 					(reg_q2520 AND symb_decoder(16#a7#)) OR
 					(reg_q2520 AND symb_decoder(16#0a#)) OR
 					(reg_q2520 AND symb_decoder(16#69#)) OR
 					(reg_q2520 AND symb_decoder(16#55#)) OR
 					(reg_q2520 AND symb_decoder(16#c2#)) OR
 					(reg_q2520 AND symb_decoder(16#f7#)) OR
 					(reg_q2520 AND symb_decoder(16#05#)) OR
 					(reg_q2520 AND symb_decoder(16#fe#)) OR
 					(reg_q2520 AND symb_decoder(16#a3#)) OR
 					(reg_q2520 AND symb_decoder(16#40#)) OR
 					(reg_q2520 AND symb_decoder(16#19#)) OR
 					(reg_q2520 AND symb_decoder(16#70#)) OR
 					(reg_q2520 AND symb_decoder(16#8f#)) OR
 					(reg_q2520 AND symb_decoder(16#67#)) OR
 					(reg_q2520 AND symb_decoder(16#96#)) OR
 					(reg_q2520 AND symb_decoder(16#d9#)) OR
 					(reg_q2520 AND symb_decoder(16#3a#)) OR
 					(reg_q2520 AND symb_decoder(16#aa#)) OR
 					(reg_q2520 AND symb_decoder(16#bb#)) OR
 					(reg_q2520 AND symb_decoder(16#81#)) OR
 					(reg_q2520 AND symb_decoder(16#e5#)) OR
 					(reg_q2520 AND symb_decoder(16#fc#)) OR
 					(reg_q2520 AND symb_decoder(16#17#)) OR
 					(reg_q2520 AND symb_decoder(16#ce#)) OR
 					(reg_q2520 AND symb_decoder(16#fa#)) OR
 					(reg_q2520 AND symb_decoder(16#25#)) OR
 					(reg_q2520 AND symb_decoder(16#d3#)) OR
 					(reg_q2520 AND symb_decoder(16#de#)) OR
 					(reg_q2520 AND symb_decoder(16#ff#)) OR
 					(reg_q2520 AND symb_decoder(16#4e#)) OR
 					(reg_q2520 AND symb_decoder(16#18#)) OR
 					(reg_q2520 AND symb_decoder(16#c4#)) OR
 					(reg_q2520 AND symb_decoder(16#59#)) OR
 					(reg_q2520 AND symb_decoder(16#0f#)) OR
 					(reg_q2520 AND symb_decoder(16#36#)) OR
 					(reg_q2520 AND symb_decoder(16#91#)) OR
 					(reg_q2520 AND symb_decoder(16#85#)) OR
 					(reg_q2520 AND symb_decoder(16#be#)) OR
 					(reg_q2520 AND symb_decoder(16#0e#)) OR
 					(reg_q2520 AND symb_decoder(16#71#)) OR
 					(reg_q2520 AND symb_decoder(16#ca#)) OR
 					(reg_q2520 AND symb_decoder(16#2b#)) OR
 					(reg_q2520 AND symb_decoder(16#79#)) OR
 					(reg_q2520 AND symb_decoder(16#f3#)) OR
 					(reg_q2520 AND symb_decoder(16#6e#)) OR
 					(reg_q2520 AND symb_decoder(16#90#)) OR
 					(reg_q2520 AND symb_decoder(16#ec#)) OR
 					(reg_q2520 AND symb_decoder(16#bc#)) OR
 					(reg_q2520 AND symb_decoder(16#2e#)) OR
 					(reg_q2520 AND symb_decoder(16#83#)) OR
 					(reg_q2520 AND symb_decoder(16#bd#)) OR
 					(reg_q2520 AND symb_decoder(16#dd#)) OR
 					(reg_q2520 AND symb_decoder(16#d6#)) OR
 					(reg_q2520 AND symb_decoder(16#8b#)) OR
 					(reg_q2520 AND symb_decoder(16#5b#)) OR
 					(reg_q2520 AND symb_decoder(16#c3#)) OR
 					(reg_q2520 AND symb_decoder(16#1f#)) OR
 					(reg_q2520 AND symb_decoder(16#41#)) OR
 					(reg_q2520 AND symb_decoder(16#6a#)) OR
 					(reg_q2520 AND symb_decoder(16#13#)) OR
 					(reg_q2520 AND symb_decoder(16#8e#)) OR
 					(reg_q2520 AND symb_decoder(16#39#)) OR
 					(reg_q2520 AND symb_decoder(16#0d#)) OR
 					(reg_q2520 AND symb_decoder(16#f6#)) OR
 					(reg_q2520 AND symb_decoder(16#8d#)) OR
 					(reg_q2520 AND symb_decoder(16#ae#)) OR
 					(reg_q2520 AND symb_decoder(16#94#)) OR
 					(reg_q2520 AND symb_decoder(16#49#)) OR
 					(reg_q2520 AND symb_decoder(16#56#)) OR
 					(reg_q2520 AND symb_decoder(16#78#)) OR
 					(reg_q2520 AND symb_decoder(16#2f#)) OR
 					(reg_q2520 AND symb_decoder(16#42#)) OR
 					(reg_q2520 AND symb_decoder(16#0c#)) OR
 					(reg_q2520 AND symb_decoder(16#b2#)) OR
 					(reg_q2520 AND symb_decoder(16#df#)) OR
 					(reg_q2520 AND symb_decoder(16#35#)) OR
 					(reg_q2520 AND symb_decoder(16#c9#)) OR
 					(reg_q2520 AND symb_decoder(16#f1#)) OR
 					(reg_q2520 AND symb_decoder(16#6c#)) OR
 					(reg_q2520 AND symb_decoder(16#30#)) OR
 					(reg_q2520 AND symb_decoder(16#58#)) OR
 					(reg_q2520 AND symb_decoder(16#b7#)) OR
 					(reg_q2520 AND symb_decoder(16#97#)) OR
 					(reg_q2520 AND symb_decoder(16#48#)) OR
 					(reg_q2520 AND symb_decoder(16#60#)) OR
 					(reg_q2520 AND symb_decoder(16#68#)) OR
 					(reg_q2520 AND symb_decoder(16#72#)) OR
 					(reg_q2520 AND symb_decoder(16#22#)) OR
 					(reg_q2520 AND symb_decoder(16#9c#)) OR
 					(reg_q2520 AND symb_decoder(16#73#)) OR
 					(reg_q2520 AND symb_decoder(16#e4#)) OR
 					(reg_q2520 AND symb_decoder(16#b9#)) OR
 					(reg_q2520 AND symb_decoder(16#c7#)) OR
 					(reg_q2520 AND symb_decoder(16#a4#)) OR
 					(reg_q2520 AND symb_decoder(16#c1#)) OR
 					(reg_q2520 AND symb_decoder(16#15#)) OR
 					(reg_q2520 AND symb_decoder(16#01#)) OR
 					(reg_q2520 AND symb_decoder(16#b1#)) OR
 					(reg_q2520 AND symb_decoder(16#86#)) OR
 					(reg_q2520 AND symb_decoder(16#9d#)) OR
 					(reg_q2520 AND symb_decoder(16#16#)) OR
 					(reg_q2520 AND symb_decoder(16#44#)) OR
 					(reg_q2520 AND symb_decoder(16#d5#)) OR
 					(reg_q2520 AND symb_decoder(16#fd#)) OR
 					(reg_q2520 AND symb_decoder(16#cb#)) OR
 					(reg_q2520 AND symb_decoder(16#09#)) OR
 					(reg_q2520 AND symb_decoder(16#cd#)) OR
 					(reg_q2520 AND symb_decoder(16#1c#)) OR
 					(reg_q2520 AND symb_decoder(16#65#)) OR
 					(reg_q2520 AND symb_decoder(16#4c#)) OR
 					(reg_q2520 AND symb_decoder(16#63#)) OR
 					(reg_q2520 AND symb_decoder(16#5d#)) OR
 					(reg_q2520 AND symb_decoder(16#64#)) OR
 					(reg_q2520 AND symb_decoder(16#e2#)) OR
 					(reg_q2520 AND symb_decoder(16#14#)) OR
 					(reg_q2520 AND symb_decoder(16#29#)) OR
 					(reg_q2520 AND symb_decoder(16#95#)) OR
 					(reg_q2520 AND symb_decoder(16#75#)) OR
 					(reg_q2520 AND symb_decoder(16#37#)) OR
 					(reg_q2520 AND symb_decoder(16#6f#)) OR
 					(reg_q2520 AND symb_decoder(16#61#)) OR
 					(reg_q2520 AND symb_decoder(16#11#)) OR
 					(reg_q2520 AND symb_decoder(16#4f#)) OR
 					(reg_q2520 AND symb_decoder(16#10#)) OR
 					(reg_q2520 AND symb_decoder(16#3c#)) OR
 					(reg_q2520 AND symb_decoder(16#e1#)) OR
 					(reg_q2520 AND symb_decoder(16#33#)) OR
 					(reg_q2520 AND symb_decoder(16#07#)) OR
 					(reg_q2520 AND symb_decoder(16#e0#)) OR
 					(reg_q2520 AND symb_decoder(16#c0#)) OR
 					(reg_q2520 AND symb_decoder(16#00#)) OR
 					(reg_q2520 AND symb_decoder(16#9f#)) OR
 					(reg_q2520 AND symb_decoder(16#02#)) OR
 					(reg_q2520 AND symb_decoder(16#e3#)) OR
 					(reg_q2520 AND symb_decoder(16#98#)) OR
 					(reg_q2520 AND symb_decoder(16#7c#)) OR
 					(reg_q2520 AND symb_decoder(16#f9#)) OR
 					(reg_q2520 AND symb_decoder(16#a1#)) OR
 					(reg_q2520 AND symb_decoder(16#52#)) OR
 					(reg_q2520 AND symb_decoder(16#28#)) OR
 					(reg_q2520 AND symb_decoder(16#6b#)) OR
 					(reg_q2520 AND symb_decoder(16#04#)) OR
 					(reg_q2520 AND symb_decoder(16#ac#)) OR
 					(reg_q2520 AND symb_decoder(16#da#)) OR
 					(reg_q2520 AND symb_decoder(16#38#)) OR
 					(reg_q2520 AND symb_decoder(16#06#)) OR
 					(reg_q2520 AND symb_decoder(16#5e#)) OR
 					(reg_q2520 AND symb_decoder(16#5a#)) OR
 					(reg_q2520 AND symb_decoder(16#f8#)) OR
 					(reg_q2520 AND symb_decoder(16#66#)) OR
 					(reg_q2520 AND symb_decoder(16#93#)) OR
 					(reg_q2520 AND symb_decoder(16#43#)) OR
 					(reg_q2520 AND symb_decoder(16#1a#)) OR
 					(reg_q2520 AND symb_decoder(16#47#)) OR
 					(reg_q2520 AND symb_decoder(16#34#)) OR
 					(reg_q2520 AND symb_decoder(16#1d#)) OR
 					(reg_q2520 AND symb_decoder(16#a5#)) OR
 					(reg_q2520 AND symb_decoder(16#5f#)) OR
 					(reg_q2520 AND symb_decoder(16#3b#)) OR
 					(reg_q2520 AND symb_decoder(16#c5#)) OR
 					(reg_q2520 AND symb_decoder(16#54#)) OR
 					(reg_q2520 AND symb_decoder(16#e9#)) OR
 					(reg_q2520 AND symb_decoder(16#db#)) OR
 					(reg_q2520 AND symb_decoder(16#ea#)) OR
 					(reg_q2520 AND symb_decoder(16#62#)) OR
 					(reg_q2520 AND symb_decoder(16#24#)) OR
 					(reg_q2520 AND symb_decoder(16#08#)) OR
 					(reg_q2520 AND symb_decoder(16#3f#)) OR
 					(reg_q2520 AND symb_decoder(16#9e#)) OR
 					(reg_q2520 AND symb_decoder(16#80#)) OR
 					(reg_q2520 AND symb_decoder(16#d2#)) OR
 					(reg_q2520 AND symb_decoder(16#45#)) OR
 					(reg_q2520 AND symb_decoder(16#e8#)) OR
 					(reg_q2520 AND symb_decoder(16#d1#)) OR
 					(reg_q2520 AND symb_decoder(16#ba#)) OR
 					(reg_q2520 AND symb_decoder(16#ee#)) OR
 					(reg_q2520 AND symb_decoder(16#7d#)) OR
 					(reg_q2520 AND symb_decoder(16#87#)) OR
 					(reg_q2520 AND symb_decoder(16#89#)) OR
 					(reg_q2520 AND symb_decoder(16#bf#)) OR
 					(reg_q2520 AND symb_decoder(16#af#)) OR
 					(reg_q2520 AND symb_decoder(16#1b#)) OR
 					(reg_q2520 AND symb_decoder(16#ef#)) OR
 					(reg_q2520 AND symb_decoder(16#82#)) OR
 					(reg_q2520 AND symb_decoder(16#8c#)) OR
 					(reg_q2520 AND symb_decoder(16#ab#)) OR
 					(reg_q2520 AND symb_decoder(16#4b#)) OR
 					(reg_q2520 AND symb_decoder(16#6d#)) OR
 					(reg_q2520 AND symb_decoder(16#2d#)) OR
 					(reg_q2520 AND symb_decoder(16#03#)) OR
 					(reg_q2520 AND symb_decoder(16#7f#)) OR
 					(reg_q2520 AND symb_decoder(16#2a#)) OR
 					(reg_q2520 AND symb_decoder(16#ed#)) OR
 					(reg_q2520 AND symb_decoder(16#21#)) OR
 					(reg_q2520 AND symb_decoder(16#cf#)) OR
 					(reg_q2520 AND symb_decoder(16#f0#)) OR
 					(reg_q2520 AND symb_decoder(16#9a#)) OR
 					(reg_q2520 AND symb_decoder(16#27#)) OR
 					(reg_q2520 AND symb_decoder(16#f2#)) OR
 					(reg_q2520 AND symb_decoder(16#a6#)) OR
 					(reg_q2520 AND symb_decoder(16#e7#)) OR
 					(reg_q2520 AND symb_decoder(16#0b#)) OR
 					(reg_q2520 AND symb_decoder(16#d8#)) OR
 					(reg_q2520 AND symb_decoder(16#b6#)) OR
 					(reg_q2520 AND symb_decoder(16#51#)) OR
 					(reg_q2520 AND symb_decoder(16#d4#)) OR
 					(reg_q2520 AND symb_decoder(16#99#)) OR
 					(reg_q2520 AND symb_decoder(16#a8#)) OR
 					(reg_q2520 AND symb_decoder(16#8a#)) OR
 					(reg_q2520 AND symb_decoder(16#b0#)) OR
 					(reg_q2520 AND symb_decoder(16#7a#)) OR
 					(reg_q2520 AND symb_decoder(16#f4#)) OR
 					(reg_q2520 AND symb_decoder(16#5c#)) OR
 					(reg_q2520 AND symb_decoder(16#7e#)) OR
 					(reg_q2520 AND symb_decoder(16#88#)) OR
 					(reg_q2520 AND symb_decoder(16#b3#)) OR
 					(reg_q2520 AND symb_decoder(16#eb#)) OR
 					(reg_q2520 AND symb_decoder(16#26#)) OR
 					(reg_q2520 AND symb_decoder(16#3e#)) OR
 					(reg_q2520 AND symb_decoder(16#1e#)) OR
 					(reg_q2520 AND symb_decoder(16#cc#)) OR
 					(reg_q2520 AND symb_decoder(16#84#)) OR
 					(reg_q2520 AND symb_decoder(16#d7#)) OR
 					(reg_q2520 AND symb_decoder(16#ad#)) OR
 					(reg_q2520 AND symb_decoder(16#53#)) OR
 					(reg_q2520 AND symb_decoder(16#b5#)) OR
 					(reg_q2520 AND symb_decoder(16#a0#)) OR
 					(reg_q2520 AND symb_decoder(16#92#)) OR
 					(reg_q2520 AND symb_decoder(16#e6#)) OR
 					(reg_q2520 AND symb_decoder(16#7b#)) OR
 					(reg_q2520 AND symb_decoder(16#c6#)) OR
 					(reg_q2520 AND symb_decoder(16#a2#)) OR
 					(reg_q2520 AND symb_decoder(16#76#)) OR
 					(reg_q2520 AND symb_decoder(16#74#)) OR
 					(reg_q2520 AND symb_decoder(16#3d#)) OR
 					(reg_q2520 AND symb_decoder(16#23#)) OR
 					(reg_q2520 AND symb_decoder(16#b8#));
reg_q2520_init <= '0' ;
	p_reg_q2520: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2520 <= reg_q2520_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2520 <= reg_q2520_init;
        else
          reg_q2520 <= reg_q2520_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph22

reg_q2447_in <= (reg_q2429 AND symb_decoder(16#e7#)) OR
 					(reg_q2429 AND symb_decoder(16#7e#)) OR
 					(reg_q2429 AND symb_decoder(16#90#)) OR
 					(reg_q2429 AND symb_decoder(16#fa#)) OR
 					(reg_q2429 AND symb_decoder(16#33#)) OR
 					(reg_q2429 AND symb_decoder(16#4e#)) OR
 					(reg_q2429 AND symb_decoder(16#5f#)) OR
 					(reg_q2429 AND symb_decoder(16#9e#)) OR
 					(reg_q2429 AND symb_decoder(16#fd#)) OR
 					(reg_q2429 AND symb_decoder(16#ec#)) OR
 					(reg_q2429 AND symb_decoder(16#9f#)) OR
 					(reg_q2429 AND symb_decoder(16#96#)) OR
 					(reg_q2429 AND symb_decoder(16#40#)) OR
 					(reg_q2429 AND symb_decoder(16#72#)) OR
 					(reg_q2429 AND symb_decoder(16#ed#)) OR
 					(reg_q2429 AND symb_decoder(16#a6#)) OR
 					(reg_q2429 AND symb_decoder(16#34#)) OR
 					(reg_q2429 AND symb_decoder(16#56#)) OR
 					(reg_q2429 AND symb_decoder(16#44#)) OR
 					(reg_q2429 AND symb_decoder(16#a0#)) OR
 					(reg_q2429 AND symb_decoder(16#e6#)) OR
 					(reg_q2429 AND symb_decoder(16#b0#)) OR
 					(reg_q2429 AND symb_decoder(16#85#)) OR
 					(reg_q2429 AND symb_decoder(16#0f#)) OR
 					(reg_q2429 AND symb_decoder(16#06#)) OR
 					(reg_q2429 AND symb_decoder(16#8c#)) OR
 					(reg_q2429 AND symb_decoder(16#1b#)) OR
 					(reg_q2429 AND symb_decoder(16#30#)) OR
 					(reg_q2429 AND symb_decoder(16#93#)) OR
 					(reg_q2429 AND symb_decoder(16#71#)) OR
 					(reg_q2429 AND symb_decoder(16#50#)) OR
 					(reg_q2429 AND symb_decoder(16#79#)) OR
 					(reg_q2429 AND symb_decoder(16#4c#)) OR
 					(reg_q2429 AND symb_decoder(16#25#)) OR
 					(reg_q2429 AND symb_decoder(16#b5#)) OR
 					(reg_q2429 AND symb_decoder(16#bc#)) OR
 					(reg_q2429 AND symb_decoder(16#7c#)) OR
 					(reg_q2429 AND symb_decoder(16#e4#)) OR
 					(reg_q2429 AND symb_decoder(16#43#)) OR
 					(reg_q2429 AND symb_decoder(16#64#)) OR
 					(reg_q2429 AND symb_decoder(16#cd#)) OR
 					(reg_q2429 AND symb_decoder(16#f5#)) OR
 					(reg_q2429 AND symb_decoder(16#1f#)) OR
 					(reg_q2429 AND symb_decoder(16#b1#)) OR
 					(reg_q2429 AND symb_decoder(16#da#)) OR
 					(reg_q2429 AND symb_decoder(16#95#)) OR
 					(reg_q2429 AND symb_decoder(16#a3#)) OR
 					(reg_q2429 AND symb_decoder(16#78#)) OR
 					(reg_q2429 AND symb_decoder(16#66#)) OR
 					(reg_q2429 AND symb_decoder(16#f8#)) OR
 					(reg_q2429 AND symb_decoder(16#38#)) OR
 					(reg_q2429 AND symb_decoder(16#d4#)) OR
 					(reg_q2429 AND symb_decoder(16#af#)) OR
 					(reg_q2429 AND symb_decoder(16#f3#)) OR
 					(reg_q2429 AND symb_decoder(16#97#)) OR
 					(reg_q2429 AND symb_decoder(16#5b#)) OR
 					(reg_q2429 AND symb_decoder(16#5c#)) OR
 					(reg_q2429 AND symb_decoder(16#24#)) OR
 					(reg_q2429 AND symb_decoder(16#1d#)) OR
 					(reg_q2429 AND symb_decoder(16#57#)) OR
 					(reg_q2429 AND symb_decoder(16#2c#)) OR
 					(reg_q2429 AND symb_decoder(16#17#)) OR
 					(reg_q2429 AND symb_decoder(16#2a#)) OR
 					(reg_q2429 AND symb_decoder(16#6d#)) OR
 					(reg_q2429 AND symb_decoder(16#89#)) OR
 					(reg_q2429 AND symb_decoder(16#2e#)) OR
 					(reg_q2429 AND symb_decoder(16#c4#)) OR
 					(reg_q2429 AND symb_decoder(16#dc#)) OR
 					(reg_q2429 AND symb_decoder(16#58#)) OR
 					(reg_q2429 AND symb_decoder(16#37#)) OR
 					(reg_q2429 AND symb_decoder(16#9a#)) OR
 					(reg_q2429 AND symb_decoder(16#04#)) OR
 					(reg_q2429 AND symb_decoder(16#3f#)) OR
 					(reg_q2429 AND symb_decoder(16#7f#)) OR
 					(reg_q2429 AND symb_decoder(16#7d#)) OR
 					(reg_q2429 AND symb_decoder(16#1a#)) OR
 					(reg_q2429 AND symb_decoder(16#6b#)) OR
 					(reg_q2429 AND symb_decoder(16#8a#)) OR
 					(reg_q2429 AND symb_decoder(16#0b#)) OR
 					(reg_q2429 AND symb_decoder(16#be#)) OR
 					(reg_q2429 AND symb_decoder(16#99#)) OR
 					(reg_q2429 AND symb_decoder(16#b9#)) OR
 					(reg_q2429 AND symb_decoder(16#2b#)) OR
 					(reg_q2429 AND symb_decoder(16#11#)) OR
 					(reg_q2429 AND symb_decoder(16#67#)) OR
 					(reg_q2429 AND symb_decoder(16#26#)) OR
 					(reg_q2429 AND symb_decoder(16#f9#)) OR
 					(reg_q2429 AND symb_decoder(16#c5#)) OR
 					(reg_q2429 AND symb_decoder(16#ac#)) OR
 					(reg_q2429 AND symb_decoder(16#9d#)) OR
 					(reg_q2429 AND symb_decoder(16#62#)) OR
 					(reg_q2429 AND symb_decoder(16#29#)) OR
 					(reg_q2429 AND symb_decoder(16#ee#)) OR
 					(reg_q2429 AND symb_decoder(16#7b#)) OR
 					(reg_q2429 AND symb_decoder(16#ae#)) OR
 					(reg_q2429 AND symb_decoder(16#f1#)) OR
 					(reg_q2429 AND symb_decoder(16#e9#)) OR
 					(reg_q2429 AND symb_decoder(16#0c#)) OR
 					(reg_q2429 AND symb_decoder(16#9b#)) OR
 					(reg_q2429 AND symb_decoder(16#09#)) OR
 					(reg_q2429 AND symb_decoder(16#6c#)) OR
 					(reg_q2429 AND symb_decoder(16#32#)) OR
 					(reg_q2429 AND symb_decoder(16#e3#)) OR
 					(reg_q2429 AND symb_decoder(16#54#)) OR
 					(reg_q2429 AND symb_decoder(16#1e#)) OR
 					(reg_q2429 AND symb_decoder(16#74#)) OR
 					(reg_q2429 AND symb_decoder(16#a9#)) OR
 					(reg_q2429 AND symb_decoder(16#69#)) OR
 					(reg_q2429 AND symb_decoder(16#3d#)) OR
 					(reg_q2429 AND symb_decoder(16#16#)) OR
 					(reg_q2429 AND symb_decoder(16#51#)) OR
 					(reg_q2429 AND symb_decoder(16#12#)) OR
 					(reg_q2429 AND symb_decoder(16#b6#)) OR
 					(reg_q2429 AND symb_decoder(16#0e#)) OR
 					(reg_q2429 AND symb_decoder(16#81#)) OR
 					(reg_q2429 AND symb_decoder(16#03#)) OR
 					(reg_q2429 AND symb_decoder(16#27#)) OR
 					(reg_q2429 AND symb_decoder(16#52#)) OR
 					(reg_q2429 AND symb_decoder(16#02#)) OR
 					(reg_q2429 AND symb_decoder(16#83#)) OR
 					(reg_q2429 AND symb_decoder(16#e1#)) OR
 					(reg_q2429 AND symb_decoder(16#c0#)) OR
 					(reg_q2429 AND symb_decoder(16#08#)) OR
 					(reg_q2429 AND symb_decoder(16#4a#)) OR
 					(reg_q2429 AND symb_decoder(16#00#)) OR
 					(reg_q2429 AND symb_decoder(16#cf#)) OR
 					(reg_q2429 AND symb_decoder(16#db#)) OR
 					(reg_q2429 AND symb_decoder(16#46#)) OR
 					(reg_q2429 AND symb_decoder(16#59#)) OR
 					(reg_q2429 AND symb_decoder(16#c1#)) OR
 					(reg_q2429 AND symb_decoder(16#36#)) OR
 					(reg_q2429 AND symb_decoder(16#f0#)) OR
 					(reg_q2429 AND symb_decoder(16#3a#)) OR
 					(reg_q2429 AND symb_decoder(16#d3#)) OR
 					(reg_q2429 AND symb_decoder(16#88#)) OR
 					(reg_q2429 AND symb_decoder(16#77#)) OR
 					(reg_q2429 AND symb_decoder(16#65#)) OR
 					(reg_q2429 AND symb_decoder(16#4d#)) OR
 					(reg_q2429 AND symb_decoder(16#63#)) OR
 					(reg_q2429 AND symb_decoder(16#68#)) OR
 					(reg_q2429 AND symb_decoder(16#82#)) OR
 					(reg_q2429 AND symb_decoder(16#e2#)) OR
 					(reg_q2429 AND symb_decoder(16#fb#)) OR
 					(reg_q2429 AND symb_decoder(16#18#)) OR
 					(reg_q2429 AND symb_decoder(16#d7#)) OR
 					(reg_q2429 AND symb_decoder(16#f4#)) OR
 					(reg_q2429 AND symb_decoder(16#3b#)) OR
 					(reg_q2429 AND symb_decoder(16#ff#)) OR
 					(reg_q2429 AND symb_decoder(16#8e#)) OR
 					(reg_q2429 AND symb_decoder(16#35#)) OR
 					(reg_q2429 AND symb_decoder(16#9c#)) OR
 					(reg_q2429 AND symb_decoder(16#60#)) OR
 					(reg_q2429 AND symb_decoder(16#7a#)) OR
 					(reg_q2429 AND symb_decoder(16#b4#)) OR
 					(reg_q2429 AND symb_decoder(16#5a#)) OR
 					(reg_q2429 AND symb_decoder(16#87#)) OR
 					(reg_q2429 AND symb_decoder(16#55#)) OR
 					(reg_q2429 AND symb_decoder(16#bd#)) OR
 					(reg_q2429 AND symb_decoder(16#01#)) OR
 					(reg_q2429 AND symb_decoder(16#d9#)) OR
 					(reg_q2429 AND symb_decoder(16#d5#)) OR
 					(reg_q2429 AND symb_decoder(16#5e#)) OR
 					(reg_q2429 AND symb_decoder(16#41#)) OR
 					(reg_q2429 AND symb_decoder(16#22#)) OR
 					(reg_q2429 AND symb_decoder(16#19#)) OR
 					(reg_q2429 AND symb_decoder(16#31#)) OR
 					(reg_q2429 AND symb_decoder(16#c7#)) OR
 					(reg_q2429 AND symb_decoder(16#86#)) OR
 					(reg_q2429 AND symb_decoder(16#75#)) OR
 					(reg_q2429 AND symb_decoder(16#e8#)) OR
 					(reg_q2429 AND symb_decoder(16#70#)) OR
 					(reg_q2429 AND symb_decoder(16#d8#)) OR
 					(reg_q2429 AND symb_decoder(16#c2#)) OR
 					(reg_q2429 AND symb_decoder(16#98#)) OR
 					(reg_q2429 AND symb_decoder(16#45#)) OR
 					(reg_q2429 AND symb_decoder(16#2f#)) OR
 					(reg_q2429 AND symb_decoder(16#b3#)) OR
 					(reg_q2429 AND symb_decoder(16#84#)) OR
 					(reg_q2429 AND symb_decoder(16#bb#)) OR
 					(reg_q2429 AND symb_decoder(16#23#)) OR
 					(reg_q2429 AND symb_decoder(16#10#)) OR
 					(reg_q2429 AND symb_decoder(16#8f#)) OR
 					(reg_q2429 AND symb_decoder(16#61#)) OR
 					(reg_q2429 AND symb_decoder(16#42#)) OR
 					(reg_q2429 AND symb_decoder(16#e5#)) OR
 					(reg_q2429 AND symb_decoder(16#05#)) OR
 					(reg_q2429 AND symb_decoder(16#3e#)) OR
 					(reg_q2429 AND symb_decoder(16#bf#)) OR
 					(reg_q2429 AND symb_decoder(16#a1#)) OR
 					(reg_q2429 AND symb_decoder(16#4f#)) OR
 					(reg_q2429 AND symb_decoder(16#eb#)) OR
 					(reg_q2429 AND symb_decoder(16#c9#)) OR
 					(reg_q2429 AND symb_decoder(16#b2#)) OR
 					(reg_q2429 AND symb_decoder(16#14#)) OR
 					(reg_q2429 AND symb_decoder(16#39#)) OR
 					(reg_q2429 AND symb_decoder(16#cb#)) OR
 					(reg_q2429 AND symb_decoder(16#fe#)) OR
 					(reg_q2429 AND symb_decoder(16#94#)) OR
 					(reg_q2429 AND symb_decoder(16#a4#)) OR
 					(reg_q2429 AND symb_decoder(16#d0#)) OR
 					(reg_q2429 AND symb_decoder(16#c8#)) OR
 					(reg_q2429 AND symb_decoder(16#f7#)) OR
 					(reg_q2429 AND symb_decoder(16#73#)) OR
 					(reg_q2429 AND symb_decoder(16#a7#)) OR
 					(reg_q2429 AND symb_decoder(16#48#)) OR
 					(reg_q2429 AND symb_decoder(16#ce#)) OR
 					(reg_q2429 AND symb_decoder(16#ad#)) OR
 					(reg_q2429 AND symb_decoder(16#4b#)) OR
 					(reg_q2429 AND symb_decoder(16#de#)) OR
 					(reg_q2429 AND symb_decoder(16#47#)) OR
 					(reg_q2429 AND symb_decoder(16#dd#)) OR
 					(reg_q2429 AND symb_decoder(16#21#)) OR
 					(reg_q2429 AND symb_decoder(16#6e#)) OR
 					(reg_q2429 AND symb_decoder(16#3c#)) OR
 					(reg_q2429 AND symb_decoder(16#d1#)) OR
 					(reg_q2429 AND symb_decoder(16#d2#)) OR
 					(reg_q2429 AND symb_decoder(16#6f#)) OR
 					(reg_q2429 AND symb_decoder(16#c6#)) OR
 					(reg_q2429 AND symb_decoder(16#b7#)) OR
 					(reg_q2429 AND symb_decoder(16#df#)) OR
 					(reg_q2429 AND symb_decoder(16#f2#)) OR
 					(reg_q2429 AND symb_decoder(16#aa#)) OR
 					(reg_q2429 AND symb_decoder(16#5d#)) OR
 					(reg_q2429 AND symb_decoder(16#6a#)) OR
 					(reg_q2429 AND symb_decoder(16#15#)) OR
 					(reg_q2429 AND symb_decoder(16#ab#)) OR
 					(reg_q2429 AND symb_decoder(16#cc#)) OR
 					(reg_q2429 AND symb_decoder(16#ea#)) OR
 					(reg_q2429 AND symb_decoder(16#c3#)) OR
 					(reg_q2429 AND symb_decoder(16#20#)) OR
 					(reg_q2429 AND symb_decoder(16#07#)) OR
 					(reg_q2429 AND symb_decoder(16#ca#)) OR
 					(reg_q2429 AND symb_decoder(16#8b#)) OR
 					(reg_q2429 AND symb_decoder(16#28#)) OR
 					(reg_q2429 AND symb_decoder(16#a2#)) OR
 					(reg_q2429 AND symb_decoder(16#53#)) OR
 					(reg_q2429 AND symb_decoder(16#fc#)) OR
 					(reg_q2429 AND symb_decoder(16#49#)) OR
 					(reg_q2429 AND symb_decoder(16#a5#)) OR
 					(reg_q2429 AND symb_decoder(16#91#)) OR
 					(reg_q2429 AND symb_decoder(16#ef#)) OR
 					(reg_q2429 AND symb_decoder(16#d6#)) OR
 					(reg_q2429 AND symb_decoder(16#2d#)) OR
 					(reg_q2429 AND symb_decoder(16#1c#)) OR
 					(reg_q2429 AND symb_decoder(16#ba#)) OR
 					(reg_q2429 AND symb_decoder(16#b8#)) OR
 					(reg_q2429 AND symb_decoder(16#a8#)) OR
 					(reg_q2429 AND symb_decoder(16#f6#)) OR
 					(reg_q2429 AND symb_decoder(16#76#)) OR
 					(reg_q2429 AND symb_decoder(16#92#)) OR
 					(reg_q2429 AND symb_decoder(16#e0#)) OR
 					(reg_q2429 AND symb_decoder(16#8d#)) OR
 					(reg_q2429 AND symb_decoder(16#80#)) OR
 					(reg_q2429 AND symb_decoder(16#13#)) OR
 					(reg_q2447 AND symb_decoder(16#d2#)) OR
 					(reg_q2447 AND symb_decoder(16#f7#)) OR
 					(reg_q2447 AND symb_decoder(16#6c#)) OR
 					(reg_q2447 AND symb_decoder(16#89#)) OR
 					(reg_q2447 AND symb_decoder(16#a9#)) OR
 					(reg_q2447 AND symb_decoder(16#85#)) OR
 					(reg_q2447 AND symb_decoder(16#fe#)) OR
 					(reg_q2447 AND symb_decoder(16#82#)) OR
 					(reg_q2447 AND symb_decoder(16#5d#)) OR
 					(reg_q2447 AND symb_decoder(16#d4#)) OR
 					(reg_q2447 AND symb_decoder(16#22#)) OR
 					(reg_q2447 AND symb_decoder(16#e9#)) OR
 					(reg_q2447 AND symb_decoder(16#20#)) OR
 					(reg_q2447 AND symb_decoder(16#2a#)) OR
 					(reg_q2447 AND symb_decoder(16#94#)) OR
 					(reg_q2447 AND symb_decoder(16#e2#)) OR
 					(reg_q2447 AND symb_decoder(16#0e#)) OR
 					(reg_q2447 AND symb_decoder(16#d9#)) OR
 					(reg_q2447 AND symb_decoder(16#db#)) OR
 					(reg_q2447 AND symb_decoder(16#8c#)) OR
 					(reg_q2447 AND symb_decoder(16#06#)) OR
 					(reg_q2447 AND symb_decoder(16#b6#)) OR
 					(reg_q2447 AND symb_decoder(16#96#)) OR
 					(reg_q2447 AND symb_decoder(16#3b#)) OR
 					(reg_q2447 AND symb_decoder(16#f0#)) OR
 					(reg_q2447 AND symb_decoder(16#2e#)) OR
 					(reg_q2447 AND symb_decoder(16#25#)) OR
 					(reg_q2447 AND symb_decoder(16#9e#)) OR
 					(reg_q2447 AND symb_decoder(16#d3#)) OR
 					(reg_q2447 AND symb_decoder(16#ec#)) OR
 					(reg_q2447 AND symb_decoder(16#39#)) OR
 					(reg_q2447 AND symb_decoder(16#6f#)) OR
 					(reg_q2447 AND symb_decoder(16#d8#)) OR
 					(reg_q2447 AND symb_decoder(16#69#)) OR
 					(reg_q2447 AND symb_decoder(16#8e#)) OR
 					(reg_q2447 AND symb_decoder(16#53#)) OR
 					(reg_q2447 AND symb_decoder(16#5b#)) OR
 					(reg_q2447 AND symb_decoder(16#de#)) OR
 					(reg_q2447 AND symb_decoder(16#ed#)) OR
 					(reg_q2447 AND symb_decoder(16#4e#)) OR
 					(reg_q2447 AND symb_decoder(16#c9#)) OR
 					(reg_q2447 AND symb_decoder(16#58#)) OR
 					(reg_q2447 AND symb_decoder(16#b8#)) OR
 					(reg_q2447 AND symb_decoder(16#5f#)) OR
 					(reg_q2447 AND symb_decoder(16#6a#)) OR
 					(reg_q2447 AND symb_decoder(16#24#)) OR
 					(reg_q2447 AND symb_decoder(16#66#)) OR
 					(reg_q2447 AND symb_decoder(16#29#)) OR
 					(reg_q2447 AND symb_decoder(16#72#)) OR
 					(reg_q2447 AND symb_decoder(16#cc#)) OR
 					(reg_q2447 AND symb_decoder(16#e5#)) OR
 					(reg_q2447 AND symb_decoder(16#bb#)) OR
 					(reg_q2447 AND symb_decoder(16#98#)) OR
 					(reg_q2447 AND symb_decoder(16#3c#)) OR
 					(reg_q2447 AND symb_decoder(16#26#)) OR
 					(reg_q2447 AND symb_decoder(16#97#)) OR
 					(reg_q2447 AND symb_decoder(16#3f#)) OR
 					(reg_q2447 AND symb_decoder(16#9d#)) OR
 					(reg_q2447 AND symb_decoder(16#45#)) OR
 					(reg_q2447 AND symb_decoder(16#4a#)) OR
 					(reg_q2447 AND symb_decoder(16#0b#)) OR
 					(reg_q2447 AND symb_decoder(16#51#)) OR
 					(reg_q2447 AND symb_decoder(16#a4#)) OR
 					(reg_q2447 AND symb_decoder(16#5e#)) OR
 					(reg_q2447 AND symb_decoder(16#73#)) OR
 					(reg_q2447 AND symb_decoder(16#23#)) OR
 					(reg_q2447 AND symb_decoder(16#18#)) OR
 					(reg_q2447 AND symb_decoder(16#76#)) OR
 					(reg_q2447 AND symb_decoder(16#ce#)) OR
 					(reg_q2447 AND symb_decoder(16#17#)) OR
 					(reg_q2447 AND symb_decoder(16#ae#)) OR
 					(reg_q2447 AND symb_decoder(16#55#)) OR
 					(reg_q2447 AND symb_decoder(16#36#)) OR
 					(reg_q2447 AND symb_decoder(16#44#)) OR
 					(reg_q2447 AND symb_decoder(16#7b#)) OR
 					(reg_q2447 AND symb_decoder(16#4f#)) OR
 					(reg_q2447 AND symb_decoder(16#15#)) OR
 					(reg_q2447 AND symb_decoder(16#67#)) OR
 					(reg_q2447 AND symb_decoder(16#8a#)) OR
 					(reg_q2447 AND symb_decoder(16#03#)) OR
 					(reg_q2447 AND symb_decoder(16#cf#)) OR
 					(reg_q2447 AND symb_decoder(16#2f#)) OR
 					(reg_q2447 AND symb_decoder(16#30#)) OR
 					(reg_q2447 AND symb_decoder(16#43#)) OR
 					(reg_q2447 AND symb_decoder(16#bc#)) OR
 					(reg_q2447 AND symb_decoder(16#59#)) OR
 					(reg_q2447 AND symb_decoder(16#63#)) OR
 					(reg_q2447 AND symb_decoder(16#f8#)) OR
 					(reg_q2447 AND symb_decoder(16#11#)) OR
 					(reg_q2447 AND symb_decoder(16#52#)) OR
 					(reg_q2447 AND symb_decoder(16#13#)) OR
 					(reg_q2447 AND symb_decoder(16#a2#)) OR
 					(reg_q2447 AND symb_decoder(16#40#)) OR
 					(reg_q2447 AND symb_decoder(16#8d#)) OR
 					(reg_q2447 AND symb_decoder(16#92#)) OR
 					(reg_q2447 AND symb_decoder(16#9a#)) OR
 					(reg_q2447 AND symb_decoder(16#7f#)) OR
 					(reg_q2447 AND symb_decoder(16#f3#)) OR
 					(reg_q2447 AND symb_decoder(16#ad#)) OR
 					(reg_q2447 AND symb_decoder(16#af#)) OR
 					(reg_q2447 AND symb_decoder(16#56#)) OR
 					(reg_q2447 AND symb_decoder(16#ac#)) OR
 					(reg_q2447 AND symb_decoder(16#b5#)) OR
 					(reg_q2447 AND symb_decoder(16#e4#)) OR
 					(reg_q2447 AND symb_decoder(16#b3#)) OR
 					(reg_q2447 AND symb_decoder(16#ef#)) OR
 					(reg_q2447 AND symb_decoder(16#b2#)) OR
 					(reg_q2447 AND symb_decoder(16#41#)) OR
 					(reg_q2447 AND symb_decoder(16#b9#)) OR
 					(reg_q2447 AND symb_decoder(16#62#)) OR
 					(reg_q2447 AND symb_decoder(16#ca#)) OR
 					(reg_q2447 AND symb_decoder(16#61#)) OR
 					(reg_q2447 AND symb_decoder(16#fa#)) OR
 					(reg_q2447 AND symb_decoder(16#ab#)) OR
 					(reg_q2447 AND symb_decoder(16#70#)) OR
 					(reg_q2447 AND symb_decoder(16#07#)) OR
 					(reg_q2447 AND symb_decoder(16#38#)) OR
 					(reg_q2447 AND symb_decoder(16#9b#)) OR
 					(reg_q2447 AND symb_decoder(16#1d#)) OR
 					(reg_q2447 AND symb_decoder(16#b0#)) OR
 					(reg_q2447 AND symb_decoder(16#3d#)) OR
 					(reg_q2447 AND symb_decoder(16#f5#)) OR
 					(reg_q2447 AND symb_decoder(16#7e#)) OR
 					(reg_q2447 AND symb_decoder(16#b7#)) OR
 					(reg_q2447 AND symb_decoder(16#1a#)) OR
 					(reg_q2447 AND symb_decoder(16#1b#)) OR
 					(reg_q2447 AND symb_decoder(16#4b#)) OR
 					(reg_q2447 AND symb_decoder(16#c6#)) OR
 					(reg_q2447 AND symb_decoder(16#95#)) OR
 					(reg_q2447 AND symb_decoder(16#10#)) OR
 					(reg_q2447 AND symb_decoder(16#a8#)) OR
 					(reg_q2447 AND symb_decoder(16#f1#)) OR
 					(reg_q2447 AND symb_decoder(16#9c#)) OR
 					(reg_q2447 AND symb_decoder(16#cb#)) OR
 					(reg_q2447 AND symb_decoder(16#00#)) OR
 					(reg_q2447 AND symb_decoder(16#75#)) OR
 					(reg_q2447 AND symb_decoder(16#57#)) OR
 					(reg_q2447 AND symb_decoder(16#8f#)) OR
 					(reg_q2447 AND symb_decoder(16#dd#)) OR
 					(reg_q2447 AND symb_decoder(16#80#)) OR
 					(reg_q2447 AND symb_decoder(16#d0#)) OR
 					(reg_q2447 AND symb_decoder(16#34#)) OR
 					(reg_q2447 AND symb_decoder(16#df#)) OR
 					(reg_q2447 AND symb_decoder(16#91#)) OR
 					(reg_q2447 AND symb_decoder(16#05#)) OR
 					(reg_q2447 AND symb_decoder(16#0c#)) OR
 					(reg_q2447 AND symb_decoder(16#02#)) OR
 					(reg_q2447 AND symb_decoder(16#c4#)) OR
 					(reg_q2447 AND symb_decoder(16#32#)) OR
 					(reg_q2447 AND symb_decoder(16#c8#)) OR
 					(reg_q2447 AND symb_decoder(16#c3#)) OR
 					(reg_q2447 AND symb_decoder(16#a6#)) OR
 					(reg_q2447 AND symb_decoder(16#e1#)) OR
 					(reg_q2447 AND symb_decoder(16#3a#)) OR
 					(reg_q2447 AND symb_decoder(16#09#)) OR
 					(reg_q2447 AND symb_decoder(16#01#)) OR
 					(reg_q2447 AND symb_decoder(16#90#)) OR
 					(reg_q2447 AND symb_decoder(16#b1#)) OR
 					(reg_q2447 AND symb_decoder(16#6e#)) OR
 					(reg_q2447 AND symb_decoder(16#16#)) OR
 					(reg_q2447 AND symb_decoder(16#21#)) OR
 					(reg_q2447 AND symb_decoder(16#ea#)) OR
 					(reg_q2447 AND symb_decoder(16#9f#)) OR
 					(reg_q2447 AND symb_decoder(16#93#)) OR
 					(reg_q2447 AND symb_decoder(16#c2#)) OR
 					(reg_q2447 AND symb_decoder(16#e7#)) OR
 					(reg_q2447 AND symb_decoder(16#71#)) OR
 					(reg_q2447 AND symb_decoder(16#04#)) OR
 					(reg_q2447 AND symb_decoder(16#50#)) OR
 					(reg_q2447 AND symb_decoder(16#e6#)) OR
 					(reg_q2447 AND symb_decoder(16#1e#)) OR
 					(reg_q2447 AND symb_decoder(16#65#)) OR
 					(reg_q2447 AND symb_decoder(16#b4#)) OR
 					(reg_q2447 AND symb_decoder(16#6d#)) OR
 					(reg_q2447 AND symb_decoder(16#c5#)) OR
 					(reg_q2447 AND symb_decoder(16#dc#)) OR
 					(reg_q2447 AND symb_decoder(16#88#)) OR
 					(reg_q2447 AND symb_decoder(16#14#)) OR
 					(reg_q2447 AND symb_decoder(16#28#)) OR
 					(reg_q2447 AND symb_decoder(16#d6#)) OR
 					(reg_q2447 AND symb_decoder(16#7c#)) OR
 					(reg_q2447 AND symb_decoder(16#fd#)) OR
 					(reg_q2447 AND symb_decoder(16#a0#)) OR
 					(reg_q2447 AND symb_decoder(16#a7#)) OR
 					(reg_q2447 AND symb_decoder(16#4c#)) OR
 					(reg_q2447 AND symb_decoder(16#ba#)) OR
 					(reg_q2447 AND symb_decoder(16#2b#)) OR
 					(reg_q2447 AND symb_decoder(16#64#)) OR
 					(reg_q2447 AND symb_decoder(16#c7#)) OR
 					(reg_q2447 AND symb_decoder(16#aa#)) OR
 					(reg_q2447 AND symb_decoder(16#bd#)) OR
 					(reg_q2447 AND symb_decoder(16#a1#)) OR
 					(reg_q2447 AND symb_decoder(16#c1#)) OR
 					(reg_q2447 AND symb_decoder(16#d7#)) OR
 					(reg_q2447 AND symb_decoder(16#19#)) OR
 					(reg_q2447 AND symb_decoder(16#da#)) OR
 					(reg_q2447 AND symb_decoder(16#f6#)) OR
 					(reg_q2447 AND symb_decoder(16#77#)) OR
 					(reg_q2447 AND symb_decoder(16#d1#)) OR
 					(reg_q2447 AND symb_decoder(16#fb#)) OR
 					(reg_q2447 AND symb_decoder(16#83#)) OR
 					(reg_q2447 AND symb_decoder(16#a5#)) OR
 					(reg_q2447 AND symb_decoder(16#f9#)) OR
 					(reg_q2447 AND symb_decoder(16#1f#)) OR
 					(reg_q2447 AND symb_decoder(16#bf#)) OR
 					(reg_q2447 AND symb_decoder(16#eb#)) OR
 					(reg_q2447 AND symb_decoder(16#31#)) OR
 					(reg_q2447 AND symb_decoder(16#46#)) OR
 					(reg_q2447 AND symb_decoder(16#33#)) OR
 					(reg_q2447 AND symb_decoder(16#fc#)) OR
 					(reg_q2447 AND symb_decoder(16#ee#)) OR
 					(reg_q2447 AND symb_decoder(16#79#)) OR
 					(reg_q2447 AND symb_decoder(16#f4#)) OR
 					(reg_q2447 AND symb_decoder(16#42#)) OR
 					(reg_q2447 AND symb_decoder(16#e0#)) OR
 					(reg_q2447 AND symb_decoder(16#1c#)) OR
 					(reg_q2447 AND symb_decoder(16#a3#)) OR
 					(reg_q2447 AND symb_decoder(16#81#)) OR
 					(reg_q2447 AND symb_decoder(16#be#)) OR
 					(reg_q2447 AND symb_decoder(16#12#)) OR
 					(reg_q2447 AND symb_decoder(16#c0#)) OR
 					(reg_q2447 AND symb_decoder(16#54#)) OR
 					(reg_q2447 AND symb_decoder(16#8b#)) OR
 					(reg_q2447 AND symb_decoder(16#08#)) OR
 					(reg_q2447 AND symb_decoder(16#68#)) OR
 					(reg_q2447 AND symb_decoder(16#0f#)) OR
 					(reg_q2447 AND symb_decoder(16#6b#)) OR
 					(reg_q2447 AND symb_decoder(16#7d#)) OR
 					(reg_q2447 AND symb_decoder(16#49#)) OR
 					(reg_q2447 AND symb_decoder(16#47#)) OR
 					(reg_q2447 AND symb_decoder(16#37#)) OR
 					(reg_q2447 AND symb_decoder(16#f2#)) OR
 					(reg_q2447 AND symb_decoder(16#7a#)) OR
 					(reg_q2447 AND symb_decoder(16#35#)) OR
 					(reg_q2447 AND symb_decoder(16#87#)) OR
 					(reg_q2447 AND symb_decoder(16#5a#)) OR
 					(reg_q2447 AND symb_decoder(16#60#)) OR
 					(reg_q2447 AND symb_decoder(16#d5#)) OR
 					(reg_q2447 AND symb_decoder(16#e8#)) OR
 					(reg_q2447 AND symb_decoder(16#27#)) OR
 					(reg_q2447 AND symb_decoder(16#ff#)) OR
 					(reg_q2447 AND symb_decoder(16#5c#)) OR
 					(reg_q2447 AND symb_decoder(16#e3#)) OR
 					(reg_q2447 AND symb_decoder(16#3e#)) OR
 					(reg_q2447 AND symb_decoder(16#99#)) OR
 					(reg_q2447 AND symb_decoder(16#2d#)) OR
 					(reg_q2447 AND symb_decoder(16#86#)) OR
 					(reg_q2447 AND symb_decoder(16#48#)) OR
 					(reg_q2447 AND symb_decoder(16#74#)) OR
 					(reg_q2447 AND symb_decoder(16#78#)) OR
 					(reg_q2447 AND symb_decoder(16#4d#)) OR
 					(reg_q2447 AND symb_decoder(16#2c#)) OR
 					(reg_q2447 AND symb_decoder(16#84#)) OR
 					(reg_q2447 AND symb_decoder(16#cd#));
reg_q773_in <= (reg_q772 AND symb_decoder(16#0a#)) OR
 					(reg_q772 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#));
reg_q472_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q471 AND symb_decoder(16#53#)) OR
 					(reg_q471 AND symb_decoder(16#73#));
reg_fullgraph22_init <= "00";

reg_fullgraph22_sel <= "0" & reg_q472_in & reg_q773_in & reg_q2447_in;

	--coder fullgraph22
with reg_fullgraph22_sel select
reg_fullgraph22_in <=
	"01" when "0001",
	"10" when "0010",
	"11" when "0100",
	"00" when others;
 --end coder

	p_reg_fullgraph22: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph22 <= reg_fullgraph22_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph22 <= reg_fullgraph22_init;
        else
          reg_fullgraph22 <= reg_fullgraph22_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph22

		reg_q2447 <= '1' when reg_fullgraph22 = "01" else '0'; 
		reg_q773 <= '1' when reg_fullgraph22 = "10" else '0'; 
		reg_q472 <= '1' when reg_fullgraph22 = "11" else '0'; 
--end decoder 

reg_q1218_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1218 AND symb_decoder(16#f5#)) OR
 					(reg_q1218 AND symb_decoder(16#9d#)) OR
 					(reg_q1218 AND symb_decoder(16#f3#)) OR
 					(reg_q1218 AND symb_decoder(16#f9#)) OR
 					(reg_q1218 AND symb_decoder(16#8f#)) OR
 					(reg_q1218 AND symb_decoder(16#12#)) OR
 					(reg_q1218 AND symb_decoder(16#09#)) OR
 					(reg_q1218 AND symb_decoder(16#81#)) OR
 					(reg_q1218 AND symb_decoder(16#84#)) OR
 					(reg_q1218 AND symb_decoder(16#c0#)) OR
 					(reg_q1218 AND symb_decoder(16#ce#)) OR
 					(reg_q1218 AND symb_decoder(16#31#)) OR
 					(reg_q1218 AND symb_decoder(16#b1#)) OR
 					(reg_q1218 AND symb_decoder(16#89#)) OR
 					(reg_q1218 AND symb_decoder(16#04#)) OR
 					(reg_q1218 AND symb_decoder(16#af#)) OR
 					(reg_q1218 AND symb_decoder(16#01#)) OR
 					(reg_q1218 AND symb_decoder(16#ec#)) OR
 					(reg_q1218 AND symb_decoder(16#cc#)) OR
 					(reg_q1218 AND symb_decoder(16#b3#)) OR
 					(reg_q1218 AND symb_decoder(16#de#)) OR
 					(reg_q1218 AND symb_decoder(16#0d#)) OR
 					(reg_q1218 AND symb_decoder(16#0f#)) OR
 					(reg_q1218 AND symb_decoder(16#e9#)) OR
 					(reg_q1218 AND symb_decoder(16#b5#)) OR
 					(reg_q1218 AND symb_decoder(16#2b#)) OR
 					(reg_q1218 AND symb_decoder(16#70#)) OR
 					(reg_q1218 AND symb_decoder(16#4f#)) OR
 					(reg_q1218 AND symb_decoder(16#ab#)) OR
 					(reg_q1218 AND symb_decoder(16#67#)) OR
 					(reg_q1218 AND symb_decoder(16#8b#)) OR
 					(reg_q1218 AND symb_decoder(16#15#)) OR
 					(reg_q1218 AND symb_decoder(16#07#)) OR
 					(reg_q1218 AND symb_decoder(16#10#)) OR
 					(reg_q1218 AND symb_decoder(16#dc#)) OR
 					(reg_q1218 AND symb_decoder(16#df#)) OR
 					(reg_q1218 AND symb_decoder(16#e3#)) OR
 					(reg_q1218 AND symb_decoder(16#23#)) OR
 					(reg_q1218 AND symb_decoder(16#ef#)) OR
 					(reg_q1218 AND symb_decoder(16#c5#)) OR
 					(reg_q1218 AND symb_decoder(16#cd#)) OR
 					(reg_q1218 AND symb_decoder(16#d4#)) OR
 					(reg_q1218 AND symb_decoder(16#bf#)) OR
 					(reg_q1218 AND symb_decoder(16#3f#)) OR
 					(reg_q1218 AND symb_decoder(16#4c#)) OR
 					(reg_q1218 AND symb_decoder(16#63#)) OR
 					(reg_q1218 AND symb_decoder(16#4e#)) OR
 					(reg_q1218 AND symb_decoder(16#7b#)) OR
 					(reg_q1218 AND symb_decoder(16#14#)) OR
 					(reg_q1218 AND symb_decoder(16#03#)) OR
 					(reg_q1218 AND symb_decoder(16#2c#)) OR
 					(reg_q1218 AND symb_decoder(16#65#)) OR
 					(reg_q1218 AND symb_decoder(16#0e#)) OR
 					(reg_q1218 AND symb_decoder(16#71#)) OR
 					(reg_q1218 AND symb_decoder(16#f1#)) OR
 					(reg_q1218 AND symb_decoder(16#fc#)) OR
 					(reg_q1218 AND symb_decoder(16#6a#)) OR
 					(reg_q1218 AND symb_decoder(16#5a#)) OR
 					(reg_q1218 AND symb_decoder(16#e5#)) OR
 					(reg_q1218 AND symb_decoder(16#58#)) OR
 					(reg_q1218 AND symb_decoder(16#87#)) OR
 					(reg_q1218 AND symb_decoder(16#a1#)) OR
 					(reg_q1218 AND symb_decoder(16#9a#)) OR
 					(reg_q1218 AND symb_decoder(16#3b#)) OR
 					(reg_q1218 AND symb_decoder(16#f2#)) OR
 					(reg_q1218 AND symb_decoder(16#8a#)) OR
 					(reg_q1218 AND symb_decoder(16#a3#)) OR
 					(reg_q1218 AND symb_decoder(16#45#)) OR
 					(reg_q1218 AND symb_decoder(16#78#)) OR
 					(reg_q1218 AND symb_decoder(16#7d#)) OR
 					(reg_q1218 AND symb_decoder(16#9b#)) OR
 					(reg_q1218 AND symb_decoder(16#c4#)) OR
 					(reg_q1218 AND symb_decoder(16#e0#)) OR
 					(reg_q1218 AND symb_decoder(16#c2#)) OR
 					(reg_q1218 AND symb_decoder(16#d3#)) OR
 					(reg_q1218 AND symb_decoder(16#3e#)) OR
 					(reg_q1218 AND symb_decoder(16#18#)) OR
 					(reg_q1218 AND symb_decoder(16#08#)) OR
 					(reg_q1218 AND symb_decoder(16#61#)) OR
 					(reg_q1218 AND symb_decoder(16#60#)) OR
 					(reg_q1218 AND symb_decoder(16#a2#)) OR
 					(reg_q1218 AND symb_decoder(16#59#)) OR
 					(reg_q1218 AND symb_decoder(16#d9#)) OR
 					(reg_q1218 AND symb_decoder(16#eb#)) OR
 					(reg_q1218 AND symb_decoder(16#5b#)) OR
 					(reg_q1218 AND symb_decoder(16#6e#)) OR
 					(reg_q1218 AND symb_decoder(16#16#)) OR
 					(reg_q1218 AND symb_decoder(16#99#)) OR
 					(reg_q1218 AND symb_decoder(16#4a#)) OR
 					(reg_q1218 AND symb_decoder(16#29#)) OR
 					(reg_q1218 AND symb_decoder(16#1d#)) OR
 					(reg_q1218 AND symb_decoder(16#53#)) OR
 					(reg_q1218 AND symb_decoder(16#d7#)) OR
 					(reg_q1218 AND symb_decoder(16#38#)) OR
 					(reg_q1218 AND symb_decoder(16#f8#)) OR
 					(reg_q1218 AND symb_decoder(16#34#)) OR
 					(reg_q1218 AND symb_decoder(16#a0#)) OR
 					(reg_q1218 AND symb_decoder(16#ea#)) OR
 					(reg_q1218 AND symb_decoder(16#48#)) OR
 					(reg_q1218 AND symb_decoder(16#80#)) OR
 					(reg_q1218 AND symb_decoder(16#11#)) OR
 					(reg_q1218 AND symb_decoder(16#5d#)) OR
 					(reg_q1218 AND symb_decoder(16#5f#)) OR
 					(reg_q1218 AND symb_decoder(16#43#)) OR
 					(reg_q1218 AND symb_decoder(16#96#)) OR
 					(reg_q1218 AND symb_decoder(16#64#)) OR
 					(reg_q1218 AND symb_decoder(16#1f#)) OR
 					(reg_q1218 AND symb_decoder(16#bd#)) OR
 					(reg_q1218 AND symb_decoder(16#2f#)) OR
 					(reg_q1218 AND symb_decoder(16#1e#)) OR
 					(reg_q1218 AND symb_decoder(16#db#)) OR
 					(reg_q1218 AND symb_decoder(16#57#)) OR
 					(reg_q1218 AND symb_decoder(16#8c#)) OR
 					(reg_q1218 AND symb_decoder(16#ac#)) OR
 					(reg_q1218 AND symb_decoder(16#f6#)) OR
 					(reg_q1218 AND symb_decoder(16#aa#)) OR
 					(reg_q1218 AND symb_decoder(16#e7#)) OR
 					(reg_q1218 AND symb_decoder(16#52#)) OR
 					(reg_q1218 AND symb_decoder(16#d1#)) OR
 					(reg_q1218 AND symb_decoder(16#21#)) OR
 					(reg_q1218 AND symb_decoder(16#a4#)) OR
 					(reg_q1218 AND symb_decoder(16#fe#)) OR
 					(reg_q1218 AND symb_decoder(16#6f#)) OR
 					(reg_q1218 AND symb_decoder(16#b6#)) OR
 					(reg_q1218 AND symb_decoder(16#90#)) OR
 					(reg_q1218 AND symb_decoder(16#3a#)) OR
 					(reg_q1218 AND symb_decoder(16#02#)) OR
 					(reg_q1218 AND symb_decoder(16#b0#)) OR
 					(reg_q1218 AND symb_decoder(16#a6#)) OR
 					(reg_q1218 AND symb_decoder(16#30#)) OR
 					(reg_q1218 AND symb_decoder(16#13#)) OR
 					(reg_q1218 AND symb_decoder(16#98#)) OR
 					(reg_q1218 AND symb_decoder(16#51#)) OR
 					(reg_q1218 AND symb_decoder(16#bc#)) OR
 					(reg_q1218 AND symb_decoder(16#e6#)) OR
 					(reg_q1218 AND symb_decoder(16#55#)) OR
 					(reg_q1218 AND symb_decoder(16#b9#)) OR
 					(reg_q1218 AND symb_decoder(16#92#)) OR
 					(reg_q1218 AND symb_decoder(16#d0#)) OR
 					(reg_q1218 AND symb_decoder(16#7e#)) OR
 					(reg_q1218 AND symb_decoder(16#fd#)) OR
 					(reg_q1218 AND symb_decoder(16#a8#)) OR
 					(reg_q1218 AND symb_decoder(16#26#)) OR
 					(reg_q1218 AND symb_decoder(16#b2#)) OR
 					(reg_q1218 AND symb_decoder(16#82#)) OR
 					(reg_q1218 AND symb_decoder(16#76#)) OR
 					(reg_q1218 AND symb_decoder(16#ca#)) OR
 					(reg_q1218 AND symb_decoder(16#66#)) OR
 					(reg_q1218 AND symb_decoder(16#c3#)) OR
 					(reg_q1218 AND symb_decoder(16#33#)) OR
 					(reg_q1218 AND symb_decoder(16#a9#)) OR
 					(reg_q1218 AND symb_decoder(16#2e#)) OR
 					(reg_q1218 AND symb_decoder(16#72#)) OR
 					(reg_q1218 AND symb_decoder(16#9c#)) OR
 					(reg_q1218 AND symb_decoder(16#cf#)) OR
 					(reg_q1218 AND symb_decoder(16#5c#)) OR
 					(reg_q1218 AND symb_decoder(16#39#)) OR
 					(reg_q1218 AND symb_decoder(16#0b#)) OR
 					(reg_q1218 AND symb_decoder(16#c7#)) OR
 					(reg_q1218 AND symb_decoder(16#ff#)) OR
 					(reg_q1218 AND symb_decoder(16#24#)) OR
 					(reg_q1218 AND symb_decoder(16#a7#)) OR
 					(reg_q1218 AND symb_decoder(16#69#)) OR
 					(reg_q1218 AND symb_decoder(16#85#)) OR
 					(reg_q1218 AND symb_decoder(16#f7#)) OR
 					(reg_q1218 AND symb_decoder(16#40#)) OR
 					(reg_q1218 AND symb_decoder(16#c9#)) OR
 					(reg_q1218 AND symb_decoder(16#1c#)) OR
 					(reg_q1218 AND symb_decoder(16#0c#)) OR
 					(reg_q1218 AND symb_decoder(16#79#)) OR
 					(reg_q1218 AND symb_decoder(16#3d#)) OR
 					(reg_q1218 AND symb_decoder(16#95#)) OR
 					(reg_q1218 AND symb_decoder(16#b7#)) OR
 					(reg_q1218 AND symb_decoder(16#91#)) OR
 					(reg_q1218 AND symb_decoder(16#1b#)) OR
 					(reg_q1218 AND symb_decoder(16#e1#)) OR
 					(reg_q1218 AND symb_decoder(16#35#)) OR
 					(reg_q1218 AND symb_decoder(16#62#)) OR
 					(reg_q1218 AND symb_decoder(16#9f#)) OR
 					(reg_q1218 AND symb_decoder(16#6c#)) OR
 					(reg_q1218 AND symb_decoder(16#8e#)) OR
 					(reg_q1218 AND symb_decoder(16#22#)) OR
 					(reg_q1218 AND symb_decoder(16#17#)) OR
 					(reg_q1218 AND symb_decoder(16#32#)) OR
 					(reg_q1218 AND symb_decoder(16#7f#)) OR
 					(reg_q1218 AND symb_decoder(16#e2#)) OR
 					(reg_q1218 AND symb_decoder(16#b8#)) OR
 					(reg_q1218 AND symb_decoder(16#97#)) OR
 					(reg_q1218 AND symb_decoder(16#d6#)) OR
 					(reg_q1218 AND symb_decoder(16#28#)) OR
 					(reg_q1218 AND symb_decoder(16#68#)) OR
 					(reg_q1218 AND symb_decoder(16#37#)) OR
 					(reg_q1218 AND symb_decoder(16#bb#)) OR
 					(reg_q1218 AND symb_decoder(16#fb#)) OR
 					(reg_q1218 AND symb_decoder(16#88#)) OR
 					(reg_q1218 AND symb_decoder(16#27#)) OR
 					(reg_q1218 AND symb_decoder(16#44#)) OR
 					(reg_q1218 AND symb_decoder(16#77#)) OR
 					(reg_q1218 AND symb_decoder(16#7c#)) OR
 					(reg_q1218 AND symb_decoder(16#ae#)) OR
 					(reg_q1218 AND symb_decoder(16#4b#)) OR
 					(reg_q1218 AND symb_decoder(16#da#)) OR
 					(reg_q1218 AND symb_decoder(16#1a#)) OR
 					(reg_q1218 AND symb_decoder(16#3c#)) OR
 					(reg_q1218 AND symb_decoder(16#ed#)) OR
 					(reg_q1218 AND symb_decoder(16#05#)) OR
 					(reg_q1218 AND symb_decoder(16#d2#)) OR
 					(reg_q1218 AND symb_decoder(16#00#)) OR
 					(reg_q1218 AND symb_decoder(16#36#)) OR
 					(reg_q1218 AND symb_decoder(16#ad#)) OR
 					(reg_q1218 AND symb_decoder(16#fa#)) OR
 					(reg_q1218 AND symb_decoder(16#8d#)) OR
 					(reg_q1218 AND symb_decoder(16#2a#)) OR
 					(reg_q1218 AND symb_decoder(16#b4#)) OR
 					(reg_q1218 AND symb_decoder(16#ee#)) OR
 					(reg_q1218 AND symb_decoder(16#f0#)) OR
 					(reg_q1218 AND symb_decoder(16#74#)) OR
 					(reg_q1218 AND symb_decoder(16#49#)) OR
 					(reg_q1218 AND symb_decoder(16#41#)) OR
 					(reg_q1218 AND symb_decoder(16#93#)) OR
 					(reg_q1218 AND symb_decoder(16#c6#)) OR
 					(reg_q1218 AND symb_decoder(16#5e#)) OR
 					(reg_q1218 AND symb_decoder(16#7a#)) OR
 					(reg_q1218 AND symb_decoder(16#83#)) OR
 					(reg_q1218 AND symb_decoder(16#c1#)) OR
 					(reg_q1218 AND symb_decoder(16#06#)) OR
 					(reg_q1218 AND symb_decoder(16#f4#)) OR
 					(reg_q1218 AND symb_decoder(16#42#)) OR
 					(reg_q1218 AND symb_decoder(16#cb#)) OR
 					(reg_q1218 AND symb_decoder(16#25#)) OR
 					(reg_q1218 AND symb_decoder(16#dd#)) OR
 					(reg_q1218 AND symb_decoder(16#4d#)) OR
 					(reg_q1218 AND symb_decoder(16#94#)) OR
 					(reg_q1218 AND symb_decoder(16#54#)) OR
 					(reg_q1218 AND symb_decoder(16#c8#)) OR
 					(reg_q1218 AND symb_decoder(16#0a#)) OR
 					(reg_q1218 AND symb_decoder(16#86#)) OR
 					(reg_q1218 AND symb_decoder(16#2d#)) OR
 					(reg_q1218 AND symb_decoder(16#73#)) OR
 					(reg_q1218 AND symb_decoder(16#6b#)) OR
 					(reg_q1218 AND symb_decoder(16#19#)) OR
 					(reg_q1218 AND symb_decoder(16#be#)) OR
 					(reg_q1218 AND symb_decoder(16#75#)) OR
 					(reg_q1218 AND symb_decoder(16#a5#)) OR
 					(reg_q1218 AND symb_decoder(16#d8#)) OR
 					(reg_q1218 AND symb_decoder(16#47#)) OR
 					(reg_q1218 AND symb_decoder(16#20#)) OR
 					(reg_q1218 AND symb_decoder(16#d5#)) OR
 					(reg_q1218 AND symb_decoder(16#e4#)) OR
 					(reg_q1218 AND symb_decoder(16#e8#)) OR
 					(reg_q1218 AND symb_decoder(16#46#)) OR
 					(reg_q1218 AND symb_decoder(16#ba#)) OR
 					(reg_q1218 AND symb_decoder(16#50#)) OR
 					(reg_q1218 AND symb_decoder(16#56#)) OR
 					(reg_q1218 AND symb_decoder(16#9e#)) OR
 					(reg_q1218 AND symb_decoder(16#6d#));
reg_q1218_init <= '0' ;
	p_reg_q1218: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1218 <= reg_q1218_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1218 <= reg_q1218_init;
        else
          reg_q1218 <= reg_q1218_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1061_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1061 AND symb_decoder(16#ee#)) OR
 					(reg_q1061 AND symb_decoder(16#2c#)) OR
 					(reg_q1061 AND symb_decoder(16#45#)) OR
 					(reg_q1061 AND symb_decoder(16#72#)) OR
 					(reg_q1061 AND symb_decoder(16#e3#)) OR
 					(reg_q1061 AND symb_decoder(16#fa#)) OR
 					(reg_q1061 AND symb_decoder(16#89#)) OR
 					(reg_q1061 AND symb_decoder(16#29#)) OR
 					(reg_q1061 AND symb_decoder(16#7f#)) OR
 					(reg_q1061 AND symb_decoder(16#c2#)) OR
 					(reg_q1061 AND symb_decoder(16#79#)) OR
 					(reg_q1061 AND symb_decoder(16#81#)) OR
 					(reg_q1061 AND symb_decoder(16#25#)) OR
 					(reg_q1061 AND symb_decoder(16#35#)) OR
 					(reg_q1061 AND symb_decoder(16#08#)) OR
 					(reg_q1061 AND symb_decoder(16#d3#)) OR
 					(reg_q1061 AND symb_decoder(16#a6#)) OR
 					(reg_q1061 AND symb_decoder(16#a2#)) OR
 					(reg_q1061 AND symb_decoder(16#6b#)) OR
 					(reg_q1061 AND symb_decoder(16#71#)) OR
 					(reg_q1061 AND symb_decoder(16#37#)) OR
 					(reg_q1061 AND symb_decoder(16#06#)) OR
 					(reg_q1061 AND symb_decoder(16#95#)) OR
 					(reg_q1061 AND symb_decoder(16#18#)) OR
 					(reg_q1061 AND symb_decoder(16#57#)) OR
 					(reg_q1061 AND symb_decoder(16#7e#)) OR
 					(reg_q1061 AND symb_decoder(16#f2#)) OR
 					(reg_q1061 AND symb_decoder(16#43#)) OR
 					(reg_q1061 AND symb_decoder(16#93#)) OR
 					(reg_q1061 AND symb_decoder(16#68#)) OR
 					(reg_q1061 AND symb_decoder(16#f8#)) OR
 					(reg_q1061 AND symb_decoder(16#3b#)) OR
 					(reg_q1061 AND symb_decoder(16#28#)) OR
 					(reg_q1061 AND symb_decoder(16#ca#)) OR
 					(reg_q1061 AND symb_decoder(16#ba#)) OR
 					(reg_q1061 AND symb_decoder(16#1c#)) OR
 					(reg_q1061 AND symb_decoder(16#44#)) OR
 					(reg_q1061 AND symb_decoder(16#76#)) OR
 					(reg_q1061 AND symb_decoder(16#05#)) OR
 					(reg_q1061 AND symb_decoder(16#f1#)) OR
 					(reg_q1061 AND symb_decoder(16#3d#)) OR
 					(reg_q1061 AND symb_decoder(16#ae#)) OR
 					(reg_q1061 AND symb_decoder(16#38#)) OR
 					(reg_q1061 AND symb_decoder(16#02#)) OR
 					(reg_q1061 AND symb_decoder(16#ec#)) OR
 					(reg_q1061 AND symb_decoder(16#26#)) OR
 					(reg_q1061 AND symb_decoder(16#61#)) OR
 					(reg_q1061 AND symb_decoder(16#70#)) OR
 					(reg_q1061 AND symb_decoder(16#84#)) OR
 					(reg_q1061 AND symb_decoder(16#34#)) OR
 					(reg_q1061 AND symb_decoder(16#85#)) OR
 					(reg_q1061 AND symb_decoder(16#eb#)) OR
 					(reg_q1061 AND symb_decoder(16#8e#)) OR
 					(reg_q1061 AND symb_decoder(16#60#)) OR
 					(reg_q1061 AND symb_decoder(16#9c#)) OR
 					(reg_q1061 AND symb_decoder(16#83#)) OR
 					(reg_q1061 AND symb_decoder(16#3c#)) OR
 					(reg_q1061 AND symb_decoder(16#32#)) OR
 					(reg_q1061 AND symb_decoder(16#49#)) OR
 					(reg_q1061 AND symb_decoder(16#be#)) OR
 					(reg_q1061 AND symb_decoder(16#52#)) OR
 					(reg_q1061 AND symb_decoder(16#de#)) OR
 					(reg_q1061 AND symb_decoder(16#f3#)) OR
 					(reg_q1061 AND symb_decoder(16#f6#)) OR
 					(reg_q1061 AND symb_decoder(16#a5#)) OR
 					(reg_q1061 AND symb_decoder(16#36#)) OR
 					(reg_q1061 AND symb_decoder(16#03#)) OR
 					(reg_q1061 AND symb_decoder(16#62#)) OR
 					(reg_q1061 AND symb_decoder(16#c9#)) OR
 					(reg_q1061 AND symb_decoder(16#16#)) OR
 					(reg_q1061 AND symb_decoder(16#7a#)) OR
 					(reg_q1061 AND symb_decoder(16#dd#)) OR
 					(reg_q1061 AND symb_decoder(16#87#)) OR
 					(reg_q1061 AND symb_decoder(16#0c#)) OR
 					(reg_q1061 AND symb_decoder(16#ff#)) OR
 					(reg_q1061 AND symb_decoder(16#aa#)) OR
 					(reg_q1061 AND symb_decoder(16#a3#)) OR
 					(reg_q1061 AND symb_decoder(16#65#)) OR
 					(reg_q1061 AND symb_decoder(16#59#)) OR
 					(reg_q1061 AND symb_decoder(16#50#)) OR
 					(reg_q1061 AND symb_decoder(16#64#)) OR
 					(reg_q1061 AND symb_decoder(16#8b#)) OR
 					(reg_q1061 AND symb_decoder(16#4f#)) OR
 					(reg_q1061 AND symb_decoder(16#c5#)) OR
 					(reg_q1061 AND symb_decoder(16#7d#)) OR
 					(reg_q1061 AND symb_decoder(16#ea#)) OR
 					(reg_q1061 AND symb_decoder(16#ac#)) OR
 					(reg_q1061 AND symb_decoder(16#9f#)) OR
 					(reg_q1061 AND symb_decoder(16#4d#)) OR
 					(reg_q1061 AND symb_decoder(16#98#)) OR
 					(reg_q1061 AND symb_decoder(16#bf#)) OR
 					(reg_q1061 AND symb_decoder(16#1b#)) OR
 					(reg_q1061 AND symb_decoder(16#2b#)) OR
 					(reg_q1061 AND symb_decoder(16#9a#)) OR
 					(reg_q1061 AND symb_decoder(16#19#)) OR
 					(reg_q1061 AND symb_decoder(16#a0#)) OR
 					(reg_q1061 AND symb_decoder(16#c4#)) OR
 					(reg_q1061 AND symb_decoder(16#8d#)) OR
 					(reg_q1061 AND symb_decoder(16#c6#)) OR
 					(reg_q1061 AND symb_decoder(16#0d#)) OR
 					(reg_q1061 AND symb_decoder(16#b5#)) OR
 					(reg_q1061 AND symb_decoder(16#d5#)) OR
 					(reg_q1061 AND symb_decoder(16#f0#)) OR
 					(reg_q1061 AND symb_decoder(16#74#)) OR
 					(reg_q1061 AND symb_decoder(16#8f#)) OR
 					(reg_q1061 AND symb_decoder(16#00#)) OR
 					(reg_q1061 AND symb_decoder(16#dc#)) OR
 					(reg_q1061 AND symb_decoder(16#17#)) OR
 					(reg_q1061 AND symb_decoder(16#5c#)) OR
 					(reg_q1061 AND symb_decoder(16#63#)) OR
 					(reg_q1061 AND symb_decoder(16#b3#)) OR
 					(reg_q1061 AND symb_decoder(16#d1#)) OR
 					(reg_q1061 AND symb_decoder(16#b7#)) OR
 					(reg_q1061 AND symb_decoder(16#bd#)) OR
 					(reg_q1061 AND symb_decoder(16#c7#)) OR
 					(reg_q1061 AND symb_decoder(16#d0#)) OR
 					(reg_q1061 AND symb_decoder(16#47#)) OR
 					(reg_q1061 AND symb_decoder(16#1f#)) OR
 					(reg_q1061 AND symb_decoder(16#a9#)) OR
 					(reg_q1061 AND symb_decoder(16#3e#)) OR
 					(reg_q1061 AND symb_decoder(16#b9#)) OR
 					(reg_q1061 AND symb_decoder(16#f7#)) OR
 					(reg_q1061 AND symb_decoder(16#f5#)) OR
 					(reg_q1061 AND symb_decoder(16#6d#)) OR
 					(reg_q1061 AND symb_decoder(16#20#)) OR
 					(reg_q1061 AND symb_decoder(16#91#)) OR
 					(reg_q1061 AND symb_decoder(16#9e#)) OR
 					(reg_q1061 AND symb_decoder(16#12#)) OR
 					(reg_q1061 AND symb_decoder(16#bb#)) OR
 					(reg_q1061 AND symb_decoder(16#0f#)) OR
 					(reg_q1061 AND symb_decoder(16#4a#)) OR
 					(reg_q1061 AND symb_decoder(16#df#)) OR
 					(reg_q1061 AND symb_decoder(16#41#)) OR
 					(reg_q1061 AND symb_decoder(16#90#)) OR
 					(reg_q1061 AND symb_decoder(16#fd#)) OR
 					(reg_q1061 AND symb_decoder(16#fe#)) OR
 					(reg_q1061 AND symb_decoder(16#b4#)) OR
 					(reg_q1061 AND symb_decoder(16#ce#)) OR
 					(reg_q1061 AND symb_decoder(16#31#)) OR
 					(reg_q1061 AND symb_decoder(16#8a#)) OR
 					(reg_q1061 AND symb_decoder(16#cc#)) OR
 					(reg_q1061 AND symb_decoder(16#9b#)) OR
 					(reg_q1061 AND symb_decoder(16#1d#)) OR
 					(reg_q1061 AND symb_decoder(16#80#)) OR
 					(reg_q1061 AND symb_decoder(16#13#)) OR
 					(reg_q1061 AND symb_decoder(16#a4#)) OR
 					(reg_q1061 AND symb_decoder(16#94#)) OR
 					(reg_q1061 AND symb_decoder(16#42#)) OR
 					(reg_q1061 AND symb_decoder(16#27#)) OR
 					(reg_q1061 AND symb_decoder(16#d8#)) OR
 					(reg_q1061 AND symb_decoder(16#0a#)) OR
 					(reg_q1061 AND symb_decoder(16#09#)) OR
 					(reg_q1061 AND symb_decoder(16#75#)) OR
 					(reg_q1061 AND symb_decoder(16#bc#)) OR
 					(reg_q1061 AND symb_decoder(16#a1#)) OR
 					(reg_q1061 AND symb_decoder(16#e1#)) OR
 					(reg_q1061 AND symb_decoder(16#f4#)) OR
 					(reg_q1061 AND symb_decoder(16#96#)) OR
 					(reg_q1061 AND symb_decoder(16#e8#)) OR
 					(reg_q1061 AND symb_decoder(16#e2#)) OR
 					(reg_q1061 AND symb_decoder(16#56#)) OR
 					(reg_q1061 AND symb_decoder(16#2d#)) OR
 					(reg_q1061 AND symb_decoder(16#b8#)) OR
 					(reg_q1061 AND symb_decoder(16#2f#)) OR
 					(reg_q1061 AND symb_decoder(16#23#)) OR
 					(reg_q1061 AND symb_decoder(16#54#)) OR
 					(reg_q1061 AND symb_decoder(16#ad#)) OR
 					(reg_q1061 AND symb_decoder(16#e9#)) OR
 					(reg_q1061 AND symb_decoder(16#e7#)) OR
 					(reg_q1061 AND symb_decoder(16#48#)) OR
 					(reg_q1061 AND symb_decoder(16#7c#)) OR
 					(reg_q1061 AND symb_decoder(16#53#)) OR
 					(reg_q1061 AND symb_decoder(16#55#)) OR
 					(reg_q1061 AND symb_decoder(16#1a#)) OR
 					(reg_q1061 AND symb_decoder(16#2e#)) OR
 					(reg_q1061 AND symb_decoder(16#2a#)) OR
 					(reg_q1061 AND symb_decoder(16#15#)) OR
 					(reg_q1061 AND symb_decoder(16#ab#)) OR
 					(reg_q1061 AND symb_decoder(16#78#)) OR
 					(reg_q1061 AND symb_decoder(16#7b#)) OR
 					(reg_q1061 AND symb_decoder(16#ef#)) OR
 					(reg_q1061 AND symb_decoder(16#11#)) OR
 					(reg_q1061 AND symb_decoder(16#da#)) OR
 					(reg_q1061 AND symb_decoder(16#22#)) OR
 					(reg_q1061 AND symb_decoder(16#fc#)) OR
 					(reg_q1061 AND symb_decoder(16#9d#)) OR
 					(reg_q1061 AND symb_decoder(16#b6#)) OR
 					(reg_q1061 AND symb_decoder(16#01#)) OR
 					(reg_q1061 AND symb_decoder(16#58#)) OR
 					(reg_q1061 AND symb_decoder(16#f9#)) OR
 					(reg_q1061 AND symb_decoder(16#07#)) OR
 					(reg_q1061 AND symb_decoder(16#51#)) OR
 					(reg_q1061 AND symb_decoder(16#4c#)) OR
 					(reg_q1061 AND symb_decoder(16#40#)) OR
 					(reg_q1061 AND symb_decoder(16#e6#)) OR
 					(reg_q1061 AND symb_decoder(16#86#)) OR
 					(reg_q1061 AND symb_decoder(16#c0#)) OR
 					(reg_q1061 AND symb_decoder(16#5e#)) OR
 					(reg_q1061 AND symb_decoder(16#b0#)) OR
 					(reg_q1061 AND symb_decoder(16#4e#)) OR
 					(reg_q1061 AND symb_decoder(16#82#)) OR
 					(reg_q1061 AND symb_decoder(16#ed#)) OR
 					(reg_q1061 AND symb_decoder(16#69#)) OR
 					(reg_q1061 AND symb_decoder(16#4b#)) OR
 					(reg_q1061 AND symb_decoder(16#92#)) OR
 					(reg_q1061 AND symb_decoder(16#88#)) OR
 					(reg_q1061 AND symb_decoder(16#e0#)) OR
 					(reg_q1061 AND symb_decoder(16#c3#)) OR
 					(reg_q1061 AND symb_decoder(16#30#)) OR
 					(reg_q1061 AND symb_decoder(16#97#)) OR
 					(reg_q1061 AND symb_decoder(16#6a#)) OR
 					(reg_q1061 AND symb_decoder(16#d2#)) OR
 					(reg_q1061 AND symb_decoder(16#b1#)) OR
 					(reg_q1061 AND symb_decoder(16#e5#)) OR
 					(reg_q1061 AND symb_decoder(16#10#)) OR
 					(reg_q1061 AND symb_decoder(16#a8#)) OR
 					(reg_q1061 AND symb_decoder(16#8c#)) OR
 					(reg_q1061 AND symb_decoder(16#73#)) OR
 					(reg_q1061 AND symb_decoder(16#24#)) OR
 					(reg_q1061 AND symb_decoder(16#3a#)) OR
 					(reg_q1061 AND symb_decoder(16#04#)) OR
 					(reg_q1061 AND symb_decoder(16#14#)) OR
 					(reg_q1061 AND symb_decoder(16#db#)) OR
 					(reg_q1061 AND symb_decoder(16#99#)) OR
 					(reg_q1061 AND symb_decoder(16#66#)) OR
 					(reg_q1061 AND symb_decoder(16#d4#)) OR
 					(reg_q1061 AND symb_decoder(16#39#)) OR
 					(reg_q1061 AND symb_decoder(16#cf#)) OR
 					(reg_q1061 AND symb_decoder(16#b2#)) OR
 					(reg_q1061 AND symb_decoder(16#e4#)) OR
 					(reg_q1061 AND symb_decoder(16#5f#)) OR
 					(reg_q1061 AND symb_decoder(16#cb#)) OR
 					(reg_q1061 AND symb_decoder(16#d7#)) OR
 					(reg_q1061 AND symb_decoder(16#5a#)) OR
 					(reg_q1061 AND symb_decoder(16#fb#)) OR
 					(reg_q1061 AND symb_decoder(16#6f#)) OR
 					(reg_q1061 AND symb_decoder(16#1e#)) OR
 					(reg_q1061 AND symb_decoder(16#46#)) OR
 					(reg_q1061 AND symb_decoder(16#a7#)) OR
 					(reg_q1061 AND symb_decoder(16#67#)) OR
 					(reg_q1061 AND symb_decoder(16#77#)) OR
 					(reg_q1061 AND symb_decoder(16#c8#)) OR
 					(reg_q1061 AND symb_decoder(16#33#)) OR
 					(reg_q1061 AND symb_decoder(16#6e#)) OR
 					(reg_q1061 AND symb_decoder(16#d6#)) OR
 					(reg_q1061 AND symb_decoder(16#5b#)) OR
 					(reg_q1061 AND symb_decoder(16#3f#)) OR
 					(reg_q1061 AND symb_decoder(16#21#)) OR
 					(reg_q1061 AND symb_decoder(16#d9#)) OR
 					(reg_q1061 AND symb_decoder(16#0e#)) OR
 					(reg_q1061 AND symb_decoder(16#af#)) OR
 					(reg_q1061 AND symb_decoder(16#0b#)) OR
 					(reg_q1061 AND symb_decoder(16#cd#)) OR
 					(reg_q1061 AND symb_decoder(16#c1#)) OR
 					(reg_q1061 AND symb_decoder(16#5d#)) OR
 					(reg_q1061 AND symb_decoder(16#6c#));
reg_q1061_init <= '0' ;
	p_reg_q1061: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1061 <= reg_q1061_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1061 <= reg_q1061_init;
        else
          reg_q1061 <= reg_q1061_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2449_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q2449 AND symb_decoder(16#bd#)) OR
 					(reg_q2449 AND symb_decoder(16#cf#)) OR
 					(reg_q2449 AND symb_decoder(16#61#)) OR
 					(reg_q2449 AND symb_decoder(16#79#)) OR
 					(reg_q2449 AND symb_decoder(16#47#)) OR
 					(reg_q2449 AND symb_decoder(16#f3#)) OR
 					(reg_q2449 AND symb_decoder(16#bf#)) OR
 					(reg_q2449 AND symb_decoder(16#69#)) OR
 					(reg_q2449 AND symb_decoder(16#cc#)) OR
 					(reg_q2449 AND symb_decoder(16#9c#)) OR
 					(reg_q2449 AND symb_decoder(16#95#)) OR
 					(reg_q2449 AND symb_decoder(16#46#)) OR
 					(reg_q2449 AND symb_decoder(16#13#)) OR
 					(reg_q2449 AND symb_decoder(16#b9#)) OR
 					(reg_q2449 AND symb_decoder(16#91#)) OR
 					(reg_q2449 AND symb_decoder(16#01#)) OR
 					(reg_q2449 AND symb_decoder(16#11#)) OR
 					(reg_q2449 AND symb_decoder(16#0f#)) OR
 					(reg_q2449 AND symb_decoder(16#96#)) OR
 					(reg_q2449 AND symb_decoder(16#24#)) OR
 					(reg_q2449 AND symb_decoder(16#6d#)) OR
 					(reg_q2449 AND symb_decoder(16#d7#)) OR
 					(reg_q2449 AND symb_decoder(16#e3#)) OR
 					(reg_q2449 AND symb_decoder(16#52#)) OR
 					(reg_q2449 AND symb_decoder(16#ed#)) OR
 					(reg_q2449 AND symb_decoder(16#1b#)) OR
 					(reg_q2449 AND symb_decoder(16#d9#)) OR
 					(reg_q2449 AND symb_decoder(16#dc#)) OR
 					(reg_q2449 AND symb_decoder(16#d0#)) OR
 					(reg_q2449 AND symb_decoder(16#c6#)) OR
 					(reg_q2449 AND symb_decoder(16#b4#)) OR
 					(reg_q2449 AND symb_decoder(16#ef#)) OR
 					(reg_q2449 AND symb_decoder(16#67#)) OR
 					(reg_q2449 AND symb_decoder(16#17#)) OR
 					(reg_q2449 AND symb_decoder(16#de#)) OR
 					(reg_q2449 AND symb_decoder(16#fa#)) OR
 					(reg_q2449 AND symb_decoder(16#31#)) OR
 					(reg_q2449 AND symb_decoder(16#e2#)) OR
 					(reg_q2449 AND symb_decoder(16#f0#)) OR
 					(reg_q2449 AND symb_decoder(16#a7#)) OR
 					(reg_q2449 AND symb_decoder(16#5e#)) OR
 					(reg_q2449 AND symb_decoder(16#b7#)) OR
 					(reg_q2449 AND symb_decoder(16#90#)) OR
 					(reg_q2449 AND symb_decoder(16#6f#)) OR
 					(reg_q2449 AND symb_decoder(16#a2#)) OR
 					(reg_q2449 AND symb_decoder(16#1c#)) OR
 					(reg_q2449 AND symb_decoder(16#7d#)) OR
 					(reg_q2449 AND symb_decoder(16#c8#)) OR
 					(reg_q2449 AND symb_decoder(16#4f#)) OR
 					(reg_q2449 AND symb_decoder(16#b1#)) OR
 					(reg_q2449 AND symb_decoder(16#40#)) OR
 					(reg_q2449 AND symb_decoder(16#19#)) OR
 					(reg_q2449 AND symb_decoder(16#da#)) OR
 					(reg_q2449 AND symb_decoder(16#db#)) OR
 					(reg_q2449 AND symb_decoder(16#9d#)) OR
 					(reg_q2449 AND symb_decoder(16#8f#)) OR
 					(reg_q2449 AND symb_decoder(16#26#)) OR
 					(reg_q2449 AND symb_decoder(16#55#)) OR
 					(reg_q2449 AND symb_decoder(16#4a#)) OR
 					(reg_q2449 AND symb_decoder(16#99#)) OR
 					(reg_q2449 AND symb_decoder(16#b5#)) OR
 					(reg_q2449 AND symb_decoder(16#18#)) OR
 					(reg_q2449 AND symb_decoder(16#5b#)) OR
 					(reg_q2449 AND symb_decoder(16#ba#)) OR
 					(reg_q2449 AND symb_decoder(16#27#)) OR
 					(reg_q2449 AND symb_decoder(16#92#)) OR
 					(reg_q2449 AND symb_decoder(16#4c#)) OR
 					(reg_q2449 AND symb_decoder(16#10#)) OR
 					(reg_q2449 AND symb_decoder(16#35#)) OR
 					(reg_q2449 AND symb_decoder(16#3c#)) OR
 					(reg_q2449 AND symb_decoder(16#45#)) OR
 					(reg_q2449 AND symb_decoder(16#d2#)) OR
 					(reg_q2449 AND symb_decoder(16#64#)) OR
 					(reg_q2449 AND symb_decoder(16#06#)) OR
 					(reg_q2449 AND symb_decoder(16#9b#)) OR
 					(reg_q2449 AND symb_decoder(16#3a#)) OR
 					(reg_q2449 AND symb_decoder(16#d5#)) OR
 					(reg_q2449 AND symb_decoder(16#fd#)) OR
 					(reg_q2449 AND symb_decoder(16#f4#)) OR
 					(reg_q2449 AND symb_decoder(16#4b#)) OR
 					(reg_q2449 AND symb_decoder(16#63#)) OR
 					(reg_q2449 AND symb_decoder(16#ca#)) OR
 					(reg_q2449 AND symb_decoder(16#3e#)) OR
 					(reg_q2449 AND symb_decoder(16#c2#)) OR
 					(reg_q2449 AND symb_decoder(16#89#)) OR
 					(reg_q2449 AND symb_decoder(16#0b#)) OR
 					(reg_q2449 AND symb_decoder(16#be#)) OR
 					(reg_q2449 AND symb_decoder(16#23#)) OR
 					(reg_q2449 AND symb_decoder(16#ae#)) OR
 					(reg_q2449 AND symb_decoder(16#a5#)) OR
 					(reg_q2449 AND symb_decoder(16#f8#)) OR
 					(reg_q2449 AND symb_decoder(16#07#)) OR
 					(reg_q2449 AND symb_decoder(16#05#)) OR
 					(reg_q2449 AND symb_decoder(16#f7#)) OR
 					(reg_q2449 AND symb_decoder(16#0a#)) OR
 					(reg_q2449 AND symb_decoder(16#30#)) OR
 					(reg_q2449 AND symb_decoder(16#00#)) OR
 					(reg_q2449 AND symb_decoder(16#76#)) OR
 					(reg_q2449 AND symb_decoder(16#ad#)) OR
 					(reg_q2449 AND symb_decoder(16#8e#)) OR
 					(reg_q2449 AND symb_decoder(16#d8#)) OR
 					(reg_q2449 AND symb_decoder(16#70#)) OR
 					(reg_q2449 AND symb_decoder(16#1d#)) OR
 					(reg_q2449 AND symb_decoder(16#ff#)) OR
 					(reg_q2449 AND symb_decoder(16#f2#)) OR
 					(reg_q2449 AND symb_decoder(16#62#)) OR
 					(reg_q2449 AND symb_decoder(16#41#)) OR
 					(reg_q2449 AND symb_decoder(16#81#)) OR
 					(reg_q2449 AND symb_decoder(16#2d#)) OR
 					(reg_q2449 AND symb_decoder(16#37#)) OR
 					(reg_q2449 AND symb_decoder(16#0c#)) OR
 					(reg_q2449 AND symb_decoder(16#c0#)) OR
 					(reg_q2449 AND symb_decoder(16#e5#)) OR
 					(reg_q2449 AND symb_decoder(16#f1#)) OR
 					(reg_q2449 AND symb_decoder(16#e1#)) OR
 					(reg_q2449 AND symb_decoder(16#4d#)) OR
 					(reg_q2449 AND symb_decoder(16#14#)) OR
 					(reg_q2449 AND symb_decoder(16#49#)) OR
 					(reg_q2449 AND symb_decoder(16#2c#)) OR
 					(reg_q2449 AND symb_decoder(16#53#)) OR
 					(reg_q2449 AND symb_decoder(16#42#)) OR
 					(reg_q2449 AND symb_decoder(16#bc#)) OR
 					(reg_q2449 AND symb_decoder(16#04#)) OR
 					(reg_q2449 AND symb_decoder(16#78#)) OR
 					(reg_q2449 AND symb_decoder(16#58#)) OR
 					(reg_q2449 AND symb_decoder(16#54#)) OR
 					(reg_q2449 AND symb_decoder(16#b2#)) OR
 					(reg_q2449 AND symb_decoder(16#9e#)) OR
 					(reg_q2449 AND symb_decoder(16#50#)) OR
 					(reg_q2449 AND symb_decoder(16#84#)) OR
 					(reg_q2449 AND symb_decoder(16#4e#)) OR
 					(reg_q2449 AND symb_decoder(16#ea#)) OR
 					(reg_q2449 AND symb_decoder(16#e0#)) OR
 					(reg_q2449 AND symb_decoder(16#f6#)) OR
 					(reg_q2449 AND symb_decoder(16#2e#)) OR
 					(reg_q2449 AND symb_decoder(16#e4#)) OR
 					(reg_q2449 AND symb_decoder(16#5c#)) OR
 					(reg_q2449 AND symb_decoder(16#7b#)) OR
 					(reg_q2449 AND symb_decoder(16#72#)) OR
 					(reg_q2449 AND symb_decoder(16#66#)) OR
 					(reg_q2449 AND symb_decoder(16#8b#)) OR
 					(reg_q2449 AND symb_decoder(16#15#)) OR
 					(reg_q2449 AND symb_decoder(16#ee#)) OR
 					(reg_q2449 AND symb_decoder(16#29#)) OR
 					(reg_q2449 AND symb_decoder(16#a0#)) OR
 					(reg_q2449 AND symb_decoder(16#5d#)) OR
 					(reg_q2449 AND symb_decoder(16#38#)) OR
 					(reg_q2449 AND symb_decoder(16#eb#)) OR
 					(reg_q2449 AND symb_decoder(16#b6#)) OR
 					(reg_q2449 AND symb_decoder(16#60#)) OR
 					(reg_q2449 AND symb_decoder(16#a6#)) OR
 					(reg_q2449 AND symb_decoder(16#2f#)) OR
 					(reg_q2449 AND symb_decoder(16#aa#)) OR
 					(reg_q2449 AND symb_decoder(16#75#)) OR
 					(reg_q2449 AND symb_decoder(16#1f#)) OR
 					(reg_q2449 AND symb_decoder(16#a1#)) OR
 					(reg_q2449 AND symb_decoder(16#85#)) OR
 					(reg_q2449 AND symb_decoder(16#ec#)) OR
 					(reg_q2449 AND symb_decoder(16#ab#)) OR
 					(reg_q2449 AND symb_decoder(16#25#)) OR
 					(reg_q2449 AND symb_decoder(16#cb#)) OR
 					(reg_q2449 AND symb_decoder(16#88#)) OR
 					(reg_q2449 AND symb_decoder(16#7c#)) OR
 					(reg_q2449 AND symb_decoder(16#2b#)) OR
 					(reg_q2449 AND symb_decoder(16#6b#)) OR
 					(reg_q2449 AND symb_decoder(16#a8#)) OR
 					(reg_q2449 AND symb_decoder(16#82#)) OR
 					(reg_q2449 AND symb_decoder(16#c4#)) OR
 					(reg_q2449 AND symb_decoder(16#87#)) OR
 					(reg_q2449 AND symb_decoder(16#16#)) OR
 					(reg_q2449 AND symb_decoder(16#c1#)) OR
 					(reg_q2449 AND symb_decoder(16#b3#)) OR
 					(reg_q2449 AND symb_decoder(16#3b#)) OR
 					(reg_q2449 AND symb_decoder(16#22#)) OR
 					(reg_q2449 AND symb_decoder(16#98#)) OR
 					(reg_q2449 AND symb_decoder(16#1a#)) OR
 					(reg_q2449 AND symb_decoder(16#a9#)) OR
 					(reg_q2449 AND symb_decoder(16#59#)) OR
 					(reg_q2449 AND symb_decoder(16#dd#)) OR
 					(reg_q2449 AND symb_decoder(16#d1#)) OR
 					(reg_q2449 AND symb_decoder(16#20#)) OR
 					(reg_q2449 AND symb_decoder(16#9a#)) OR
 					(reg_q2449 AND symb_decoder(16#c3#)) OR
 					(reg_q2449 AND symb_decoder(16#34#)) OR
 					(reg_q2449 AND symb_decoder(16#21#)) OR
 					(reg_q2449 AND symb_decoder(16#c9#)) OR
 					(reg_q2449 AND symb_decoder(16#a3#)) OR
 					(reg_q2449 AND symb_decoder(16#5a#)) OR
 					(reg_q2449 AND symb_decoder(16#28#)) OR
 					(reg_q2449 AND symb_decoder(16#f5#)) OR
 					(reg_q2449 AND symb_decoder(16#e8#)) OR
 					(reg_q2449 AND symb_decoder(16#bb#)) OR
 					(reg_q2449 AND symb_decoder(16#7e#)) OR
 					(reg_q2449 AND symb_decoder(16#b8#)) OR
 					(reg_q2449 AND symb_decoder(16#fe#)) OR
 					(reg_q2449 AND symb_decoder(16#df#)) OR
 					(reg_q2449 AND symb_decoder(16#8a#)) OR
 					(reg_q2449 AND symb_decoder(16#93#)) OR
 					(reg_q2449 AND symb_decoder(16#0d#)) OR
 					(reg_q2449 AND symb_decoder(16#6a#)) OR
 					(reg_q2449 AND symb_decoder(16#0e#)) OR
 					(reg_q2449 AND symb_decoder(16#09#)) OR
 					(reg_q2449 AND symb_decoder(16#36#)) OR
 					(reg_q2449 AND symb_decoder(16#8d#)) OR
 					(reg_q2449 AND symb_decoder(16#48#)) OR
 					(reg_q2449 AND symb_decoder(16#7a#)) OR
 					(reg_q2449 AND symb_decoder(16#39#)) OR
 					(reg_q2449 AND symb_decoder(16#e7#)) OR
 					(reg_q2449 AND symb_decoder(16#8c#)) OR
 					(reg_q2449 AND symb_decoder(16#02#)) OR
 					(reg_q2449 AND symb_decoder(16#ac#)) OR
 					(reg_q2449 AND symb_decoder(16#71#)) OR
 					(reg_q2449 AND symb_decoder(16#3f#)) OR
 					(reg_q2449 AND symb_decoder(16#73#)) OR
 					(reg_q2449 AND symb_decoder(16#c5#)) OR
 					(reg_q2449 AND symb_decoder(16#57#)) OR
 					(reg_q2449 AND symb_decoder(16#d6#)) OR
 					(reg_q2449 AND symb_decoder(16#6c#)) OR
 					(reg_q2449 AND symb_decoder(16#51#)) OR
 					(reg_q2449 AND symb_decoder(16#e6#)) OR
 					(reg_q2449 AND symb_decoder(16#7f#)) OR
 					(reg_q2449 AND symb_decoder(16#fb#)) OR
 					(reg_q2449 AND symb_decoder(16#56#)) OR
 					(reg_q2449 AND symb_decoder(16#ce#)) OR
 					(reg_q2449 AND symb_decoder(16#94#)) OR
 					(reg_q2449 AND symb_decoder(16#32#)) OR
 					(reg_q2449 AND symb_decoder(16#86#)) OR
 					(reg_q2449 AND symb_decoder(16#83#)) OR
 					(reg_q2449 AND symb_decoder(16#77#)) OR
 					(reg_q2449 AND symb_decoder(16#a4#)) OR
 					(reg_q2449 AND symb_decoder(16#6e#)) OR
 					(reg_q2449 AND symb_decoder(16#12#)) OR
 					(reg_q2449 AND symb_decoder(16#9f#)) OR
 					(reg_q2449 AND symb_decoder(16#3d#)) OR
 					(reg_q2449 AND symb_decoder(16#cd#)) OR
 					(reg_q2449 AND symb_decoder(16#44#)) OR
 					(reg_q2449 AND symb_decoder(16#68#)) OR
 					(reg_q2449 AND symb_decoder(16#b0#)) OR
 					(reg_q2449 AND symb_decoder(16#f9#)) OR
 					(reg_q2449 AND symb_decoder(16#5f#)) OR
 					(reg_q2449 AND symb_decoder(16#c7#)) OR
 					(reg_q2449 AND symb_decoder(16#74#)) OR
 					(reg_q2449 AND symb_decoder(16#af#)) OR
 					(reg_q2449 AND symb_decoder(16#d3#)) OR
 					(reg_q2449 AND symb_decoder(16#d4#)) OR
 					(reg_q2449 AND symb_decoder(16#80#)) OR
 					(reg_q2449 AND symb_decoder(16#e9#)) OR
 					(reg_q2449 AND symb_decoder(16#97#)) OR
 					(reg_q2449 AND symb_decoder(16#08#)) OR
 					(reg_q2449 AND symb_decoder(16#1e#)) OR
 					(reg_q2449 AND symb_decoder(16#65#)) OR
 					(reg_q2449 AND symb_decoder(16#43#)) OR
 					(reg_q2449 AND symb_decoder(16#2a#)) OR
 					(reg_q2449 AND symb_decoder(16#33#)) OR
 					(reg_q2449 AND symb_decoder(16#03#)) OR
 					(reg_q2449 AND symb_decoder(16#fc#));
reg_q2449_init <= '0' ;
	p_reg_q2449: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2449 <= reg_q2449_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2449 <= reg_q2449_init;
        else
          reg_q2449 <= reg_q2449_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q497_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q497 AND symb_decoder(16#20#)) OR
 					(reg_q497 AND symb_decoder(16#40#)) OR
 					(reg_q497 AND symb_decoder(16#8c#)) OR
 					(reg_q497 AND symb_decoder(16#9e#)) OR
 					(reg_q497 AND symb_decoder(16#9d#)) OR
 					(reg_q497 AND symb_decoder(16#af#)) OR
 					(reg_q497 AND symb_decoder(16#2e#)) OR
 					(reg_q497 AND symb_decoder(16#e9#)) OR
 					(reg_q497 AND symb_decoder(16#b4#)) OR
 					(reg_q497 AND symb_decoder(16#fe#)) OR
 					(reg_q497 AND symb_decoder(16#0b#)) OR
 					(reg_q497 AND symb_decoder(16#1d#)) OR
 					(reg_q497 AND symb_decoder(16#f2#)) OR
 					(reg_q497 AND symb_decoder(16#6a#)) OR
 					(reg_q497 AND symb_decoder(16#0d#)) OR
 					(reg_q497 AND symb_decoder(16#8f#)) OR
 					(reg_q497 AND symb_decoder(16#54#)) OR
 					(reg_q497 AND symb_decoder(16#73#)) OR
 					(reg_q497 AND symb_decoder(16#ec#)) OR
 					(reg_q497 AND symb_decoder(16#13#)) OR
 					(reg_q497 AND symb_decoder(16#12#)) OR
 					(reg_q497 AND symb_decoder(16#7a#)) OR
 					(reg_q497 AND symb_decoder(16#74#)) OR
 					(reg_q497 AND symb_decoder(16#4d#)) OR
 					(reg_q497 AND symb_decoder(16#57#)) OR
 					(reg_q497 AND symb_decoder(16#fc#)) OR
 					(reg_q497 AND symb_decoder(16#f1#)) OR
 					(reg_q497 AND symb_decoder(16#a8#)) OR
 					(reg_q497 AND symb_decoder(16#59#)) OR
 					(reg_q497 AND symb_decoder(16#a3#)) OR
 					(reg_q497 AND symb_decoder(16#23#)) OR
 					(reg_q497 AND symb_decoder(16#8b#)) OR
 					(reg_q497 AND symb_decoder(16#85#)) OR
 					(reg_q497 AND symb_decoder(16#53#)) OR
 					(reg_q497 AND symb_decoder(16#6b#)) OR
 					(reg_q497 AND symb_decoder(16#5f#)) OR
 					(reg_q497 AND symb_decoder(16#1c#)) OR
 					(reg_q497 AND symb_decoder(16#9f#)) OR
 					(reg_q497 AND symb_decoder(16#62#)) OR
 					(reg_q497 AND symb_decoder(16#58#)) OR
 					(reg_q497 AND symb_decoder(16#49#)) OR
 					(reg_q497 AND symb_decoder(16#c8#)) OR
 					(reg_q497 AND symb_decoder(16#c9#)) OR
 					(reg_q497 AND symb_decoder(16#03#)) OR
 					(reg_q497 AND symb_decoder(16#c4#)) OR
 					(reg_q497 AND symb_decoder(16#35#)) OR
 					(reg_q497 AND symb_decoder(16#dc#)) OR
 					(reg_q497 AND symb_decoder(16#88#)) OR
 					(reg_q497 AND symb_decoder(16#8d#)) OR
 					(reg_q497 AND symb_decoder(16#e5#)) OR
 					(reg_q497 AND symb_decoder(16#c2#)) OR
 					(reg_q497 AND symb_decoder(16#cd#)) OR
 					(reg_q497 AND symb_decoder(16#e8#)) OR
 					(reg_q497 AND symb_decoder(16#55#)) OR
 					(reg_q497 AND symb_decoder(16#fb#)) OR
 					(reg_q497 AND symb_decoder(16#7f#)) OR
 					(reg_q497 AND symb_decoder(16#45#)) OR
 					(reg_q497 AND symb_decoder(16#c7#)) OR
 					(reg_q497 AND symb_decoder(16#0a#)) OR
 					(reg_q497 AND symb_decoder(16#68#)) OR
 					(reg_q497 AND symb_decoder(16#5c#)) OR
 					(reg_q497 AND symb_decoder(16#ab#)) OR
 					(reg_q497 AND symb_decoder(16#91#)) OR
 					(reg_q497 AND symb_decoder(16#b1#)) OR
 					(reg_q497 AND symb_decoder(16#37#)) OR
 					(reg_q497 AND symb_decoder(16#a6#)) OR
 					(reg_q497 AND symb_decoder(16#ee#)) OR
 					(reg_q497 AND symb_decoder(16#94#)) OR
 					(reg_q497 AND symb_decoder(16#9b#)) OR
 					(reg_q497 AND symb_decoder(16#ae#)) OR
 					(reg_q497 AND symb_decoder(16#04#)) OR
 					(reg_q497 AND symb_decoder(16#66#)) OR
 					(reg_q497 AND symb_decoder(16#ce#)) OR
 					(reg_q497 AND symb_decoder(16#a9#)) OR
 					(reg_q497 AND symb_decoder(16#e0#)) OR
 					(reg_q497 AND symb_decoder(16#f0#)) OR
 					(reg_q497 AND symb_decoder(16#07#)) OR
 					(reg_q497 AND symb_decoder(16#ef#)) OR
 					(reg_q497 AND symb_decoder(16#d3#)) OR
 					(reg_q497 AND symb_decoder(16#eb#)) OR
 					(reg_q497 AND symb_decoder(16#bc#)) OR
 					(reg_q497 AND symb_decoder(16#38#)) OR
 					(reg_q497 AND symb_decoder(16#48#)) OR
 					(reg_q497 AND symb_decoder(16#51#)) OR
 					(reg_q497 AND symb_decoder(16#d0#)) OR
 					(reg_q497 AND symb_decoder(16#3e#)) OR
 					(reg_q497 AND symb_decoder(16#76#)) OR
 					(reg_q497 AND symb_decoder(16#5d#)) OR
 					(reg_q497 AND symb_decoder(16#be#)) OR
 					(reg_q497 AND symb_decoder(16#70#)) OR
 					(reg_q497 AND symb_decoder(16#6d#)) OR
 					(reg_q497 AND symb_decoder(16#21#)) OR
 					(reg_q497 AND symb_decoder(16#d4#)) OR
 					(reg_q497 AND symb_decoder(16#1f#)) OR
 					(reg_q497 AND symb_decoder(16#c5#)) OR
 					(reg_q497 AND symb_decoder(16#a4#)) OR
 					(reg_q497 AND symb_decoder(16#cb#)) OR
 					(reg_q497 AND symb_decoder(16#a7#)) OR
 					(reg_q497 AND symb_decoder(16#47#)) OR
 					(reg_q497 AND symb_decoder(16#b9#)) OR
 					(reg_q497 AND symb_decoder(16#69#)) OR
 					(reg_q497 AND symb_decoder(16#bf#)) OR
 					(reg_q497 AND symb_decoder(16#a0#)) OR
 					(reg_q497 AND symb_decoder(16#97#)) OR
 					(reg_q497 AND symb_decoder(16#02#)) OR
 					(reg_q497 AND symb_decoder(16#80#)) OR
 					(reg_q497 AND symb_decoder(16#33#)) OR
 					(reg_q497 AND symb_decoder(16#b0#)) OR
 					(reg_q497 AND symb_decoder(16#15#)) OR
 					(reg_q497 AND symb_decoder(16#3d#)) OR
 					(reg_q497 AND symb_decoder(16#4c#)) OR
 					(reg_q497 AND symb_decoder(16#46#)) OR
 					(reg_q497 AND symb_decoder(16#44#)) OR
 					(reg_q497 AND symb_decoder(16#79#)) OR
 					(reg_q497 AND symb_decoder(16#e7#)) OR
 					(reg_q497 AND symb_decoder(16#7d#)) OR
 					(reg_q497 AND symb_decoder(16#72#)) OR
 					(reg_q497 AND symb_decoder(16#78#)) OR
 					(reg_q497 AND symb_decoder(16#34#)) OR
 					(reg_q497 AND symb_decoder(16#29#)) OR
 					(reg_q497 AND symb_decoder(16#31#)) OR
 					(reg_q497 AND symb_decoder(16#c6#)) OR
 					(reg_q497 AND symb_decoder(16#c0#)) OR
 					(reg_q497 AND symb_decoder(16#9c#)) OR
 					(reg_q497 AND symb_decoder(16#d8#)) OR
 					(reg_q497 AND symb_decoder(16#50#)) OR
 					(reg_q497 AND symb_decoder(16#6c#)) OR
 					(reg_q497 AND symb_decoder(16#5b#)) OR
 					(reg_q497 AND symb_decoder(16#87#)) OR
 					(reg_q497 AND symb_decoder(16#8a#)) OR
 					(reg_q497 AND symb_decoder(16#4a#)) OR
 					(reg_q497 AND symb_decoder(16#d7#)) OR
 					(reg_q497 AND symb_decoder(16#96#)) OR
 					(reg_q497 AND symb_decoder(16#f5#)) OR
 					(reg_q497 AND symb_decoder(16#3c#)) OR
 					(reg_q497 AND symb_decoder(16#24#)) OR
 					(reg_q497 AND symb_decoder(16#bd#)) OR
 					(reg_q497 AND symb_decoder(16#32#)) OR
 					(reg_q497 AND symb_decoder(16#2a#)) OR
 					(reg_q497 AND symb_decoder(16#cf#)) OR
 					(reg_q497 AND symb_decoder(16#2b#)) OR
 					(reg_q497 AND symb_decoder(16#d9#)) OR
 					(reg_q497 AND symb_decoder(16#ff#)) OR
 					(reg_q497 AND symb_decoder(16#cc#)) OR
 					(reg_q497 AND symb_decoder(16#42#)) OR
 					(reg_q497 AND symb_decoder(16#a5#)) OR
 					(reg_q497 AND symb_decoder(16#86#)) OR
 					(reg_q497 AND symb_decoder(16#83#)) OR
 					(reg_q497 AND symb_decoder(16#b3#)) OR
 					(reg_q497 AND symb_decoder(16#92#)) OR
 					(reg_q497 AND symb_decoder(16#95#)) OR
 					(reg_q497 AND symb_decoder(16#aa#)) OR
 					(reg_q497 AND symb_decoder(16#fa#)) OR
 					(reg_q497 AND symb_decoder(16#6e#)) OR
 					(reg_q497 AND symb_decoder(16#82#)) OR
 					(reg_q497 AND symb_decoder(16#64#)) OR
 					(reg_q497 AND symb_decoder(16#22#)) OR
 					(reg_q497 AND symb_decoder(16#7b#)) OR
 					(reg_q497 AND symb_decoder(16#d6#)) OR
 					(reg_q497 AND symb_decoder(16#09#)) OR
 					(reg_q497 AND symb_decoder(16#ed#)) OR
 					(reg_q497 AND symb_decoder(16#4f#)) OR
 					(reg_q497 AND symb_decoder(16#a1#)) OR
 					(reg_q497 AND symb_decoder(16#c3#)) OR
 					(reg_q497 AND symb_decoder(16#28#)) OR
 					(reg_q497 AND symb_decoder(16#65#)) OR
 					(reg_q497 AND symb_decoder(16#5e#)) OR
 					(reg_q497 AND symb_decoder(16#63#)) OR
 					(reg_q497 AND symb_decoder(16#14#)) OR
 					(reg_q497 AND symb_decoder(16#1e#)) OR
 					(reg_q497 AND symb_decoder(16#71#)) OR
 					(reg_q497 AND symb_decoder(16#0e#)) OR
 					(reg_q497 AND symb_decoder(16#2d#)) OR
 					(reg_q497 AND symb_decoder(16#b6#)) OR
 					(reg_q497 AND symb_decoder(16#7c#)) OR
 					(reg_q497 AND symb_decoder(16#d1#)) OR
 					(reg_q497 AND symb_decoder(16#4b#)) OR
 					(reg_q497 AND symb_decoder(16#ca#)) OR
 					(reg_q497 AND symb_decoder(16#d2#)) OR
 					(reg_q497 AND symb_decoder(16#4e#)) OR
 					(reg_q497 AND symb_decoder(16#f4#)) OR
 					(reg_q497 AND symb_decoder(16#fd#)) OR
 					(reg_q497 AND symb_decoder(16#17#)) OR
 					(reg_q497 AND symb_decoder(16#bb#)) OR
 					(reg_q497 AND symb_decoder(16#25#)) OR
 					(reg_q497 AND symb_decoder(16#b8#)) OR
 					(reg_q497 AND symb_decoder(16#52#)) OR
 					(reg_q497 AND symb_decoder(16#e1#)) OR
 					(reg_q497 AND symb_decoder(16#90#)) OR
 					(reg_q497 AND symb_decoder(16#da#)) OR
 					(reg_q497 AND symb_decoder(16#27#)) OR
 					(reg_q497 AND symb_decoder(16#01#)) OR
 					(reg_q497 AND symb_decoder(16#9a#)) OR
 					(reg_q497 AND symb_decoder(16#b2#)) OR
 					(reg_q497 AND symb_decoder(16#89#)) OR
 					(reg_q497 AND symb_decoder(16#a2#)) OR
 					(reg_q497 AND symb_decoder(16#67#)) OR
 					(reg_q497 AND symb_decoder(16#5a#)) OR
 					(reg_q497 AND symb_decoder(16#39#)) OR
 					(reg_q497 AND symb_decoder(16#7e#)) OR
 					(reg_q497 AND symb_decoder(16#05#)) OR
 					(reg_q497 AND symb_decoder(16#dd#)) OR
 					(reg_q497 AND symb_decoder(16#36#)) OR
 					(reg_q497 AND symb_decoder(16#06#)) OR
 					(reg_q497 AND symb_decoder(16#1a#)) OR
 					(reg_q497 AND symb_decoder(16#df#)) OR
 					(reg_q497 AND symb_decoder(16#61#)) OR
 					(reg_q497 AND symb_decoder(16#81#)) OR
 					(reg_q497 AND symb_decoder(16#f9#)) OR
 					(reg_q497 AND symb_decoder(16#98#)) OR
 					(reg_q497 AND symb_decoder(16#30#)) OR
 					(reg_q497 AND symb_decoder(16#99#)) OR
 					(reg_q497 AND symb_decoder(16#00#)) OR
 					(reg_q497 AND symb_decoder(16#3b#)) OR
 					(reg_q497 AND symb_decoder(16#b7#)) OR
 					(reg_q497 AND symb_decoder(16#3f#)) OR
 					(reg_q497 AND symb_decoder(16#60#)) OR
 					(reg_q497 AND symb_decoder(16#1b#)) OR
 					(reg_q497 AND symb_decoder(16#93#)) OR
 					(reg_q497 AND symb_decoder(16#26#)) OR
 					(reg_q497 AND symb_decoder(16#f6#)) OR
 					(reg_q497 AND symb_decoder(16#e4#)) OR
 					(reg_q497 AND symb_decoder(16#ea#)) OR
 					(reg_q497 AND symb_decoder(16#08#)) OR
 					(reg_q497 AND symb_decoder(16#2f#)) OR
 					(reg_q497 AND symb_decoder(16#ba#)) OR
 					(reg_q497 AND symb_decoder(16#e3#)) OR
 					(reg_q497 AND symb_decoder(16#0f#)) OR
 					(reg_q497 AND symb_decoder(16#c1#)) OR
 					(reg_q497 AND symb_decoder(16#b5#)) OR
 					(reg_q497 AND symb_decoder(16#43#)) OR
 					(reg_q497 AND symb_decoder(16#ad#)) OR
 					(reg_q497 AND symb_decoder(16#0c#)) OR
 					(reg_q497 AND symb_decoder(16#e2#)) OR
 					(reg_q497 AND symb_decoder(16#75#)) OR
 					(reg_q497 AND symb_decoder(16#16#)) OR
 					(reg_q497 AND symb_decoder(16#84#)) OR
 					(reg_q497 AND symb_decoder(16#11#)) OR
 					(reg_q497 AND symb_decoder(16#2c#)) OR
 					(reg_q497 AND symb_decoder(16#19#)) OR
 					(reg_q497 AND symb_decoder(16#6f#)) OR
 					(reg_q497 AND symb_decoder(16#de#)) OR
 					(reg_q497 AND symb_decoder(16#41#)) OR
 					(reg_q497 AND symb_decoder(16#8e#)) OR
 					(reg_q497 AND symb_decoder(16#ac#)) OR
 					(reg_q497 AND symb_decoder(16#f7#)) OR
 					(reg_q497 AND symb_decoder(16#77#)) OR
 					(reg_q497 AND symb_decoder(16#e6#)) OR
 					(reg_q497 AND symb_decoder(16#f3#)) OR
 					(reg_q497 AND symb_decoder(16#db#)) OR
 					(reg_q497 AND symb_decoder(16#f8#)) OR
 					(reg_q497 AND symb_decoder(16#3a#)) OR
 					(reg_q497 AND symb_decoder(16#18#)) OR
 					(reg_q497 AND symb_decoder(16#56#)) OR
 					(reg_q497 AND symb_decoder(16#10#)) OR
 					(reg_q497 AND symb_decoder(16#d5#));
reg_q497_init <= '0' ;
	p_reg_q497: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q497 <= reg_q497_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q497 <= reg_q497_init;
        else
          reg_q497 <= reg_q497_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q757_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q757 AND symb_decoder(16#b4#)) OR
 					(reg_q757 AND symb_decoder(16#cc#)) OR
 					(reg_q757 AND symb_decoder(16#8e#)) OR
 					(reg_q757 AND symb_decoder(16#53#)) OR
 					(reg_q757 AND symb_decoder(16#2f#)) OR
 					(reg_q757 AND symb_decoder(16#b9#)) OR
 					(reg_q757 AND symb_decoder(16#14#)) OR
 					(reg_q757 AND symb_decoder(16#86#)) OR
 					(reg_q757 AND symb_decoder(16#30#)) OR
 					(reg_q757 AND symb_decoder(16#7a#)) OR
 					(reg_q757 AND symb_decoder(16#a0#)) OR
 					(reg_q757 AND symb_decoder(16#5b#)) OR
 					(reg_q757 AND symb_decoder(16#07#)) OR
 					(reg_q757 AND symb_decoder(16#5d#)) OR
 					(reg_q757 AND symb_decoder(16#10#)) OR
 					(reg_q757 AND symb_decoder(16#47#)) OR
 					(reg_q757 AND symb_decoder(16#88#)) OR
 					(reg_q757 AND symb_decoder(16#73#)) OR
 					(reg_q757 AND symb_decoder(16#3f#)) OR
 					(reg_q757 AND symb_decoder(16#9e#)) OR
 					(reg_q757 AND symb_decoder(16#d9#)) OR
 					(reg_q757 AND symb_decoder(16#65#)) OR
 					(reg_q757 AND symb_decoder(16#b8#)) OR
 					(reg_q757 AND symb_decoder(16#8f#)) OR
 					(reg_q757 AND symb_decoder(16#ce#)) OR
 					(reg_q757 AND symb_decoder(16#e0#)) OR
 					(reg_q757 AND symb_decoder(16#87#)) OR
 					(reg_q757 AND symb_decoder(16#ba#)) OR
 					(reg_q757 AND symb_decoder(16#04#)) OR
 					(reg_q757 AND symb_decoder(16#e7#)) OR
 					(reg_q757 AND symb_decoder(16#ed#)) OR
 					(reg_q757 AND symb_decoder(16#c3#)) OR
 					(reg_q757 AND symb_decoder(16#6b#)) OR
 					(reg_q757 AND symb_decoder(16#1e#)) OR
 					(reg_q757 AND symb_decoder(16#f9#)) OR
 					(reg_q757 AND symb_decoder(16#8a#)) OR
 					(reg_q757 AND symb_decoder(16#f4#)) OR
 					(reg_q757 AND symb_decoder(16#70#)) OR
 					(reg_q757 AND symb_decoder(16#90#)) OR
 					(reg_q757 AND symb_decoder(16#ec#)) OR
 					(reg_q757 AND symb_decoder(16#c0#)) OR
 					(reg_q757 AND symb_decoder(16#d4#)) OR
 					(reg_q757 AND symb_decoder(16#0a#)) OR
 					(reg_q757 AND symb_decoder(16#59#)) OR
 					(reg_q757 AND symb_decoder(16#e8#)) OR
 					(reg_q757 AND symb_decoder(16#6d#)) OR
 					(reg_q757 AND symb_decoder(16#e2#)) OR
 					(reg_q757 AND symb_decoder(16#08#)) OR
 					(reg_q757 AND symb_decoder(16#8c#)) OR
 					(reg_q757 AND symb_decoder(16#7d#)) OR
 					(reg_q757 AND symb_decoder(16#3a#)) OR
 					(reg_q757 AND symb_decoder(16#d6#)) OR
 					(reg_q757 AND symb_decoder(16#28#)) OR
 					(reg_q757 AND symb_decoder(16#7b#)) OR
 					(reg_q757 AND symb_decoder(16#0e#)) OR
 					(reg_q757 AND symb_decoder(16#f8#)) OR
 					(reg_q757 AND symb_decoder(16#bd#)) OR
 					(reg_q757 AND symb_decoder(16#24#)) OR
 					(reg_q757 AND symb_decoder(16#e9#)) OR
 					(reg_q757 AND symb_decoder(16#02#)) OR
 					(reg_q757 AND symb_decoder(16#80#)) OR
 					(reg_q757 AND symb_decoder(16#df#)) OR
 					(reg_q757 AND symb_decoder(16#18#)) OR
 					(reg_q757 AND symb_decoder(16#f2#)) OR
 					(reg_q757 AND symb_decoder(16#97#)) OR
 					(reg_q757 AND symb_decoder(16#05#)) OR
 					(reg_q757 AND symb_decoder(16#bf#)) OR
 					(reg_q757 AND symb_decoder(16#4b#)) OR
 					(reg_q757 AND symb_decoder(16#a3#)) OR
 					(reg_q757 AND symb_decoder(16#29#)) OR
 					(reg_q757 AND symb_decoder(16#a5#)) OR
 					(reg_q757 AND symb_decoder(16#fb#)) OR
 					(reg_q757 AND symb_decoder(16#f0#)) OR
 					(reg_q757 AND symb_decoder(16#49#)) OR
 					(reg_q757 AND symb_decoder(16#d0#)) OR
 					(reg_q757 AND symb_decoder(16#0c#)) OR
 					(reg_q757 AND symb_decoder(16#46#)) OR
 					(reg_q757 AND symb_decoder(16#8d#)) OR
 					(reg_q757 AND symb_decoder(16#be#)) OR
 					(reg_q757 AND symb_decoder(16#fd#)) OR
 					(reg_q757 AND symb_decoder(16#d1#)) OR
 					(reg_q757 AND symb_decoder(16#f5#)) OR
 					(reg_q757 AND symb_decoder(16#c9#)) OR
 					(reg_q757 AND symb_decoder(16#a4#)) OR
 					(reg_q757 AND symb_decoder(16#a7#)) OR
 					(reg_q757 AND symb_decoder(16#1c#)) OR
 					(reg_q757 AND symb_decoder(16#45#)) OR
 					(reg_q757 AND symb_decoder(16#21#)) OR
 					(reg_q757 AND symb_decoder(16#01#)) OR
 					(reg_q757 AND symb_decoder(16#b2#)) OR
 					(reg_q757 AND symb_decoder(16#58#)) OR
 					(reg_q757 AND symb_decoder(16#2c#)) OR
 					(reg_q757 AND symb_decoder(16#f1#)) OR
 					(reg_q757 AND symb_decoder(16#61#)) OR
 					(reg_q757 AND symb_decoder(16#12#)) OR
 					(reg_q757 AND symb_decoder(16#6c#)) OR
 					(reg_q757 AND symb_decoder(16#e6#)) OR
 					(reg_q757 AND symb_decoder(16#ee#)) OR
 					(reg_q757 AND symb_decoder(16#1d#)) OR
 					(reg_q757 AND symb_decoder(16#ac#)) OR
 					(reg_q757 AND symb_decoder(16#c5#)) OR
 					(reg_q757 AND symb_decoder(16#5e#)) OR
 					(reg_q757 AND symb_decoder(16#d8#)) OR
 					(reg_q757 AND symb_decoder(16#a8#)) OR
 					(reg_q757 AND symb_decoder(16#2e#)) OR
 					(reg_q757 AND symb_decoder(16#93#)) OR
 					(reg_q757 AND symb_decoder(16#7e#)) OR
 					(reg_q757 AND symb_decoder(16#23#)) OR
 					(reg_q757 AND symb_decoder(16#8b#)) OR
 					(reg_q757 AND symb_decoder(16#44#)) OR
 					(reg_q757 AND symb_decoder(16#0d#)) OR
 					(reg_q757 AND symb_decoder(16#9a#)) OR
 					(reg_q757 AND symb_decoder(16#d2#)) OR
 					(reg_q757 AND symb_decoder(16#85#)) OR
 					(reg_q757 AND symb_decoder(16#09#)) OR
 					(reg_q757 AND symb_decoder(16#d7#)) OR
 					(reg_q757 AND symb_decoder(16#de#)) OR
 					(reg_q757 AND symb_decoder(16#99#)) OR
 					(reg_q757 AND symb_decoder(16#62#)) OR
 					(reg_q757 AND symb_decoder(16#4e#)) OR
 					(reg_q757 AND symb_decoder(16#94#)) OR
 					(reg_q757 AND symb_decoder(16#22#)) OR
 					(reg_q757 AND symb_decoder(16#43#)) OR
 					(reg_q757 AND symb_decoder(16#eb#)) OR
 					(reg_q757 AND symb_decoder(16#3b#)) OR
 					(reg_q757 AND symb_decoder(16#76#)) OR
 					(reg_q757 AND symb_decoder(16#f7#)) OR
 					(reg_q757 AND symb_decoder(16#da#)) OR
 					(reg_q757 AND symb_decoder(16#6e#)) OR
 					(reg_q757 AND symb_decoder(16#71#)) OR
 					(reg_q757 AND symb_decoder(16#c4#)) OR
 					(reg_q757 AND symb_decoder(16#cb#)) OR
 					(reg_q757 AND symb_decoder(16#13#)) OR
 					(reg_q757 AND symb_decoder(16#31#)) OR
 					(reg_q757 AND symb_decoder(16#48#)) OR
 					(reg_q757 AND symb_decoder(16#11#)) OR
 					(reg_q757 AND symb_decoder(16#72#)) OR
 					(reg_q757 AND symb_decoder(16#75#)) OR
 					(reg_q757 AND symb_decoder(16#2d#)) OR
 					(reg_q757 AND symb_decoder(16#42#)) OR
 					(reg_q757 AND symb_decoder(16#41#)) OR
 					(reg_q757 AND symb_decoder(16#af#)) OR
 					(reg_q757 AND symb_decoder(16#3d#)) OR
 					(reg_q757 AND symb_decoder(16#fe#)) OR
 					(reg_q757 AND symb_decoder(16#17#)) OR
 					(reg_q757 AND symb_decoder(16#ea#)) OR
 					(reg_q757 AND symb_decoder(16#dc#)) OR
 					(reg_q757 AND symb_decoder(16#f6#)) OR
 					(reg_q757 AND symb_decoder(16#db#)) OR
 					(reg_q757 AND symb_decoder(16#15#)) OR
 					(reg_q757 AND symb_decoder(16#64#)) OR
 					(reg_q757 AND symb_decoder(16#d3#)) OR
 					(reg_q757 AND symb_decoder(16#4a#)) OR
 					(reg_q757 AND symb_decoder(16#60#)) OR
 					(reg_q757 AND symb_decoder(16#83#)) OR
 					(reg_q757 AND symb_decoder(16#cf#)) OR
 					(reg_q757 AND symb_decoder(16#6a#)) OR
 					(reg_q757 AND symb_decoder(16#9c#)) OR
 					(reg_q757 AND symb_decoder(16#9d#)) OR
 					(reg_q757 AND symb_decoder(16#03#)) OR
 					(reg_q757 AND symb_decoder(16#92#)) OR
 					(reg_q757 AND symb_decoder(16#9b#)) OR
 					(reg_q757 AND symb_decoder(16#67#)) OR
 					(reg_q757 AND symb_decoder(16#1b#)) OR
 					(reg_q757 AND symb_decoder(16#bb#)) OR
 					(reg_q757 AND symb_decoder(16#b0#)) OR
 					(reg_q757 AND symb_decoder(16#aa#)) OR
 					(reg_q757 AND symb_decoder(16#2b#)) OR
 					(reg_q757 AND symb_decoder(16#d5#)) OR
 					(reg_q757 AND symb_decoder(16#b6#)) OR
 					(reg_q757 AND symb_decoder(16#ae#)) OR
 					(reg_q757 AND symb_decoder(16#89#)) OR
 					(reg_q757 AND symb_decoder(16#c8#)) OR
 					(reg_q757 AND symb_decoder(16#ca#)) OR
 					(reg_q757 AND symb_decoder(16#3e#)) OR
 					(reg_q757 AND symb_decoder(16#79#)) OR
 					(reg_q757 AND symb_decoder(16#2a#)) OR
 					(reg_q757 AND symb_decoder(16#a9#)) OR
 					(reg_q757 AND symb_decoder(16#16#)) OR
 					(reg_q757 AND symb_decoder(16#56#)) OR
 					(reg_q757 AND symb_decoder(16#c2#)) OR
 					(reg_q757 AND symb_decoder(16#37#)) OR
 					(reg_q757 AND symb_decoder(16#66#)) OR
 					(reg_q757 AND symb_decoder(16#33#)) OR
 					(reg_q757 AND symb_decoder(16#57#)) OR
 					(reg_q757 AND symb_decoder(16#4f#)) OR
 					(reg_q757 AND symb_decoder(16#e1#)) OR
 					(reg_q757 AND symb_decoder(16#91#)) OR
 					(reg_q757 AND symb_decoder(16#f3#)) OR
 					(reg_q757 AND symb_decoder(16#39#)) OR
 					(reg_q757 AND symb_decoder(16#00#)) OR
 					(reg_q757 AND symb_decoder(16#4d#)) OR
 					(reg_q757 AND symb_decoder(16#84#)) OR
 					(reg_q757 AND symb_decoder(16#82#)) OR
 					(reg_q757 AND symb_decoder(16#34#)) OR
 					(reg_q757 AND symb_decoder(16#b3#)) OR
 					(reg_q757 AND symb_decoder(16#ef#)) OR
 					(reg_q757 AND symb_decoder(16#50#)) OR
 					(reg_q757 AND symb_decoder(16#55#)) OR
 					(reg_q757 AND symb_decoder(16#74#)) OR
 					(reg_q757 AND symb_decoder(16#54#)) OR
 					(reg_q757 AND symb_decoder(16#77#)) OR
 					(reg_q757 AND symb_decoder(16#9f#)) OR
 					(reg_q757 AND symb_decoder(16#51#)) OR
 					(reg_q757 AND symb_decoder(16#4c#)) OR
 					(reg_q757 AND symb_decoder(16#0b#)) OR
 					(reg_q757 AND symb_decoder(16#63#)) OR
 					(reg_q757 AND symb_decoder(16#20#)) OR
 					(reg_q757 AND symb_decoder(16#a1#)) OR
 					(reg_q757 AND symb_decoder(16#35#)) OR
 					(reg_q757 AND symb_decoder(16#81#)) OR
 					(reg_q757 AND symb_decoder(16#19#)) OR
 					(reg_q757 AND symb_decoder(16#b5#)) OR
 					(reg_q757 AND symb_decoder(16#1f#)) OR
 					(reg_q757 AND symb_decoder(16#6f#)) OR
 					(reg_q757 AND symb_decoder(16#5f#)) OR
 					(reg_q757 AND symb_decoder(16#98#)) OR
 					(reg_q757 AND symb_decoder(16#25#)) OR
 					(reg_q757 AND symb_decoder(16#fc#)) OR
 					(reg_q757 AND symb_decoder(16#ab#)) OR
 					(reg_q757 AND symb_decoder(16#b1#)) OR
 					(reg_q757 AND symb_decoder(16#69#)) OR
 					(reg_q757 AND symb_decoder(16#7f#)) OR
 					(reg_q757 AND symb_decoder(16#36#)) OR
 					(reg_q757 AND symb_decoder(16#a2#)) OR
 					(reg_q757 AND symb_decoder(16#0f#)) OR
 					(reg_q757 AND symb_decoder(16#27#)) OR
 					(reg_q757 AND symb_decoder(16#cd#)) OR
 					(reg_q757 AND symb_decoder(16#68#)) OR
 					(reg_q757 AND symb_decoder(16#bc#)) OR
 					(reg_q757 AND symb_decoder(16#26#)) OR
 					(reg_q757 AND symb_decoder(16#06#)) OR
 					(reg_q757 AND symb_decoder(16#e5#)) OR
 					(reg_q757 AND symb_decoder(16#dd#)) OR
 					(reg_q757 AND symb_decoder(16#78#)) OR
 					(reg_q757 AND symb_decoder(16#52#)) OR
 					(reg_q757 AND symb_decoder(16#96#)) OR
 					(reg_q757 AND symb_decoder(16#ff#)) OR
 					(reg_q757 AND symb_decoder(16#95#)) OR
 					(reg_q757 AND symb_decoder(16#c6#)) OR
 					(reg_q757 AND symb_decoder(16#5a#)) OR
 					(reg_q757 AND symb_decoder(16#1a#)) OR
 					(reg_q757 AND symb_decoder(16#40#)) OR
 					(reg_q757 AND symb_decoder(16#fa#)) OR
 					(reg_q757 AND symb_decoder(16#c7#)) OR
 					(reg_q757 AND symb_decoder(16#3c#)) OR
 					(reg_q757 AND symb_decoder(16#c1#)) OR
 					(reg_q757 AND symb_decoder(16#ad#)) OR
 					(reg_q757 AND symb_decoder(16#a6#)) OR
 					(reg_q757 AND symb_decoder(16#5c#)) OR
 					(reg_q757 AND symb_decoder(16#38#)) OR
 					(reg_q757 AND symb_decoder(16#7c#)) OR
 					(reg_q757 AND symb_decoder(16#e3#)) OR
 					(reg_q757 AND symb_decoder(16#32#)) OR
 					(reg_q757 AND symb_decoder(16#e4#)) OR
 					(reg_q757 AND symb_decoder(16#b7#));
reg_q757_init <= '0' ;
	p_reg_q757: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q757 <= reg_q757_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q757 <= reg_q757_init;
        else
          reg_q757 <= reg_q757_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph28

reg_q1626_in <= (reg_q1626 AND symb_decoder(16#fc#)) OR
 					(reg_q1626 AND symb_decoder(16#9d#)) OR
 					(reg_q1626 AND symb_decoder(16#75#)) OR
 					(reg_q1626 AND symb_decoder(16#d2#)) OR
 					(reg_q1626 AND symb_decoder(16#31#)) OR
 					(reg_q1626 AND symb_decoder(16#1b#)) OR
 					(reg_q1626 AND symb_decoder(16#78#)) OR
 					(reg_q1626 AND symb_decoder(16#e0#)) OR
 					(reg_q1626 AND symb_decoder(16#50#)) OR
 					(reg_q1626 AND symb_decoder(16#10#)) OR
 					(reg_q1626 AND symb_decoder(16#83#)) OR
 					(reg_q1626 AND symb_decoder(16#18#)) OR
 					(reg_q1626 AND symb_decoder(16#b3#)) OR
 					(reg_q1626 AND symb_decoder(16#c1#)) OR
 					(reg_q1626 AND symb_decoder(16#2d#)) OR
 					(reg_q1626 AND symb_decoder(16#99#)) OR
 					(reg_q1626 AND symb_decoder(16#b0#)) OR
 					(reg_q1626 AND symb_decoder(16#26#)) OR
 					(reg_q1626 AND symb_decoder(16#69#)) OR
 					(reg_q1626 AND symb_decoder(16#0b#)) OR
 					(reg_q1626 AND symb_decoder(16#b9#)) OR
 					(reg_q1626 AND symb_decoder(16#ab#)) OR
 					(reg_q1626 AND symb_decoder(16#7a#)) OR
 					(reg_q1626 AND symb_decoder(16#52#)) OR
 					(reg_q1626 AND symb_decoder(16#91#)) OR
 					(reg_q1626 AND symb_decoder(16#45#)) OR
 					(reg_q1626 AND symb_decoder(16#d7#)) OR
 					(reg_q1626 AND symb_decoder(16#a2#)) OR
 					(reg_q1626 AND symb_decoder(16#cb#)) OR
 					(reg_q1626 AND symb_decoder(16#5e#)) OR
 					(reg_q1626 AND symb_decoder(16#ce#)) OR
 					(reg_q1626 AND symb_decoder(16#c5#)) OR
 					(reg_q1626 AND symb_decoder(16#bd#)) OR
 					(reg_q1626 AND symb_decoder(16#20#)) OR
 					(reg_q1626 AND symb_decoder(16#04#)) OR
 					(reg_q1626 AND symb_decoder(16#ca#)) OR
 					(reg_q1626 AND symb_decoder(16#94#)) OR
 					(reg_q1626 AND symb_decoder(16#a4#)) OR
 					(reg_q1626 AND symb_decoder(16#a1#)) OR
 					(reg_q1626 AND symb_decoder(16#39#)) OR
 					(reg_q1626 AND symb_decoder(16#fa#)) OR
 					(reg_q1626 AND symb_decoder(16#13#)) OR
 					(reg_q1626 AND symb_decoder(16#ae#)) OR
 					(reg_q1626 AND symb_decoder(16#ec#)) OR
 					(reg_q1626 AND symb_decoder(16#02#)) OR
 					(reg_q1626 AND symb_decoder(16#de#)) OR
 					(reg_q1626 AND symb_decoder(16#58#)) OR
 					(reg_q1626 AND symb_decoder(16#f6#)) OR
 					(reg_q1626 AND symb_decoder(16#79#)) OR
 					(reg_q1626 AND symb_decoder(16#e1#)) OR
 					(reg_q1626 AND symb_decoder(16#d1#)) OR
 					(reg_q1626 AND symb_decoder(16#22#)) OR
 					(reg_q1626 AND symb_decoder(16#5b#)) OR
 					(reg_q1626 AND symb_decoder(16#09#)) OR
 					(reg_q1626 AND symb_decoder(16#8d#)) OR
 					(reg_q1626 AND symb_decoder(16#f7#)) OR
 					(reg_q1626 AND symb_decoder(16#15#)) OR
 					(reg_q1626 AND symb_decoder(16#ed#)) OR
 					(reg_q1626 AND symb_decoder(16#96#)) OR
 					(reg_q1626 AND symb_decoder(16#1e#)) OR
 					(reg_q1626 AND symb_decoder(16#f3#)) OR
 					(reg_q1626 AND symb_decoder(16#84#)) OR
 					(reg_q1626 AND symb_decoder(16#7b#)) OR
 					(reg_q1626 AND symb_decoder(16#70#)) OR
 					(reg_q1626 AND symb_decoder(16#5c#)) OR
 					(reg_q1626 AND symb_decoder(16#6a#)) OR
 					(reg_q1626 AND symb_decoder(16#cc#)) OR
 					(reg_q1626 AND symb_decoder(16#b5#)) OR
 					(reg_q1626 AND symb_decoder(16#88#)) OR
 					(reg_q1626 AND symb_decoder(16#81#)) OR
 					(reg_q1626 AND symb_decoder(16#f0#)) OR
 					(reg_q1626 AND symb_decoder(16#c8#)) OR
 					(reg_q1626 AND symb_decoder(16#fd#)) OR
 					(reg_q1626 AND symb_decoder(16#66#)) OR
 					(reg_q1626 AND symb_decoder(16#08#)) OR
 					(reg_q1626 AND symb_decoder(16#0c#)) OR
 					(reg_q1626 AND symb_decoder(16#ff#)) OR
 					(reg_q1626 AND symb_decoder(16#b2#)) OR
 					(reg_q1626 AND symb_decoder(16#4e#)) OR
 					(reg_q1626 AND symb_decoder(16#ea#)) OR
 					(reg_q1626 AND symb_decoder(16#b6#)) OR
 					(reg_q1626 AND symb_decoder(16#b4#)) OR
 					(reg_q1626 AND symb_decoder(16#ac#)) OR
 					(reg_q1626 AND symb_decoder(16#54#)) OR
 					(reg_q1626 AND symb_decoder(16#d9#)) OR
 					(reg_q1626 AND symb_decoder(16#3b#)) OR
 					(reg_q1626 AND symb_decoder(16#1d#)) OR
 					(reg_q1626 AND symb_decoder(16#63#)) OR
 					(reg_q1626 AND symb_decoder(16#3a#)) OR
 					(reg_q1626 AND symb_decoder(16#bb#)) OR
 					(reg_q1626 AND symb_decoder(16#36#)) OR
 					(reg_q1626 AND symb_decoder(16#7c#)) OR
 					(reg_q1626 AND symb_decoder(16#74#)) OR
 					(reg_q1626 AND symb_decoder(16#77#)) OR
 					(reg_q1626 AND symb_decoder(16#30#)) OR
 					(reg_q1626 AND symb_decoder(16#ef#)) OR
 					(reg_q1626 AND symb_decoder(16#53#)) OR
 					(reg_q1626 AND symb_decoder(16#ee#)) OR
 					(reg_q1626 AND symb_decoder(16#64#)) OR
 					(reg_q1626 AND symb_decoder(16#e5#)) OR
 					(reg_q1626 AND symb_decoder(16#23#)) OR
 					(reg_q1626 AND symb_decoder(16#06#)) OR
 					(reg_q1626 AND symb_decoder(16#4a#)) OR
 					(reg_q1626 AND symb_decoder(16#dc#)) OR
 					(reg_q1626 AND symb_decoder(16#c9#)) OR
 					(reg_q1626 AND symb_decoder(16#da#)) OR
 					(reg_q1626 AND symb_decoder(16#12#)) OR
 					(reg_q1626 AND symb_decoder(16#72#)) OR
 					(reg_q1626 AND symb_decoder(16#9b#)) OR
 					(reg_q1626 AND symb_decoder(16#29#)) OR
 					(reg_q1626 AND symb_decoder(16#cf#)) OR
 					(reg_q1626 AND symb_decoder(16#44#)) OR
 					(reg_q1626 AND symb_decoder(16#fe#)) OR
 					(reg_q1626 AND symb_decoder(16#93#)) OR
 					(reg_q1626 AND symb_decoder(16#8a#)) OR
 					(reg_q1626 AND symb_decoder(16#a7#)) OR
 					(reg_q1626 AND symb_decoder(16#e4#)) OR
 					(reg_q1626 AND symb_decoder(16#6c#)) OR
 					(reg_q1626 AND symb_decoder(16#f9#)) OR
 					(reg_q1626 AND symb_decoder(16#4c#)) OR
 					(reg_q1626 AND symb_decoder(16#98#)) OR
 					(reg_q1626 AND symb_decoder(16#2b#)) OR
 					(reg_q1626 AND symb_decoder(16#3d#)) OR
 					(reg_q1626 AND symb_decoder(16#f8#)) OR
 					(reg_q1626 AND symb_decoder(16#1a#)) OR
 					(reg_q1626 AND symb_decoder(16#57#)) OR
 					(reg_q1626 AND symb_decoder(16#17#)) OR
 					(reg_q1626 AND symb_decoder(16#d8#)) OR
 					(reg_q1626 AND symb_decoder(16#40#)) OR
 					(reg_q1626 AND symb_decoder(16#82#)) OR
 					(reg_q1626 AND symb_decoder(16#f5#)) OR
 					(reg_q1626 AND symb_decoder(16#85#)) OR
 					(reg_q1626 AND symb_decoder(16#9c#)) OR
 					(reg_q1626 AND symb_decoder(16#bc#)) OR
 					(reg_q1626 AND symb_decoder(16#a9#)) OR
 					(reg_q1626 AND symb_decoder(16#e6#)) OR
 					(reg_q1626 AND symb_decoder(16#eb#)) OR
 					(reg_q1626 AND symb_decoder(16#aa#)) OR
 					(reg_q1626 AND symb_decoder(16#8b#)) OR
 					(reg_q1626 AND symb_decoder(16#7d#)) OR
 					(reg_q1626 AND symb_decoder(16#90#)) OR
 					(reg_q1626 AND symb_decoder(16#48#)) OR
 					(reg_q1626 AND symb_decoder(16#fb#)) OR
 					(reg_q1626 AND symb_decoder(16#a0#)) OR
 					(reg_q1626 AND symb_decoder(16#b7#)) OR
 					(reg_q1626 AND symb_decoder(16#d4#)) OR
 					(reg_q1626 AND symb_decoder(16#80#)) OR
 					(reg_q1626 AND symb_decoder(16#34#)) OR
 					(reg_q1626 AND symb_decoder(16#56#)) OR
 					(reg_q1626 AND symb_decoder(16#35#)) OR
 					(reg_q1626 AND symb_decoder(16#60#)) OR
 					(reg_q1626 AND symb_decoder(16#6b#)) OR
 					(reg_q1626 AND symb_decoder(16#e2#)) OR
 					(reg_q1626 AND symb_decoder(16#89#)) OR
 					(reg_q1626 AND symb_decoder(16#38#)) OR
 					(reg_q1626 AND symb_decoder(16#59#)) OR
 					(reg_q1626 AND symb_decoder(16#27#)) OR
 					(reg_q1626 AND symb_decoder(16#71#)) OR
 					(reg_q1626 AND symb_decoder(16#97#)) OR
 					(reg_q1626 AND symb_decoder(16#9f#)) OR
 					(reg_q1626 AND symb_decoder(16#76#)) OR
 					(reg_q1626 AND symb_decoder(16#41#)) OR
 					(reg_q1626 AND symb_decoder(16#d3#)) OR
 					(reg_q1626 AND symb_decoder(16#d5#)) OR
 					(reg_q1626 AND symb_decoder(16#3f#)) OR
 					(reg_q1626 AND symb_decoder(16#67#)) OR
 					(reg_q1626 AND symb_decoder(16#f1#)) OR
 					(reg_q1626 AND symb_decoder(16#c4#)) OR
 					(reg_q1626 AND symb_decoder(16#df#)) OR
 					(reg_q1626 AND symb_decoder(16#db#)) OR
 					(reg_q1626 AND symb_decoder(16#61#)) OR
 					(reg_q1626 AND symb_decoder(16#0e#)) OR
 					(reg_q1626 AND symb_decoder(16#42#)) OR
 					(reg_q1626 AND symb_decoder(16#62#)) OR
 					(reg_q1626 AND symb_decoder(16#4d#)) OR
 					(reg_q1626 AND symb_decoder(16#be#)) OR
 					(reg_q1626 AND symb_decoder(16#c3#)) OR
 					(reg_q1626 AND symb_decoder(16#2e#)) OR
 					(reg_q1626 AND symb_decoder(16#a3#)) OR
 					(reg_q1626 AND symb_decoder(16#b8#)) OR
 					(reg_q1626 AND symb_decoder(16#05#)) OR
 					(reg_q1626 AND symb_decoder(16#2c#)) OR
 					(reg_q1626 AND symb_decoder(16#e3#)) OR
 					(reg_q1626 AND symb_decoder(16#37#)) OR
 					(reg_q1626 AND symb_decoder(16#2a#)) OR
 					(reg_q1626 AND symb_decoder(16#68#)) OR
 					(reg_q1626 AND symb_decoder(16#73#)) OR
 					(reg_q1626 AND symb_decoder(16#af#)) OR
 					(reg_q1626 AND symb_decoder(16#c7#)) OR
 					(reg_q1626 AND symb_decoder(16#49#)) OR
 					(reg_q1626 AND symb_decoder(16#ad#)) OR
 					(reg_q1626 AND symb_decoder(16#5f#)) OR
 					(reg_q1626 AND symb_decoder(16#14#)) OR
 					(reg_q1626 AND symb_decoder(16#01#)) OR
 					(reg_q1626 AND symb_decoder(16#e8#)) OR
 					(reg_q1626 AND symb_decoder(16#00#)) OR
 					(reg_q1626 AND symb_decoder(16#43#)) OR
 					(reg_q1626 AND symb_decoder(16#0f#)) OR
 					(reg_q1626 AND symb_decoder(16#33#)) OR
 					(reg_q1626 AND symb_decoder(16#f2#)) OR
 					(reg_q1626 AND symb_decoder(16#9e#)) OR
 					(reg_q1626 AND symb_decoder(16#1f#)) OR
 					(reg_q1626 AND symb_decoder(16#92#)) OR
 					(reg_q1626 AND symb_decoder(16#7f#)) OR
 					(reg_q1626 AND symb_decoder(16#11#)) OR
 					(reg_q1626 AND symb_decoder(16#19#)) OR
 					(reg_q1626 AND symb_decoder(16#e9#)) OR
 					(reg_q1626 AND symb_decoder(16#8c#)) OR
 					(reg_q1626 AND symb_decoder(16#07#)) OR
 					(reg_q1626 AND symb_decoder(16#8f#)) OR
 					(reg_q1626 AND symb_decoder(16#dd#)) OR
 					(reg_q1626 AND symb_decoder(16#a5#)) OR
 					(reg_q1626 AND symb_decoder(16#03#)) OR
 					(reg_q1626 AND symb_decoder(16#3e#)) OR
 					(reg_q1626 AND symb_decoder(16#a6#)) OR
 					(reg_q1626 AND symb_decoder(16#2f#)) OR
 					(reg_q1626 AND symb_decoder(16#8e#)) OR
 					(reg_q1626 AND symb_decoder(16#bf#)) OR
 					(reg_q1626 AND symb_decoder(16#32#)) OR
 					(reg_q1626 AND symb_decoder(16#6f#)) OR
 					(reg_q1626 AND symb_decoder(16#28#)) OR
 					(reg_q1626 AND symb_decoder(16#5a#)) OR
 					(reg_q1626 AND symb_decoder(16#ba#)) OR
 					(reg_q1626 AND symb_decoder(16#9a#)) OR
 					(reg_q1626 AND symb_decoder(16#4f#)) OR
 					(reg_q1626 AND symb_decoder(16#c6#)) OR
 					(reg_q1626 AND symb_decoder(16#3c#)) OR
 					(reg_q1626 AND symb_decoder(16#d0#)) OR
 					(reg_q1626 AND symb_decoder(16#a8#)) OR
 					(reg_q1626 AND symb_decoder(16#55#)) OR
 					(reg_q1626 AND symb_decoder(16#47#)) OR
 					(reg_q1626 AND symb_decoder(16#f4#)) OR
 					(reg_q1626 AND symb_decoder(16#87#)) OR
 					(reg_q1626 AND symb_decoder(16#65#)) OR
 					(reg_q1626 AND symb_decoder(16#16#)) OR
 					(reg_q1626 AND symb_decoder(16#e7#)) OR
 					(reg_q1626 AND symb_decoder(16#46#)) OR
 					(reg_q1626 AND symb_decoder(16#cd#)) OR
 					(reg_q1626 AND symb_decoder(16#95#)) OR
 					(reg_q1626 AND symb_decoder(16#c2#)) OR
 					(reg_q1626 AND symb_decoder(16#d6#)) OR
 					(reg_q1626 AND symb_decoder(16#25#)) OR
 					(reg_q1626 AND symb_decoder(16#6e#)) OR
 					(reg_q1626 AND symb_decoder(16#6d#)) OR
 					(reg_q1626 AND symb_decoder(16#24#)) OR
 					(reg_q1626 AND symb_decoder(16#7e#)) OR
 					(reg_q1626 AND symb_decoder(16#21#)) OR
 					(reg_q1626 AND symb_decoder(16#86#)) OR
 					(reg_q1626 AND symb_decoder(16#1c#)) OR
 					(reg_q1626 AND symb_decoder(16#51#)) OR
 					(reg_q1626 AND symb_decoder(16#5d#)) OR
 					(reg_q1626 AND symb_decoder(16#4b#)) OR
 					(reg_q1626 AND symb_decoder(16#b1#)) OR
 					(reg_q1626 AND symb_decoder(16#c0#)) OR
 					(reg_q1616 AND symb_decoder(16#02#)) OR
 					(reg_q1616 AND symb_decoder(16#04#)) OR
 					(reg_q1616 AND symb_decoder(16#2c#)) OR
 					(reg_q1616 AND symb_decoder(16#ae#)) OR
 					(reg_q1616 AND symb_decoder(16#83#)) OR
 					(reg_q1616 AND symb_decoder(16#a6#)) OR
 					(reg_q1616 AND symb_decoder(16#74#)) OR
 					(reg_q1616 AND symb_decoder(16#72#)) OR
 					(reg_q1616 AND symb_decoder(16#fa#)) OR
 					(reg_q1616 AND symb_decoder(16#1a#)) OR
 					(reg_q1616 AND symb_decoder(16#42#)) OR
 					(reg_q1616 AND symb_decoder(16#a0#)) OR
 					(reg_q1616 AND symb_decoder(16#24#)) OR
 					(reg_q1616 AND symb_decoder(16#af#)) OR
 					(reg_q1616 AND symb_decoder(16#ec#)) OR
 					(reg_q1616 AND symb_decoder(16#1d#)) OR
 					(reg_q1616 AND symb_decoder(16#2b#)) OR
 					(reg_q1616 AND symb_decoder(16#14#)) OR
 					(reg_q1616 AND symb_decoder(16#d4#)) OR
 					(reg_q1616 AND symb_decoder(16#e7#)) OR
 					(reg_q1616 AND symb_decoder(16#82#)) OR
 					(reg_q1616 AND symb_decoder(16#cb#)) OR
 					(reg_q1616 AND symb_decoder(16#92#)) OR
 					(reg_q1616 AND symb_decoder(16#80#)) OR
 					(reg_q1616 AND symb_decoder(16#cf#)) OR
 					(reg_q1616 AND symb_decoder(16#e4#)) OR
 					(reg_q1616 AND symb_decoder(16#44#)) OR
 					(reg_q1616 AND symb_decoder(16#11#)) OR
 					(reg_q1616 AND symb_decoder(16#b9#)) OR
 					(reg_q1616 AND symb_decoder(16#19#)) OR
 					(reg_q1616 AND symb_decoder(16#d5#)) OR
 					(reg_q1616 AND symb_decoder(16#3d#)) OR
 					(reg_q1616 AND symb_decoder(16#79#)) OR
 					(reg_q1616 AND symb_decoder(16#0c#)) OR
 					(reg_q1616 AND symb_decoder(16#0f#)) OR
 					(reg_q1616 AND symb_decoder(16#60#)) OR
 					(reg_q1616 AND symb_decoder(16#b3#)) OR
 					(reg_q1616 AND symb_decoder(16#b6#)) OR
 					(reg_q1616 AND symb_decoder(16#ab#)) OR
 					(reg_q1616 AND symb_decoder(16#2a#)) OR
 					(reg_q1616 AND symb_decoder(16#3a#)) OR
 					(reg_q1616 AND symb_decoder(16#bd#)) OR
 					(reg_q1616 AND symb_decoder(16#8b#)) OR
 					(reg_q1616 AND symb_decoder(16#fb#)) OR
 					(reg_q1616 AND symb_decoder(16#a3#)) OR
 					(reg_q1616 AND symb_decoder(16#30#)) OR
 					(reg_q1616 AND symb_decoder(16#98#)) OR
 					(reg_q1616 AND symb_decoder(16#5d#)) OR
 					(reg_q1616 AND symb_decoder(16#47#)) OR
 					(reg_q1616 AND symb_decoder(16#68#)) OR
 					(reg_q1616 AND symb_decoder(16#4a#)) OR
 					(reg_q1616 AND symb_decoder(16#c4#)) OR
 					(reg_q1616 AND symb_decoder(16#6b#)) OR
 					(reg_q1616 AND symb_decoder(16#9f#)) OR
 					(reg_q1616 AND symb_decoder(16#7e#)) OR
 					(reg_q1616 AND symb_decoder(16#a1#)) OR
 					(reg_q1616 AND symb_decoder(16#e9#)) OR
 					(reg_q1616 AND symb_decoder(16#f3#)) OR
 					(reg_q1616 AND symb_decoder(16#c6#)) OR
 					(reg_q1616 AND symb_decoder(16#17#)) OR
 					(reg_q1616 AND symb_decoder(16#32#)) OR
 					(reg_q1616 AND symb_decoder(16#43#)) OR
 					(reg_q1616 AND symb_decoder(16#d9#)) OR
 					(reg_q1616 AND symb_decoder(16#16#)) OR
 					(reg_q1616 AND symb_decoder(16#97#)) OR
 					(reg_q1616 AND symb_decoder(16#bc#)) OR
 					(reg_q1616 AND symb_decoder(16#25#)) OR
 					(reg_q1616 AND symb_decoder(16#a5#)) OR
 					(reg_q1616 AND symb_decoder(16#39#)) OR
 					(reg_q1616 AND symb_decoder(16#0b#)) OR
 					(reg_q1616 AND symb_decoder(16#5a#)) OR
 					(reg_q1616 AND symb_decoder(16#34#)) OR
 					(reg_q1616 AND symb_decoder(16#4b#)) OR
 					(reg_q1616 AND symb_decoder(16#91#)) OR
 					(reg_q1616 AND symb_decoder(16#dd#)) OR
 					(reg_q1616 AND symb_decoder(16#71#)) OR
 					(reg_q1616 AND symb_decoder(16#87#)) OR
 					(reg_q1616 AND symb_decoder(16#4f#)) OR
 					(reg_q1616 AND symb_decoder(16#e8#)) OR
 					(reg_q1616 AND symb_decoder(16#96#)) OR
 					(reg_q1616 AND symb_decoder(16#9a#)) OR
 					(reg_q1616 AND symb_decoder(16#99#)) OR
 					(reg_q1616 AND symb_decoder(16#1f#)) OR
 					(reg_q1616 AND symb_decoder(16#7f#)) OR
 					(reg_q1616 AND symb_decoder(16#56#)) OR
 					(reg_q1616 AND symb_decoder(16#f2#)) OR
 					(reg_q1616 AND symb_decoder(16#88#)) OR
 					(reg_q1616 AND symb_decoder(16#4c#)) OR
 					(reg_q1616 AND symb_decoder(16#ad#)) OR
 					(reg_q1616 AND symb_decoder(16#29#)) OR
 					(reg_q1616 AND symb_decoder(16#67#)) OR
 					(reg_q1616 AND symb_decoder(16#ed#)) OR
 					(reg_q1616 AND symb_decoder(16#73#)) OR
 					(reg_q1616 AND symb_decoder(16#8e#)) OR
 					(reg_q1616 AND symb_decoder(16#a4#)) OR
 					(reg_q1616 AND symb_decoder(16#4e#)) OR
 					(reg_q1616 AND symb_decoder(16#01#)) OR
 					(reg_q1616 AND symb_decoder(16#84#)) OR
 					(reg_q1616 AND symb_decoder(16#be#)) OR
 					(reg_q1616 AND symb_decoder(16#9b#)) OR
 					(reg_q1616 AND symb_decoder(16#31#)) OR
 					(reg_q1616 AND symb_decoder(16#1b#)) OR
 					(reg_q1616 AND symb_decoder(16#ef#)) OR
 					(reg_q1616 AND symb_decoder(16#ba#)) OR
 					(reg_q1616 AND symb_decoder(16#2d#)) OR
 					(reg_q1616 AND symb_decoder(16#09#)) OR
 					(reg_q1616 AND symb_decoder(16#35#)) OR
 					(reg_q1616 AND symb_decoder(16#ce#)) OR
 					(reg_q1616 AND symb_decoder(16#c7#)) OR
 					(reg_q1616 AND symb_decoder(16#f6#)) OR
 					(reg_q1616 AND symb_decoder(16#c0#)) OR
 					(reg_q1616 AND symb_decoder(16#eb#)) OR
 					(reg_q1616 AND symb_decoder(16#bf#)) OR
 					(reg_q1616 AND symb_decoder(16#8c#)) OR
 					(reg_q1616 AND symb_decoder(16#15#)) OR
 					(reg_q1616 AND symb_decoder(16#e6#)) OR
 					(reg_q1616 AND symb_decoder(16#55#)) OR
 					(reg_q1616 AND symb_decoder(16#62#)) OR
 					(reg_q1616 AND symb_decoder(16#77#)) OR
 					(reg_q1616 AND symb_decoder(16#f0#)) OR
 					(reg_q1616 AND symb_decoder(16#c3#)) OR
 					(reg_q1616 AND symb_decoder(16#20#)) OR
 					(reg_q1616 AND symb_decoder(16#e1#)) OR
 					(reg_q1616 AND symb_decoder(16#05#)) OR
 					(reg_q1616 AND symb_decoder(16#e5#)) OR
 					(reg_q1616 AND symb_decoder(16#a9#)) OR
 					(reg_q1616 AND symb_decoder(16#70#)) OR
 					(reg_q1616 AND symb_decoder(16#d8#)) OR
 					(reg_q1616 AND symb_decoder(16#da#)) OR
 					(reg_q1616 AND symb_decoder(16#59#)) OR
 					(reg_q1616 AND symb_decoder(16#fc#)) OR
 					(reg_q1616 AND symb_decoder(16#5b#)) OR
 					(reg_q1616 AND symb_decoder(16#1e#)) OR
 					(reg_q1616 AND symb_decoder(16#7b#)) OR
 					(reg_q1616 AND symb_decoder(16#f5#)) OR
 					(reg_q1616 AND symb_decoder(16#52#)) OR
 					(reg_q1616 AND symb_decoder(16#f9#)) OR
 					(reg_q1616 AND symb_decoder(16#12#)) OR
 					(reg_q1616 AND symb_decoder(16#61#)) OR
 					(reg_q1616 AND symb_decoder(16#49#)) OR
 					(reg_q1616 AND symb_decoder(16#51#)) OR
 					(reg_q1616 AND symb_decoder(16#3e#)) OR
 					(reg_q1616 AND symb_decoder(16#94#)) OR
 					(reg_q1616 AND symb_decoder(16#50#)) OR
 					(reg_q1616 AND symb_decoder(16#78#)) OR
 					(reg_q1616 AND symb_decoder(16#df#)) OR
 					(reg_q1616 AND symb_decoder(16#85#)) OR
 					(reg_q1616 AND symb_decoder(16#28#)) OR
 					(reg_q1616 AND symb_decoder(16#10#)) OR
 					(reg_q1616 AND symb_decoder(16#db#)) OR
 					(reg_q1616 AND symb_decoder(16#41#)) OR
 					(reg_q1616 AND symb_decoder(16#64#)) OR
 					(reg_q1616 AND symb_decoder(16#53#)) OR
 					(reg_q1616 AND symb_decoder(16#b4#)) OR
 					(reg_q1616 AND symb_decoder(16#2e#)) OR
 					(reg_q1616 AND symb_decoder(16#6d#)) OR
 					(reg_q1616 AND symb_decoder(16#69#)) OR
 					(reg_q1616 AND symb_decoder(16#b8#)) OR
 					(reg_q1616 AND symb_decoder(16#ca#)) OR
 					(reg_q1616 AND symb_decoder(16#23#)) OR
 					(reg_q1616 AND symb_decoder(16#d6#)) OR
 					(reg_q1616 AND symb_decoder(16#5f#)) OR
 					(reg_q1616 AND symb_decoder(16#90#)) OR
 					(reg_q1616 AND symb_decoder(16#a2#)) OR
 					(reg_q1616 AND symb_decoder(16#b2#)) OR
 					(reg_q1616 AND symb_decoder(16#0e#)) OR
 					(reg_q1616 AND symb_decoder(16#76#)) OR
 					(reg_q1616 AND symb_decoder(16#65#)) OR
 					(reg_q1616 AND symb_decoder(16#b1#)) OR
 					(reg_q1616 AND symb_decoder(16#95#)) OR
 					(reg_q1616 AND symb_decoder(16#54#)) OR
 					(reg_q1616 AND symb_decoder(16#d1#)) OR
 					(reg_q1616 AND symb_decoder(16#46#)) OR
 					(reg_q1616 AND symb_decoder(16#6e#)) OR
 					(reg_q1616 AND symb_decoder(16#18#)) OR
 					(reg_q1616 AND symb_decoder(16#36#)) OR
 					(reg_q1616 AND symb_decoder(16#b5#)) OR
 					(reg_q1616 AND symb_decoder(16#00#)) OR
 					(reg_q1616 AND symb_decoder(16#57#)) OR
 					(reg_q1616 AND symb_decoder(16#5e#)) OR
 					(reg_q1616 AND symb_decoder(16#3c#)) OR
 					(reg_q1616 AND symb_decoder(16#7d#)) OR
 					(reg_q1616 AND symb_decoder(16#66#)) OR
 					(reg_q1616 AND symb_decoder(16#d3#)) OR
 					(reg_q1616 AND symb_decoder(16#1c#)) OR
 					(reg_q1616 AND symb_decoder(16#37#)) OR
 					(reg_q1616 AND symb_decoder(16#7c#)) OR
 					(reg_q1616 AND symb_decoder(16#fd#)) OR
 					(reg_q1616 AND symb_decoder(16#3f#)) OR
 					(reg_q1616 AND symb_decoder(16#33#)) OR
 					(reg_q1616 AND symb_decoder(16#06#)) OR
 					(reg_q1616 AND symb_decoder(16#89#)) OR
 					(reg_q1616 AND symb_decoder(16#fe#)) OR
 					(reg_q1616 AND symb_decoder(16#b0#)) OR
 					(reg_q1616 AND symb_decoder(16#ee#)) OR
 					(reg_q1616 AND symb_decoder(16#bb#)) OR
 					(reg_q1616 AND symb_decoder(16#9e#)) OR
 					(reg_q1616 AND symb_decoder(16#a7#)) OR
 					(reg_q1616 AND symb_decoder(16#7a#)) OR
 					(reg_q1616 AND symb_decoder(16#03#)) OR
 					(reg_q1616 AND symb_decoder(16#c5#)) OR
 					(reg_q1616 AND symb_decoder(16#8f#)) OR
 					(reg_q1616 AND symb_decoder(16#21#)) OR
 					(reg_q1616 AND symb_decoder(16#4d#)) OR
 					(reg_q1616 AND symb_decoder(16#d0#)) OR
 					(reg_q1616 AND symb_decoder(16#aa#)) OR
 					(reg_q1616 AND symb_decoder(16#cc#)) OR
 					(reg_q1616 AND symb_decoder(16#48#)) OR
 					(reg_q1616 AND symb_decoder(16#e0#)) OR
 					(reg_q1616 AND symb_decoder(16#f4#)) OR
 					(reg_q1616 AND symb_decoder(16#f7#)) OR
 					(reg_q1616 AND symb_decoder(16#63#)) OR
 					(reg_q1616 AND symb_decoder(16#c9#)) OR
 					(reg_q1616 AND symb_decoder(16#ff#)) OR
 					(reg_q1616 AND symb_decoder(16#ea#)) OR
 					(reg_q1616 AND symb_decoder(16#81#)) OR
 					(reg_q1616 AND symb_decoder(16#cd#)) OR
 					(reg_q1616 AND symb_decoder(16#22#)) OR
 					(reg_q1616 AND symb_decoder(16#6f#)) OR
 					(reg_q1616 AND symb_decoder(16#07#)) OR
 					(reg_q1616 AND symb_decoder(16#d7#)) OR
 					(reg_q1616 AND symb_decoder(16#c1#)) OR
 					(reg_q1616 AND symb_decoder(16#58#)) OR
 					(reg_q1616 AND symb_decoder(16#c2#)) OR
 					(reg_q1616 AND symb_decoder(16#9c#)) OR
 					(reg_q1616 AND symb_decoder(16#f8#)) OR
 					(reg_q1616 AND symb_decoder(16#f1#)) OR
 					(reg_q1616 AND symb_decoder(16#26#)) OR
 					(reg_q1616 AND symb_decoder(16#8a#)) OR
 					(reg_q1616 AND symb_decoder(16#dc#)) OR
 					(reg_q1616 AND symb_decoder(16#6c#)) OR
 					(reg_q1616 AND symb_decoder(16#27#)) OR
 					(reg_q1616 AND symb_decoder(16#e2#)) OR
 					(reg_q1616 AND symb_decoder(16#b7#)) OR
 					(reg_q1616 AND symb_decoder(16#38#)) OR
 					(reg_q1616 AND symb_decoder(16#5c#)) OR
 					(reg_q1616 AND symb_decoder(16#6a#)) OR
 					(reg_q1616 AND symb_decoder(16#93#)) OR
 					(reg_q1616 AND symb_decoder(16#2f#)) OR
 					(reg_q1616 AND symb_decoder(16#75#)) OR
 					(reg_q1616 AND symb_decoder(16#a8#)) OR
 					(reg_q1616 AND symb_decoder(16#40#)) OR
 					(reg_q1616 AND symb_decoder(16#08#)) OR
 					(reg_q1616 AND symb_decoder(16#45#)) OR
 					(reg_q1616 AND symb_decoder(16#8d#)) OR
 					(reg_q1616 AND symb_decoder(16#c8#)) OR
 					(reg_q1616 AND symb_decoder(16#ac#)) OR
 					(reg_q1616 AND symb_decoder(16#86#)) OR
 					(reg_q1616 AND symb_decoder(16#9d#)) OR
 					(reg_q1616 AND symb_decoder(16#e3#)) OR
 					(reg_q1616 AND symb_decoder(16#d2#)) OR
 					(reg_q1616 AND symb_decoder(16#13#)) OR
 					(reg_q1616 AND symb_decoder(16#de#)) OR
 					(reg_q1616 AND symb_decoder(16#3b#));
reg_q471_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q470 AND symb_decoder(16#0d#)) OR
 					(reg_q470 AND symb_decoder(16#0a#));
reg_q759_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q758 AND symb_decoder(16#53#)) OR
 					(reg_q758 AND symb_decoder(16#73#));
reg_fullgraph28_init <= "00";

reg_fullgraph28_sel <= "0" & reg_q759_in & reg_q471_in & reg_q1626_in;

	--coder fullgraph28
with reg_fullgraph28_sel select
reg_fullgraph28_in <=
	"01" when "0001",
	"10" when "0010",
	"11" when "0100",
	"00" when others;
 --end coder

	p_reg_fullgraph28: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph28 <= reg_fullgraph28_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph28 <= reg_fullgraph28_init;
        else
          reg_fullgraph28 <= reg_fullgraph28_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph28

		reg_q1626 <= '1' when reg_fullgraph28 = "01" else '0'; 
		reg_q471 <= '1' when reg_fullgraph28 = "10" else '0'; 
		reg_q759 <= '1' when reg_fullgraph28 = "11" else '0'; 
--end decoder 

reg_q1951_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1951 AND symb_decoder(16#9c#)) OR
 					(reg_q1951 AND symb_decoder(16#ec#)) OR
 					(reg_q1951 AND symb_decoder(16#81#)) OR
 					(reg_q1951 AND symb_decoder(16#d7#)) OR
 					(reg_q1951 AND symb_decoder(16#8d#)) OR
 					(reg_q1951 AND symb_decoder(16#8e#)) OR
 					(reg_q1951 AND symb_decoder(16#ea#)) OR
 					(reg_q1951 AND symb_decoder(16#44#)) OR
 					(reg_q1951 AND symb_decoder(16#01#)) OR
 					(reg_q1951 AND symb_decoder(16#89#)) OR
 					(reg_q1951 AND symb_decoder(16#67#)) OR
 					(reg_q1951 AND symb_decoder(16#be#)) OR
 					(reg_q1951 AND symb_decoder(16#5f#)) OR
 					(reg_q1951 AND symb_decoder(16#b5#)) OR
 					(reg_q1951 AND symb_decoder(16#c1#)) OR
 					(reg_q1951 AND symb_decoder(16#31#)) OR
 					(reg_q1951 AND symb_decoder(16#5b#)) OR
 					(reg_q1951 AND symb_decoder(16#66#)) OR
 					(reg_q1951 AND symb_decoder(16#e6#)) OR
 					(reg_q1951 AND symb_decoder(16#0d#)) OR
 					(reg_q1951 AND symb_decoder(16#c4#)) OR
 					(reg_q1951 AND symb_decoder(16#6e#)) OR
 					(reg_q1951 AND symb_decoder(16#14#)) OR
 					(reg_q1951 AND symb_decoder(16#a5#)) OR
 					(reg_q1951 AND symb_decoder(16#6c#)) OR
 					(reg_q1951 AND symb_decoder(16#45#)) OR
 					(reg_q1951 AND symb_decoder(16#f6#)) OR
 					(reg_q1951 AND symb_decoder(16#ee#)) OR
 					(reg_q1951 AND symb_decoder(16#2c#)) OR
 					(reg_q1951 AND symb_decoder(16#a7#)) OR
 					(reg_q1951 AND symb_decoder(16#eb#)) OR
 					(reg_q1951 AND symb_decoder(16#97#)) OR
 					(reg_q1951 AND symb_decoder(16#84#)) OR
 					(reg_q1951 AND symb_decoder(16#5c#)) OR
 					(reg_q1951 AND symb_decoder(16#1c#)) OR
 					(reg_q1951 AND symb_decoder(16#a1#)) OR
 					(reg_q1951 AND symb_decoder(16#d5#)) OR
 					(reg_q1951 AND symb_decoder(16#7c#)) OR
 					(reg_q1951 AND symb_decoder(16#86#)) OR
 					(reg_q1951 AND symb_decoder(16#43#)) OR
 					(reg_q1951 AND symb_decoder(16#20#)) OR
 					(reg_q1951 AND symb_decoder(16#f5#)) OR
 					(reg_q1951 AND symb_decoder(16#ca#)) OR
 					(reg_q1951 AND symb_decoder(16#ab#)) OR
 					(reg_q1951 AND symb_decoder(16#fc#)) OR
 					(reg_q1951 AND symb_decoder(16#6a#)) OR
 					(reg_q1951 AND symb_decoder(16#c0#)) OR
 					(reg_q1951 AND symb_decoder(16#88#)) OR
 					(reg_q1951 AND symb_decoder(16#ac#)) OR
 					(reg_q1951 AND symb_decoder(16#35#)) OR
 					(reg_q1951 AND symb_decoder(16#98#)) OR
 					(reg_q1951 AND symb_decoder(16#ef#)) OR
 					(reg_q1951 AND symb_decoder(16#2b#)) OR
 					(reg_q1951 AND symb_decoder(16#17#)) OR
 					(reg_q1951 AND symb_decoder(16#49#)) OR
 					(reg_q1951 AND symb_decoder(16#55#)) OR
 					(reg_q1951 AND symb_decoder(16#a9#)) OR
 					(reg_q1951 AND symb_decoder(16#33#)) OR
 					(reg_q1951 AND symb_decoder(16#2e#)) OR
 					(reg_q1951 AND symb_decoder(16#d0#)) OR
 					(reg_q1951 AND symb_decoder(16#b0#)) OR
 					(reg_q1951 AND symb_decoder(16#df#)) OR
 					(reg_q1951 AND symb_decoder(16#a3#)) OR
 					(reg_q1951 AND symb_decoder(16#5d#)) OR
 					(reg_q1951 AND symb_decoder(16#1b#)) OR
 					(reg_q1951 AND symb_decoder(16#f2#)) OR
 					(reg_q1951 AND symb_decoder(16#04#)) OR
 					(reg_q1951 AND symb_decoder(16#c7#)) OR
 					(reg_q1951 AND symb_decoder(16#1d#)) OR
 					(reg_q1951 AND symb_decoder(16#cf#)) OR
 					(reg_q1951 AND symb_decoder(16#06#)) OR
 					(reg_q1951 AND symb_decoder(16#aa#)) OR
 					(reg_q1951 AND symb_decoder(16#1a#)) OR
 					(reg_q1951 AND symb_decoder(16#16#)) OR
 					(reg_q1951 AND symb_decoder(16#8a#)) OR
 					(reg_q1951 AND symb_decoder(16#e4#)) OR
 					(reg_q1951 AND symb_decoder(16#21#)) OR
 					(reg_q1951 AND symb_decoder(16#4c#)) OR
 					(reg_q1951 AND symb_decoder(16#0e#)) OR
 					(reg_q1951 AND symb_decoder(16#72#)) OR
 					(reg_q1951 AND symb_decoder(16#db#)) OR
 					(reg_q1951 AND symb_decoder(16#c2#)) OR
 					(reg_q1951 AND symb_decoder(16#e1#)) OR
 					(reg_q1951 AND symb_decoder(16#74#)) OR
 					(reg_q1951 AND symb_decoder(16#f8#)) OR
 					(reg_q1951 AND symb_decoder(16#71#)) OR
 					(reg_q1951 AND symb_decoder(16#99#)) OR
 					(reg_q1951 AND symb_decoder(16#4f#)) OR
 					(reg_q1951 AND symb_decoder(16#10#)) OR
 					(reg_q1951 AND symb_decoder(16#27#)) OR
 					(reg_q1951 AND symb_decoder(16#3c#)) OR
 					(reg_q1951 AND symb_decoder(16#b6#)) OR
 					(reg_q1951 AND symb_decoder(16#b1#)) OR
 					(reg_q1951 AND symb_decoder(16#c6#)) OR
 					(reg_q1951 AND symb_decoder(16#51#)) OR
 					(reg_q1951 AND symb_decoder(16#58#)) OR
 					(reg_q1951 AND symb_decoder(16#3e#)) OR
 					(reg_q1951 AND symb_decoder(16#25#)) OR
 					(reg_q1951 AND symb_decoder(16#e8#)) OR
 					(reg_q1951 AND symb_decoder(16#90#)) OR
 					(reg_q1951 AND symb_decoder(16#6b#)) OR
 					(reg_q1951 AND symb_decoder(16#dd#)) OR
 					(reg_q1951 AND symb_decoder(16#8b#)) OR
 					(reg_q1951 AND symb_decoder(16#59#)) OR
 					(reg_q1951 AND symb_decoder(16#57#)) OR
 					(reg_q1951 AND symb_decoder(16#70#)) OR
 					(reg_q1951 AND symb_decoder(16#96#)) OR
 					(reg_q1951 AND symb_decoder(16#36#)) OR
 					(reg_q1951 AND symb_decoder(16#c5#)) OR
 					(reg_q1951 AND symb_decoder(16#76#)) OR
 					(reg_q1951 AND symb_decoder(16#b8#)) OR
 					(reg_q1951 AND symb_decoder(16#7a#)) OR
 					(reg_q1951 AND symb_decoder(16#f7#)) OR
 					(reg_q1951 AND symb_decoder(16#b4#)) OR
 					(reg_q1951 AND symb_decoder(16#8c#)) OR
 					(reg_q1951 AND symb_decoder(16#e5#)) OR
 					(reg_q1951 AND symb_decoder(16#95#)) OR
 					(reg_q1951 AND symb_decoder(16#6d#)) OR
 					(reg_q1951 AND symb_decoder(16#fe#)) OR
 					(reg_q1951 AND symb_decoder(16#a6#)) OR
 					(reg_q1951 AND symb_decoder(16#bb#)) OR
 					(reg_q1951 AND symb_decoder(16#d2#)) OR
 					(reg_q1951 AND symb_decoder(16#f0#)) OR
 					(reg_q1951 AND symb_decoder(16#a4#)) OR
 					(reg_q1951 AND symb_decoder(16#46#)) OR
 					(reg_q1951 AND symb_decoder(16#da#)) OR
 					(reg_q1951 AND symb_decoder(16#7b#)) OR
 					(reg_q1951 AND symb_decoder(16#ad#)) OR
 					(reg_q1951 AND symb_decoder(16#6f#)) OR
 					(reg_q1951 AND symb_decoder(16#30#)) OR
 					(reg_q1951 AND symb_decoder(16#9a#)) OR
 					(reg_q1951 AND symb_decoder(16#ae#)) OR
 					(reg_q1951 AND symb_decoder(16#3f#)) OR
 					(reg_q1951 AND symb_decoder(16#5a#)) OR
 					(reg_q1951 AND symb_decoder(16#08#)) OR
 					(reg_q1951 AND symb_decoder(16#42#)) OR
 					(reg_q1951 AND symb_decoder(16#3a#)) OR
 					(reg_q1951 AND symb_decoder(16#0b#)) OR
 					(reg_q1951 AND symb_decoder(16#53#)) OR
 					(reg_q1951 AND symb_decoder(16#62#)) OR
 					(reg_q1951 AND symb_decoder(16#00#)) OR
 					(reg_q1951 AND symb_decoder(16#cc#)) OR
 					(reg_q1951 AND symb_decoder(16#1f#)) OR
 					(reg_q1951 AND symb_decoder(16#41#)) OR
 					(reg_q1951 AND symb_decoder(16#2a#)) OR
 					(reg_q1951 AND symb_decoder(16#d1#)) OR
 					(reg_q1951 AND symb_decoder(16#9b#)) OR
 					(reg_q1951 AND symb_decoder(16#85#)) OR
 					(reg_q1951 AND symb_decoder(16#92#)) OR
 					(reg_q1951 AND symb_decoder(16#2d#)) OR
 					(reg_q1951 AND symb_decoder(16#d8#)) OR
 					(reg_q1951 AND symb_decoder(16#37#)) OR
 					(reg_q1951 AND symb_decoder(16#a0#)) OR
 					(reg_q1951 AND symb_decoder(16#65#)) OR
 					(reg_q1951 AND symb_decoder(16#26#)) OR
 					(reg_q1951 AND symb_decoder(16#02#)) OR
 					(reg_q1951 AND symb_decoder(16#7d#)) OR
 					(reg_q1951 AND symb_decoder(16#c9#)) OR
 					(reg_q1951 AND symb_decoder(16#f1#)) OR
 					(reg_q1951 AND symb_decoder(16#dc#)) OR
 					(reg_q1951 AND symb_decoder(16#cd#)) OR
 					(reg_q1951 AND symb_decoder(16#ce#)) OR
 					(reg_q1951 AND symb_decoder(16#80#)) OR
 					(reg_q1951 AND symb_decoder(16#9e#)) OR
 					(reg_q1951 AND symb_decoder(16#13#)) OR
 					(reg_q1951 AND symb_decoder(16#73#)) OR
 					(reg_q1951 AND symb_decoder(16#56#)) OR
 					(reg_q1951 AND symb_decoder(16#ff#)) OR
 					(reg_q1951 AND symb_decoder(16#f4#)) OR
 					(reg_q1951 AND symb_decoder(16#e0#)) OR
 					(reg_q1951 AND symb_decoder(16#79#)) OR
 					(reg_q1951 AND symb_decoder(16#63#)) OR
 					(reg_q1951 AND symb_decoder(16#78#)) OR
 					(reg_q1951 AND symb_decoder(16#28#)) OR
 					(reg_q1951 AND symb_decoder(16#e7#)) OR
 					(reg_q1951 AND symb_decoder(16#5e#)) OR
 					(reg_q1951 AND symb_decoder(16#d4#)) OR
 					(reg_q1951 AND symb_decoder(16#50#)) OR
 					(reg_q1951 AND symb_decoder(16#ed#)) OR
 					(reg_q1951 AND symb_decoder(16#d6#)) OR
 					(reg_q1951 AND symb_decoder(16#e9#)) OR
 					(reg_q1951 AND symb_decoder(16#cb#)) OR
 					(reg_q1951 AND symb_decoder(16#07#)) OR
 					(reg_q1951 AND symb_decoder(16#38#)) OR
 					(reg_q1951 AND symb_decoder(16#94#)) OR
 					(reg_q1951 AND symb_decoder(16#09#)) OR
 					(reg_q1951 AND symb_decoder(16#3d#)) OR
 					(reg_q1951 AND symb_decoder(16#0c#)) OR
 					(reg_q1951 AND symb_decoder(16#8f#)) OR
 					(reg_q1951 AND symb_decoder(16#15#)) OR
 					(reg_q1951 AND symb_decoder(16#54#)) OR
 					(reg_q1951 AND symb_decoder(16#0f#)) OR
 					(reg_q1951 AND symb_decoder(16#b3#)) OR
 					(reg_q1951 AND symb_decoder(16#4d#)) OR
 					(reg_q1951 AND symb_decoder(16#de#)) OR
 					(reg_q1951 AND symb_decoder(16#77#)) OR
 					(reg_q1951 AND symb_decoder(16#19#)) OR
 					(reg_q1951 AND symb_decoder(16#29#)) OR
 					(reg_q1951 AND symb_decoder(16#22#)) OR
 					(reg_q1951 AND symb_decoder(16#2f#)) OR
 					(reg_q1951 AND symb_decoder(16#c3#)) OR
 					(reg_q1951 AND symb_decoder(16#23#)) OR
 					(reg_q1951 AND symb_decoder(16#03#)) OR
 					(reg_q1951 AND symb_decoder(16#9d#)) OR
 					(reg_q1951 AND symb_decoder(16#e3#)) OR
 					(reg_q1951 AND symb_decoder(16#52#)) OR
 					(reg_q1951 AND symb_decoder(16#64#)) OR
 					(reg_q1951 AND symb_decoder(16#ba#)) OR
 					(reg_q1951 AND symb_decoder(16#91#)) OR
 					(reg_q1951 AND symb_decoder(16#0a#)) OR
 					(reg_q1951 AND symb_decoder(16#18#)) OR
 					(reg_q1951 AND symb_decoder(16#39#)) OR
 					(reg_q1951 AND symb_decoder(16#11#)) OR
 					(reg_q1951 AND symb_decoder(16#a8#)) OR
 					(reg_q1951 AND symb_decoder(16#87#)) OR
 					(reg_q1951 AND symb_decoder(16#d9#)) OR
 					(reg_q1951 AND symb_decoder(16#82#)) OR
 					(reg_q1951 AND symb_decoder(16#83#)) OR
 					(reg_q1951 AND symb_decoder(16#61#)) OR
 					(reg_q1951 AND symb_decoder(16#af#)) OR
 					(reg_q1951 AND symb_decoder(16#fa#)) OR
 					(reg_q1951 AND symb_decoder(16#75#)) OR
 					(reg_q1951 AND symb_decoder(16#c8#)) OR
 					(reg_q1951 AND symb_decoder(16#9f#)) OR
 					(reg_q1951 AND symb_decoder(16#60#)) OR
 					(reg_q1951 AND symb_decoder(16#bf#)) OR
 					(reg_q1951 AND symb_decoder(16#bd#)) OR
 					(reg_q1951 AND symb_decoder(16#b9#)) OR
 					(reg_q1951 AND symb_decoder(16#48#)) OR
 					(reg_q1951 AND symb_decoder(16#b2#)) OR
 					(reg_q1951 AND symb_decoder(16#bc#)) OR
 					(reg_q1951 AND symb_decoder(16#47#)) OR
 					(reg_q1951 AND symb_decoder(16#3b#)) OR
 					(reg_q1951 AND symb_decoder(16#4a#)) OR
 					(reg_q1951 AND symb_decoder(16#4b#)) OR
 					(reg_q1951 AND symb_decoder(16#d3#)) OR
 					(reg_q1951 AND symb_decoder(16#05#)) OR
 					(reg_q1951 AND symb_decoder(16#68#)) OR
 					(reg_q1951 AND symb_decoder(16#b7#)) OR
 					(reg_q1951 AND symb_decoder(16#e2#)) OR
 					(reg_q1951 AND symb_decoder(16#69#)) OR
 					(reg_q1951 AND symb_decoder(16#f9#)) OR
 					(reg_q1951 AND symb_decoder(16#93#)) OR
 					(reg_q1951 AND symb_decoder(16#1e#)) OR
 					(reg_q1951 AND symb_decoder(16#24#)) OR
 					(reg_q1951 AND symb_decoder(16#f3#)) OR
 					(reg_q1951 AND symb_decoder(16#32#)) OR
 					(reg_q1951 AND symb_decoder(16#34#)) OR
 					(reg_q1951 AND symb_decoder(16#12#)) OR
 					(reg_q1951 AND symb_decoder(16#4e#)) OR
 					(reg_q1951 AND symb_decoder(16#fb#)) OR
 					(reg_q1951 AND symb_decoder(16#fd#)) OR
 					(reg_q1951 AND symb_decoder(16#a2#)) OR
 					(reg_q1951 AND symb_decoder(16#40#)) OR
 					(reg_q1951 AND symb_decoder(16#7f#)) OR
 					(reg_q1951 AND symb_decoder(16#7e#));
reg_q1951_init <= '0' ;
	p_reg_q1951: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1951 <= reg_q1951_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1951 <= reg_q1951_init;
        else
          reg_q1951 <= reg_q1951_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2680_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q2680 AND symb_decoder(16#09#)) OR
 					(reg_q2680 AND symb_decoder(16#6c#)) OR
 					(reg_q2680 AND symb_decoder(16#41#)) OR
 					(reg_q2680 AND symb_decoder(16#29#)) OR
 					(reg_q2680 AND symb_decoder(16#87#)) OR
 					(reg_q2680 AND symb_decoder(16#0f#)) OR
 					(reg_q2680 AND symb_decoder(16#f1#)) OR
 					(reg_q2680 AND symb_decoder(16#61#)) OR
 					(reg_q2680 AND symb_decoder(16#d0#)) OR
 					(reg_q2680 AND symb_decoder(16#44#)) OR
 					(reg_q2680 AND symb_decoder(16#67#)) OR
 					(reg_q2680 AND symb_decoder(16#55#)) OR
 					(reg_q2680 AND symb_decoder(16#6b#)) OR
 					(reg_q2680 AND symb_decoder(16#bb#)) OR
 					(reg_q2680 AND symb_decoder(16#fb#)) OR
 					(reg_q2680 AND symb_decoder(16#2f#)) OR
 					(reg_q2680 AND symb_decoder(16#9a#)) OR
 					(reg_q2680 AND symb_decoder(16#a3#)) OR
 					(reg_q2680 AND symb_decoder(16#59#)) OR
 					(reg_q2680 AND symb_decoder(16#43#)) OR
 					(reg_q2680 AND symb_decoder(16#b5#)) OR
 					(reg_q2680 AND symb_decoder(16#a0#)) OR
 					(reg_q2680 AND symb_decoder(16#69#)) OR
 					(reg_q2680 AND symb_decoder(16#40#)) OR
 					(reg_q2680 AND symb_decoder(16#01#)) OR
 					(reg_q2680 AND symb_decoder(16#18#)) OR
 					(reg_q2680 AND symb_decoder(16#4d#)) OR
 					(reg_q2680 AND symb_decoder(16#bd#)) OR
 					(reg_q2680 AND symb_decoder(16#57#)) OR
 					(reg_q2680 AND symb_decoder(16#ee#)) OR
 					(reg_q2680 AND symb_decoder(16#9d#)) OR
 					(reg_q2680 AND symb_decoder(16#d3#)) OR
 					(reg_q2680 AND symb_decoder(16#39#)) OR
 					(reg_q2680 AND symb_decoder(16#93#)) OR
 					(reg_q2680 AND symb_decoder(16#07#)) OR
 					(reg_q2680 AND symb_decoder(16#98#)) OR
 					(reg_q2680 AND symb_decoder(16#fe#)) OR
 					(reg_q2680 AND symb_decoder(16#73#)) OR
 					(reg_q2680 AND symb_decoder(16#8f#)) OR
 					(reg_q2680 AND symb_decoder(16#71#)) OR
 					(reg_q2680 AND symb_decoder(16#d7#)) OR
 					(reg_q2680 AND symb_decoder(16#22#)) OR
 					(reg_q2680 AND symb_decoder(16#c7#)) OR
 					(reg_q2680 AND symb_decoder(16#33#)) OR
 					(reg_q2680 AND symb_decoder(16#62#)) OR
 					(reg_q2680 AND symb_decoder(16#e3#)) OR
 					(reg_q2680 AND symb_decoder(16#5f#)) OR
 					(reg_q2680 AND symb_decoder(16#1e#)) OR
 					(reg_q2680 AND symb_decoder(16#0a#)) OR
 					(reg_q2680 AND symb_decoder(16#cd#)) OR
 					(reg_q2680 AND symb_decoder(16#8e#)) OR
 					(reg_q2680 AND symb_decoder(16#a5#)) OR
 					(reg_q2680 AND symb_decoder(16#f0#)) OR
 					(reg_q2680 AND symb_decoder(16#bc#)) OR
 					(reg_q2680 AND symb_decoder(16#ba#)) OR
 					(reg_q2680 AND symb_decoder(16#e0#)) OR
 					(reg_q2680 AND symb_decoder(16#30#)) OR
 					(reg_q2680 AND symb_decoder(16#37#)) OR
 					(reg_q2680 AND symb_decoder(16#31#)) OR
 					(reg_q2680 AND symb_decoder(16#77#)) OR
 					(reg_q2680 AND symb_decoder(16#fd#)) OR
 					(reg_q2680 AND symb_decoder(16#3a#)) OR
 					(reg_q2680 AND symb_decoder(16#ef#)) OR
 					(reg_q2680 AND symb_decoder(16#b1#)) OR
 					(reg_q2680 AND symb_decoder(16#a8#)) OR
 					(reg_q2680 AND symb_decoder(16#f6#)) OR
 					(reg_q2680 AND symb_decoder(16#06#)) OR
 					(reg_q2680 AND symb_decoder(16#4a#)) OR
 					(reg_q2680 AND symb_decoder(16#fc#)) OR
 					(reg_q2680 AND symb_decoder(16#0b#)) OR
 					(reg_q2680 AND symb_decoder(16#e2#)) OR
 					(reg_q2680 AND symb_decoder(16#1a#)) OR
 					(reg_q2680 AND symb_decoder(16#8b#)) OR
 					(reg_q2680 AND symb_decoder(16#de#)) OR
 					(reg_q2680 AND symb_decoder(16#08#)) OR
 					(reg_q2680 AND symb_decoder(16#c5#)) OR
 					(reg_q2680 AND symb_decoder(16#ea#)) OR
 					(reg_q2680 AND symb_decoder(16#f8#)) OR
 					(reg_q2680 AND symb_decoder(16#15#)) OR
 					(reg_q2680 AND symb_decoder(16#38#)) OR
 					(reg_q2680 AND symb_decoder(16#c2#)) OR
 					(reg_q2680 AND symb_decoder(16#68#)) OR
 					(reg_q2680 AND symb_decoder(16#64#)) OR
 					(reg_q2680 AND symb_decoder(16#32#)) OR
 					(reg_q2680 AND symb_decoder(16#78#)) OR
 					(reg_q2680 AND symb_decoder(16#94#)) OR
 					(reg_q2680 AND symb_decoder(16#f9#)) OR
 					(reg_q2680 AND symb_decoder(16#97#)) OR
 					(reg_q2680 AND symb_decoder(16#36#)) OR
 					(reg_q2680 AND symb_decoder(16#90#)) OR
 					(reg_q2680 AND symb_decoder(16#af#)) OR
 					(reg_q2680 AND symb_decoder(16#1f#)) OR
 					(reg_q2680 AND symb_decoder(16#2c#)) OR
 					(reg_q2680 AND symb_decoder(16#2e#)) OR
 					(reg_q2680 AND symb_decoder(16#74#)) OR
 					(reg_q2680 AND symb_decoder(16#45#)) OR
 					(reg_q2680 AND symb_decoder(16#95#)) OR
 					(reg_q2680 AND symb_decoder(16#ae#)) OR
 					(reg_q2680 AND symb_decoder(16#9e#)) OR
 					(reg_q2680 AND symb_decoder(16#5b#)) OR
 					(reg_q2680 AND symb_decoder(16#86#)) OR
 					(reg_q2680 AND symb_decoder(16#0e#)) OR
 					(reg_q2680 AND symb_decoder(16#e4#)) OR
 					(reg_q2680 AND symb_decoder(16#7e#)) OR
 					(reg_q2680 AND symb_decoder(16#4f#)) OR
 					(reg_q2680 AND symb_decoder(16#23#)) OR
 					(reg_q2680 AND symb_decoder(16#89#)) OR
 					(reg_q2680 AND symb_decoder(16#8a#)) OR
 					(reg_q2680 AND symb_decoder(16#eb#)) OR
 					(reg_q2680 AND symb_decoder(16#ff#)) OR
 					(reg_q2680 AND symb_decoder(16#54#)) OR
 					(reg_q2680 AND symb_decoder(16#ca#)) OR
 					(reg_q2680 AND symb_decoder(16#6a#)) OR
 					(reg_q2680 AND symb_decoder(16#03#)) OR
 					(reg_q2680 AND symb_decoder(16#4b#)) OR
 					(reg_q2680 AND symb_decoder(16#a6#)) OR
 					(reg_q2680 AND symb_decoder(16#a2#)) OR
 					(reg_q2680 AND symb_decoder(16#df#)) OR
 					(reg_q2680 AND symb_decoder(16#7f#)) OR
 					(reg_q2680 AND symb_decoder(16#b0#)) OR
 					(reg_q2680 AND symb_decoder(16#91#)) OR
 					(reg_q2680 AND symb_decoder(16#76#)) OR
 					(reg_q2680 AND symb_decoder(16#81#)) OR
 					(reg_q2680 AND symb_decoder(16#da#)) OR
 					(reg_q2680 AND symb_decoder(16#05#)) OR
 					(reg_q2680 AND symb_decoder(16#b8#)) OR
 					(reg_q2680 AND symb_decoder(16#99#)) OR
 					(reg_q2680 AND symb_decoder(16#5c#)) OR
 					(reg_q2680 AND symb_decoder(16#53#)) OR
 					(reg_q2680 AND symb_decoder(16#27#)) OR
 					(reg_q2680 AND symb_decoder(16#e7#)) OR
 					(reg_q2680 AND symb_decoder(16#13#)) OR
 					(reg_q2680 AND symb_decoder(16#7a#)) OR
 					(reg_q2680 AND symb_decoder(16#a9#)) OR
 					(reg_q2680 AND symb_decoder(16#70#)) OR
 					(reg_q2680 AND symb_decoder(16#b6#)) OR
 					(reg_q2680 AND symb_decoder(16#6e#)) OR
 					(reg_q2680 AND symb_decoder(16#4c#)) OR
 					(reg_q2680 AND symb_decoder(16#00#)) OR
 					(reg_q2680 AND symb_decoder(16#b4#)) OR
 					(reg_q2680 AND symb_decoder(16#8c#)) OR
 					(reg_q2680 AND symb_decoder(16#a4#)) OR
 					(reg_q2680 AND symb_decoder(16#9c#)) OR
 					(reg_q2680 AND symb_decoder(16#dc#)) OR
 					(reg_q2680 AND symb_decoder(16#c4#)) OR
 					(reg_q2680 AND symb_decoder(16#cc#)) OR
 					(reg_q2680 AND symb_decoder(16#26#)) OR
 					(reg_q2680 AND symb_decoder(16#7c#)) OR
 					(reg_q2680 AND symb_decoder(16#0d#)) OR
 					(reg_q2680 AND symb_decoder(16#d9#)) OR
 					(reg_q2680 AND symb_decoder(16#0c#)) OR
 					(reg_q2680 AND symb_decoder(16#84#)) OR
 					(reg_q2680 AND symb_decoder(16#5a#)) OR
 					(reg_q2680 AND symb_decoder(16#ce#)) OR
 					(reg_q2680 AND symb_decoder(16#ec#)) OR
 					(reg_q2680 AND symb_decoder(16#42#)) OR
 					(reg_q2680 AND symb_decoder(16#ed#)) OR
 					(reg_q2680 AND symb_decoder(16#75#)) OR
 					(reg_q2680 AND symb_decoder(16#e5#)) OR
 					(reg_q2680 AND symb_decoder(16#c0#)) OR
 					(reg_q2680 AND symb_decoder(16#f4#)) OR
 					(reg_q2680 AND symb_decoder(16#24#)) OR
 					(reg_q2680 AND symb_decoder(16#72#)) OR
 					(reg_q2680 AND symb_decoder(16#3b#)) OR
 					(reg_q2680 AND symb_decoder(16#83#)) OR
 					(reg_q2680 AND symb_decoder(16#c6#)) OR
 					(reg_q2680 AND symb_decoder(16#25#)) OR
 					(reg_q2680 AND symb_decoder(16#51#)) OR
 					(reg_q2680 AND symb_decoder(16#6d#)) OR
 					(reg_q2680 AND symb_decoder(16#f3#)) OR
 					(reg_q2680 AND symb_decoder(16#db#)) OR
 					(reg_q2680 AND symb_decoder(16#96#)) OR
 					(reg_q2680 AND symb_decoder(16#d2#)) OR
 					(reg_q2680 AND symb_decoder(16#8d#)) OR
 					(reg_q2680 AND symb_decoder(16#63#)) OR
 					(reg_q2680 AND symb_decoder(16#56#)) OR
 					(reg_q2680 AND symb_decoder(16#e8#)) OR
 					(reg_q2680 AND symb_decoder(16#b3#)) OR
 					(reg_q2680 AND symb_decoder(16#65#)) OR
 					(reg_q2680 AND symb_decoder(16#d1#)) OR
 					(reg_q2680 AND symb_decoder(16#9f#)) OR
 					(reg_q2680 AND symb_decoder(16#be#)) OR
 					(reg_q2680 AND symb_decoder(16#3f#)) OR
 					(reg_q2680 AND symb_decoder(16#79#)) OR
 					(reg_q2680 AND symb_decoder(16#7d#)) OR
 					(reg_q2680 AND symb_decoder(16#3e#)) OR
 					(reg_q2680 AND symb_decoder(16#fa#)) OR
 					(reg_q2680 AND symb_decoder(16#46#)) OR
 					(reg_q2680 AND symb_decoder(16#47#)) OR
 					(reg_q2680 AND symb_decoder(16#3d#)) OR
 					(reg_q2680 AND symb_decoder(16#92#)) OR
 					(reg_q2680 AND symb_decoder(16#7b#)) OR
 					(reg_q2680 AND symb_decoder(16#b2#)) OR
 					(reg_q2680 AND symb_decoder(16#cb#)) OR
 					(reg_q2680 AND symb_decoder(16#28#)) OR
 					(reg_q2680 AND symb_decoder(16#2d#)) OR
 					(reg_q2680 AND symb_decoder(16#5e#)) OR
 					(reg_q2680 AND symb_decoder(16#17#)) OR
 					(reg_q2680 AND symb_decoder(16#a7#)) OR
 					(reg_q2680 AND symb_decoder(16#48#)) OR
 					(reg_q2680 AND symb_decoder(16#e6#)) OR
 					(reg_q2680 AND symb_decoder(16#10#)) OR
 					(reg_q2680 AND symb_decoder(16#80#)) OR
 					(reg_q2680 AND symb_decoder(16#19#)) OR
 					(reg_q2680 AND symb_decoder(16#11#)) OR
 					(reg_q2680 AND symb_decoder(16#cf#)) OR
 					(reg_q2680 AND symb_decoder(16#20#)) OR
 					(reg_q2680 AND symb_decoder(16#85#)) OR
 					(reg_q2680 AND symb_decoder(16#50#)) OR
 					(reg_q2680 AND symb_decoder(16#49#)) OR
 					(reg_q2680 AND symb_decoder(16#f2#)) OR
 					(reg_q2680 AND symb_decoder(16#21#)) OR
 					(reg_q2680 AND symb_decoder(16#14#)) OR
 					(reg_q2680 AND symb_decoder(16#60#)) OR
 					(reg_q2680 AND symb_decoder(16#2a#)) OR
 					(reg_q2680 AND symb_decoder(16#58#)) OR
 					(reg_q2680 AND symb_decoder(16#88#)) OR
 					(reg_q2680 AND symb_decoder(16#aa#)) OR
 					(reg_q2680 AND symb_decoder(16#4e#)) OR
 					(reg_q2680 AND symb_decoder(16#dd#)) OR
 					(reg_q2680 AND symb_decoder(16#35#)) OR
 					(reg_q2680 AND symb_decoder(16#bf#)) OR
 					(reg_q2680 AND symb_decoder(16#e9#)) OR
 					(reg_q2680 AND symb_decoder(16#d5#)) OR
 					(reg_q2680 AND symb_decoder(16#9b#)) OR
 					(reg_q2680 AND symb_decoder(16#c3#)) OR
 					(reg_q2680 AND symb_decoder(16#ad#)) OR
 					(reg_q2680 AND symb_decoder(16#6f#)) OR
 					(reg_q2680 AND symb_decoder(16#d6#)) OR
 					(reg_q2680 AND symb_decoder(16#12#)) OR
 					(reg_q2680 AND symb_decoder(16#e1#)) OR
 					(reg_q2680 AND symb_decoder(16#1b#)) OR
 					(reg_q2680 AND symb_decoder(16#a1#)) OR
 					(reg_q2680 AND symb_decoder(16#1d#)) OR
 					(reg_q2680 AND symb_decoder(16#f7#)) OR
 					(reg_q2680 AND symb_decoder(16#04#)) OR
 					(reg_q2680 AND symb_decoder(16#5d#)) OR
 					(reg_q2680 AND symb_decoder(16#ab#)) OR
 					(reg_q2680 AND symb_decoder(16#82#)) OR
 					(reg_q2680 AND symb_decoder(16#16#)) OR
 					(reg_q2680 AND symb_decoder(16#3c#)) OR
 					(reg_q2680 AND symb_decoder(16#34#)) OR
 					(reg_q2680 AND symb_decoder(16#d8#)) OR
 					(reg_q2680 AND symb_decoder(16#66#)) OR
 					(reg_q2680 AND symb_decoder(16#c1#)) OR
 					(reg_q2680 AND symb_decoder(16#52#)) OR
 					(reg_q2680 AND symb_decoder(16#b9#)) OR
 					(reg_q2680 AND symb_decoder(16#ac#)) OR
 					(reg_q2680 AND symb_decoder(16#c8#)) OR
 					(reg_q2680 AND symb_decoder(16#d4#)) OR
 					(reg_q2680 AND symb_decoder(16#1c#)) OR
 					(reg_q2680 AND symb_decoder(16#f5#)) OR
 					(reg_q2680 AND symb_decoder(16#c9#)) OR
 					(reg_q2680 AND symb_decoder(16#2b#)) OR
 					(reg_q2680 AND symb_decoder(16#b7#)) OR
 					(reg_q2680 AND symb_decoder(16#02#));
reg_q2680_init <= '0' ;
	p_reg_q2680: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2680 <= reg_q2680_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2680 <= reg_q2680_init;
        else
          reg_q2680 <= reg_q2680_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2417_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q2417 AND symb_decoder(16#de#)) OR
 					(reg_q2417 AND symb_decoder(16#46#)) OR
 					(reg_q2417 AND symb_decoder(16#cf#)) OR
 					(reg_q2417 AND symb_decoder(16#09#)) OR
 					(reg_q2417 AND symb_decoder(16#12#)) OR
 					(reg_q2417 AND symb_decoder(16#02#)) OR
 					(reg_q2417 AND symb_decoder(16#af#)) OR
 					(reg_q2417 AND symb_decoder(16#22#)) OR
 					(reg_q2417 AND symb_decoder(16#0a#)) OR
 					(reg_q2417 AND symb_decoder(16#26#)) OR
 					(reg_q2417 AND symb_decoder(16#21#)) OR
 					(reg_q2417 AND symb_decoder(16#82#)) OR
 					(reg_q2417 AND symb_decoder(16#a8#)) OR
 					(reg_q2417 AND symb_decoder(16#35#)) OR
 					(reg_q2417 AND symb_decoder(16#ca#)) OR
 					(reg_q2417 AND symb_decoder(16#90#)) OR
 					(reg_q2417 AND symb_decoder(16#d3#)) OR
 					(reg_q2417 AND symb_decoder(16#b8#)) OR
 					(reg_q2417 AND symb_decoder(16#8d#)) OR
 					(reg_q2417 AND symb_decoder(16#54#)) OR
 					(reg_q2417 AND symb_decoder(16#14#)) OR
 					(reg_q2417 AND symb_decoder(16#d4#)) OR
 					(reg_q2417 AND symb_decoder(16#f2#)) OR
 					(reg_q2417 AND symb_decoder(16#2e#)) OR
 					(reg_q2417 AND symb_decoder(16#a5#)) OR
 					(reg_q2417 AND symb_decoder(16#19#)) OR
 					(reg_q2417 AND symb_decoder(16#a6#)) OR
 					(reg_q2417 AND symb_decoder(16#6d#)) OR
 					(reg_q2417 AND symb_decoder(16#0e#)) OR
 					(reg_q2417 AND symb_decoder(16#1f#)) OR
 					(reg_q2417 AND symb_decoder(16#37#)) OR
 					(reg_q2417 AND symb_decoder(16#c6#)) OR
 					(reg_q2417 AND symb_decoder(16#6e#)) OR
 					(reg_q2417 AND symb_decoder(16#9d#)) OR
 					(reg_q2417 AND symb_decoder(16#bd#)) OR
 					(reg_q2417 AND symb_decoder(16#86#)) OR
 					(reg_q2417 AND symb_decoder(16#10#)) OR
 					(reg_q2417 AND symb_decoder(16#97#)) OR
 					(reg_q2417 AND symb_decoder(16#11#)) OR
 					(reg_q2417 AND symb_decoder(16#3c#)) OR
 					(reg_q2417 AND symb_decoder(16#88#)) OR
 					(reg_q2417 AND symb_decoder(16#61#)) OR
 					(reg_q2417 AND symb_decoder(16#91#)) OR
 					(reg_q2417 AND symb_decoder(16#7a#)) OR
 					(reg_q2417 AND symb_decoder(16#1a#)) OR
 					(reg_q2417 AND symb_decoder(16#bf#)) OR
 					(reg_q2417 AND symb_decoder(16#8c#)) OR
 					(reg_q2417 AND symb_decoder(16#c8#)) OR
 					(reg_q2417 AND symb_decoder(16#39#)) OR
 					(reg_q2417 AND symb_decoder(16#15#)) OR
 					(reg_q2417 AND symb_decoder(16#34#)) OR
 					(reg_q2417 AND symb_decoder(16#96#)) OR
 					(reg_q2417 AND symb_decoder(16#16#)) OR
 					(reg_q2417 AND symb_decoder(16#44#)) OR
 					(reg_q2417 AND symb_decoder(16#7b#)) OR
 					(reg_q2417 AND symb_decoder(16#ad#)) OR
 					(reg_q2417 AND symb_decoder(16#cd#)) OR
 					(reg_q2417 AND symb_decoder(16#9b#)) OR
 					(reg_q2417 AND symb_decoder(16#c9#)) OR
 					(reg_q2417 AND symb_decoder(16#98#)) OR
 					(reg_q2417 AND symb_decoder(16#e8#)) OR
 					(reg_q2417 AND symb_decoder(16#74#)) OR
 					(reg_q2417 AND symb_decoder(16#47#)) OR
 					(reg_q2417 AND symb_decoder(16#42#)) OR
 					(reg_q2417 AND symb_decoder(16#60#)) OR
 					(reg_q2417 AND symb_decoder(16#1e#)) OR
 					(reg_q2417 AND symb_decoder(16#a4#)) OR
 					(reg_q2417 AND symb_decoder(16#c2#)) OR
 					(reg_q2417 AND symb_decoder(16#e7#)) OR
 					(reg_q2417 AND symb_decoder(16#ed#)) OR
 					(reg_q2417 AND symb_decoder(16#06#)) OR
 					(reg_q2417 AND symb_decoder(16#58#)) OR
 					(reg_q2417 AND symb_decoder(16#57#)) OR
 					(reg_q2417 AND symb_decoder(16#e2#)) OR
 					(reg_q2417 AND symb_decoder(16#93#)) OR
 					(reg_q2417 AND symb_decoder(16#e0#)) OR
 					(reg_q2417 AND symb_decoder(16#1c#)) OR
 					(reg_q2417 AND symb_decoder(16#5e#)) OR
 					(reg_q2417 AND symb_decoder(16#9f#)) OR
 					(reg_q2417 AND symb_decoder(16#0f#)) OR
 					(reg_q2417 AND symb_decoder(16#b0#)) OR
 					(reg_q2417 AND symb_decoder(16#3d#)) OR
 					(reg_q2417 AND symb_decoder(16#b2#)) OR
 					(reg_q2417 AND symb_decoder(16#d0#)) OR
 					(reg_q2417 AND symb_decoder(16#65#)) OR
 					(reg_q2417 AND symb_decoder(16#a7#)) OR
 					(reg_q2417 AND symb_decoder(16#62#)) OR
 					(reg_q2417 AND symb_decoder(16#4d#)) OR
 					(reg_q2417 AND symb_decoder(16#f0#)) OR
 					(reg_q2417 AND symb_decoder(16#8b#)) OR
 					(reg_q2417 AND symb_decoder(16#78#)) OR
 					(reg_q2417 AND symb_decoder(16#a3#)) OR
 					(reg_q2417 AND symb_decoder(16#ec#)) OR
 					(reg_q2417 AND symb_decoder(16#40#)) OR
 					(reg_q2417 AND symb_decoder(16#83#)) OR
 					(reg_q2417 AND symb_decoder(16#2b#)) OR
 					(reg_q2417 AND symb_decoder(16#5b#)) OR
 					(reg_q2417 AND symb_decoder(16#f9#)) OR
 					(reg_q2417 AND symb_decoder(16#38#)) OR
 					(reg_q2417 AND symb_decoder(16#8a#)) OR
 					(reg_q2417 AND symb_decoder(16#4e#)) OR
 					(reg_q2417 AND symb_decoder(16#25#)) OR
 					(reg_q2417 AND symb_decoder(16#d6#)) OR
 					(reg_q2417 AND symb_decoder(16#ff#)) OR
 					(reg_q2417 AND symb_decoder(16#b1#)) OR
 					(reg_q2417 AND symb_decoder(16#d8#)) OR
 					(reg_q2417 AND symb_decoder(16#c7#)) OR
 					(reg_q2417 AND symb_decoder(16#45#)) OR
 					(reg_q2417 AND symb_decoder(16#9c#)) OR
 					(reg_q2417 AND symb_decoder(16#36#)) OR
 					(reg_q2417 AND symb_decoder(16#ce#)) OR
 					(reg_q2417 AND symb_decoder(16#7e#)) OR
 					(reg_q2417 AND symb_decoder(16#95#)) OR
 					(reg_q2417 AND symb_decoder(16#4b#)) OR
 					(reg_q2417 AND symb_decoder(16#fc#)) OR
 					(reg_q2417 AND symb_decoder(16#a0#)) OR
 					(reg_q2417 AND symb_decoder(16#67#)) OR
 					(reg_q2417 AND symb_decoder(16#d2#)) OR
 					(reg_q2417 AND symb_decoder(16#bc#)) OR
 					(reg_q2417 AND symb_decoder(16#51#)) OR
 					(reg_q2417 AND symb_decoder(16#4c#)) OR
 					(reg_q2417 AND symb_decoder(16#9e#)) OR
 					(reg_q2417 AND symb_decoder(16#52#)) OR
 					(reg_q2417 AND symb_decoder(16#00#)) OR
 					(reg_q2417 AND symb_decoder(16#20#)) OR
 					(reg_q2417 AND symb_decoder(16#3e#)) OR
 					(reg_q2417 AND symb_decoder(16#0b#)) OR
 					(reg_q2417 AND symb_decoder(16#f1#)) OR
 					(reg_q2417 AND symb_decoder(16#ae#)) OR
 					(reg_q2417 AND symb_decoder(16#df#)) OR
 					(reg_q2417 AND symb_decoder(16#72#)) OR
 					(reg_q2417 AND symb_decoder(16#53#)) OR
 					(reg_q2417 AND symb_decoder(16#27#)) OR
 					(reg_q2417 AND symb_decoder(16#fa#)) OR
 					(reg_q2417 AND symb_decoder(16#c5#)) OR
 					(reg_q2417 AND symb_decoder(16#eb#)) OR
 					(reg_q2417 AND symb_decoder(16#be#)) OR
 					(reg_q2417 AND symb_decoder(16#89#)) OR
 					(reg_q2417 AND symb_decoder(16#e1#)) OR
 					(reg_q2417 AND symb_decoder(16#7c#)) OR
 					(reg_q2417 AND symb_decoder(16#ba#)) OR
 					(reg_q2417 AND symb_decoder(16#55#)) OR
 					(reg_q2417 AND symb_decoder(16#31#)) OR
 					(reg_q2417 AND symb_decoder(16#5d#)) OR
 					(reg_q2417 AND symb_decoder(16#c4#)) OR
 					(reg_q2417 AND symb_decoder(16#3a#)) OR
 					(reg_q2417 AND symb_decoder(16#7f#)) OR
 					(reg_q2417 AND symb_decoder(16#32#)) OR
 					(reg_q2417 AND symb_decoder(16#49#)) OR
 					(reg_q2417 AND symb_decoder(16#79#)) OR
 					(reg_q2417 AND symb_decoder(16#13#)) OR
 					(reg_q2417 AND symb_decoder(16#6f#)) OR
 					(reg_q2417 AND symb_decoder(16#07#)) OR
 					(reg_q2417 AND symb_decoder(16#92#)) OR
 					(reg_q2417 AND symb_decoder(16#7d#)) OR
 					(reg_q2417 AND symb_decoder(16#59#)) OR
 					(reg_q2417 AND symb_decoder(16#50#)) OR
 					(reg_q2417 AND symb_decoder(16#73#)) OR
 					(reg_q2417 AND symb_decoder(16#2f#)) OR
 					(reg_q2417 AND symb_decoder(16#b4#)) OR
 					(reg_q2417 AND symb_decoder(16#48#)) OR
 					(reg_q2417 AND symb_decoder(16#08#)) OR
 					(reg_q2417 AND symb_decoder(16#d7#)) OR
 					(reg_q2417 AND symb_decoder(16#56#)) OR
 					(reg_q2417 AND symb_decoder(16#b5#)) OR
 					(reg_q2417 AND symb_decoder(16#1d#)) OR
 					(reg_q2417 AND symb_decoder(16#e9#)) OR
 					(reg_q2417 AND symb_decoder(16#41#)) OR
 					(reg_q2417 AND symb_decoder(16#28#)) OR
 					(reg_q2417 AND symb_decoder(16#2d#)) OR
 					(reg_q2417 AND symb_decoder(16#99#)) OR
 					(reg_q2417 AND symb_decoder(16#64#)) OR
 					(reg_q2417 AND symb_decoder(16#e3#)) OR
 					(reg_q2417 AND symb_decoder(16#63#)) OR
 					(reg_q2417 AND symb_decoder(16#f3#)) OR
 					(reg_q2417 AND symb_decoder(16#e5#)) OR
 					(reg_q2417 AND symb_decoder(16#03#)) OR
 					(reg_q2417 AND symb_decoder(16#68#)) OR
 					(reg_q2417 AND symb_decoder(16#bb#)) OR
 					(reg_q2417 AND symb_decoder(16#db#)) OR
 					(reg_q2417 AND symb_decoder(16#fb#)) OR
 					(reg_q2417 AND symb_decoder(16#f5#)) OR
 					(reg_q2417 AND symb_decoder(16#4f#)) OR
 					(reg_q2417 AND symb_decoder(16#84#)) OR
 					(reg_q2417 AND symb_decoder(16#01#)) OR
 					(reg_q2417 AND symb_decoder(16#0d#)) OR
 					(reg_q2417 AND symb_decoder(16#6b#)) OR
 					(reg_q2417 AND symb_decoder(16#f4#)) OR
 					(reg_q2417 AND symb_decoder(16#f8#)) OR
 					(reg_q2417 AND symb_decoder(16#05#)) OR
 					(reg_q2417 AND symb_decoder(16#70#)) OR
 					(reg_q2417 AND symb_decoder(16#2a#)) OR
 					(reg_q2417 AND symb_decoder(16#aa#)) OR
 					(reg_q2417 AND symb_decoder(16#33#)) OR
 					(reg_q2417 AND symb_decoder(16#cc#)) OR
 					(reg_q2417 AND symb_decoder(16#18#)) OR
 					(reg_q2417 AND symb_decoder(16#94#)) OR
 					(reg_q2417 AND symb_decoder(16#c0#)) OR
 					(reg_q2417 AND symb_decoder(16#75#)) OR
 					(reg_q2417 AND symb_decoder(16#30#)) OR
 					(reg_q2417 AND symb_decoder(16#a1#)) OR
 					(reg_q2417 AND symb_decoder(16#da#)) OR
 					(reg_q2417 AND symb_decoder(16#9a#)) OR
 					(reg_q2417 AND symb_decoder(16#69#)) OR
 					(reg_q2417 AND symb_decoder(16#66#)) OR
 					(reg_q2417 AND symb_decoder(16#ac#)) OR
 					(reg_q2417 AND symb_decoder(16#c3#)) OR
 					(reg_q2417 AND symb_decoder(16#81#)) OR
 					(reg_q2417 AND symb_decoder(16#04#)) OR
 					(reg_q2417 AND symb_decoder(16#dc#)) OR
 					(reg_q2417 AND symb_decoder(16#8e#)) OR
 					(reg_q2417 AND symb_decoder(16#ea#)) OR
 					(reg_q2417 AND symb_decoder(16#76#)) OR
 					(reg_q2417 AND symb_decoder(16#f7#)) OR
 					(reg_q2417 AND symb_decoder(16#43#)) OR
 					(reg_q2417 AND symb_decoder(16#8f#)) OR
 					(reg_q2417 AND symb_decoder(16#5a#)) OR
 					(reg_q2417 AND symb_decoder(16#fd#)) OR
 					(reg_q2417 AND symb_decoder(16#e6#)) OR
 					(reg_q2417 AND symb_decoder(16#cb#)) OR
 					(reg_q2417 AND symb_decoder(16#dd#)) OR
 					(reg_q2417 AND symb_decoder(16#c1#)) OR
 					(reg_q2417 AND symb_decoder(16#ef#)) OR
 					(reg_q2417 AND symb_decoder(16#e4#)) OR
 					(reg_q2417 AND symb_decoder(16#3f#)) OR
 					(reg_q2417 AND symb_decoder(16#23#)) OR
 					(reg_q2417 AND symb_decoder(16#f6#)) OR
 					(reg_q2417 AND symb_decoder(16#b6#)) OR
 					(reg_q2417 AND symb_decoder(16#1b#)) OR
 					(reg_q2417 AND symb_decoder(16#87#)) OR
 					(reg_q2417 AND symb_decoder(16#6a#)) OR
 					(reg_q2417 AND symb_decoder(16#5c#)) OR
 					(reg_q2417 AND symb_decoder(16#29#)) OR
 					(reg_q2417 AND symb_decoder(16#3b#)) OR
 					(reg_q2417 AND symb_decoder(16#5f#)) OR
 					(reg_q2417 AND symb_decoder(16#d9#)) OR
 					(reg_q2417 AND symb_decoder(16#6c#)) OR
 					(reg_q2417 AND symb_decoder(16#80#)) OR
 					(reg_q2417 AND symb_decoder(16#0c#)) OR
 					(reg_q2417 AND symb_decoder(16#ab#)) OR
 					(reg_q2417 AND symb_decoder(16#85#)) OR
 					(reg_q2417 AND symb_decoder(16#71#)) OR
 					(reg_q2417 AND symb_decoder(16#a2#)) OR
 					(reg_q2417 AND symb_decoder(16#fe#)) OR
 					(reg_q2417 AND symb_decoder(16#ee#)) OR
 					(reg_q2417 AND symb_decoder(16#a9#)) OR
 					(reg_q2417 AND symb_decoder(16#77#)) OR
 					(reg_q2417 AND symb_decoder(16#b3#)) OR
 					(reg_q2417 AND symb_decoder(16#2c#)) OR
 					(reg_q2417 AND symb_decoder(16#d1#)) OR
 					(reg_q2417 AND symb_decoder(16#d5#)) OR
 					(reg_q2417 AND symb_decoder(16#4a#)) OR
 					(reg_q2417 AND symb_decoder(16#b9#)) OR
 					(reg_q2417 AND symb_decoder(16#17#)) OR
 					(reg_q2417 AND symb_decoder(16#24#)) OR
 					(reg_q2417 AND symb_decoder(16#b7#));
reg_q2417_init <= '0' ;
	p_reg_q2417: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2417 <= reg_q2417_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2417 <= reg_q2417_init;
        else
          reg_q2417 <= reg_q2417_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q99_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q99 AND symb_decoder(16#2a#)) OR
 					(reg_q99 AND symb_decoder(16#05#)) OR
 					(reg_q99 AND symb_decoder(16#ed#)) OR
 					(reg_q99 AND symb_decoder(16#ce#)) OR
 					(reg_q99 AND symb_decoder(16#56#)) OR
 					(reg_q99 AND symb_decoder(16#03#)) OR
 					(reg_q99 AND symb_decoder(16#1f#)) OR
 					(reg_q99 AND symb_decoder(16#cb#)) OR
 					(reg_q99 AND symb_decoder(16#af#)) OR
 					(reg_q99 AND symb_decoder(16#4d#)) OR
 					(reg_q99 AND symb_decoder(16#27#)) OR
 					(reg_q99 AND symb_decoder(16#28#)) OR
 					(reg_q99 AND symb_decoder(16#d8#)) OR
 					(reg_q99 AND symb_decoder(16#34#)) OR
 					(reg_q99 AND symb_decoder(16#a4#)) OR
 					(reg_q99 AND symb_decoder(16#59#)) OR
 					(reg_q99 AND symb_decoder(16#f5#)) OR
 					(reg_q99 AND symb_decoder(16#8c#)) OR
 					(reg_q99 AND symb_decoder(16#fb#)) OR
 					(reg_q99 AND symb_decoder(16#e5#)) OR
 					(reg_q99 AND symb_decoder(16#eb#)) OR
 					(reg_q99 AND symb_decoder(16#50#)) OR
 					(reg_q99 AND symb_decoder(16#f6#)) OR
 					(reg_q99 AND symb_decoder(16#a9#)) OR
 					(reg_q99 AND symb_decoder(16#30#)) OR
 					(reg_q99 AND symb_decoder(16#54#)) OR
 					(reg_q99 AND symb_decoder(16#84#)) OR
 					(reg_q99 AND symb_decoder(16#9d#)) OR
 					(reg_q99 AND symb_decoder(16#7e#)) OR
 					(reg_q99 AND symb_decoder(16#6f#)) OR
 					(reg_q99 AND symb_decoder(16#f3#)) OR
 					(reg_q99 AND symb_decoder(16#68#)) OR
 					(reg_q99 AND symb_decoder(16#98#)) OR
 					(reg_q99 AND symb_decoder(16#be#)) OR
 					(reg_q99 AND symb_decoder(16#16#)) OR
 					(reg_q99 AND symb_decoder(16#9c#)) OR
 					(reg_q99 AND symb_decoder(16#18#)) OR
 					(reg_q99 AND symb_decoder(16#7b#)) OR
 					(reg_q99 AND symb_decoder(16#75#)) OR
 					(reg_q99 AND symb_decoder(16#e1#)) OR
 					(reg_q99 AND symb_decoder(16#d5#)) OR
 					(reg_q99 AND symb_decoder(16#db#)) OR
 					(reg_q99 AND symb_decoder(16#3c#)) OR
 					(reg_q99 AND symb_decoder(16#42#)) OR
 					(reg_q99 AND symb_decoder(16#bd#)) OR
 					(reg_q99 AND symb_decoder(16#0f#)) OR
 					(reg_q99 AND symb_decoder(16#6e#)) OR
 					(reg_q99 AND symb_decoder(16#f4#)) OR
 					(reg_q99 AND symb_decoder(16#8a#)) OR
 					(reg_q99 AND symb_decoder(16#a2#)) OR
 					(reg_q99 AND symb_decoder(16#c7#)) OR
 					(reg_q99 AND symb_decoder(16#fe#)) OR
 					(reg_q99 AND symb_decoder(16#c8#)) OR
 					(reg_q99 AND symb_decoder(16#7f#)) OR
 					(reg_q99 AND symb_decoder(16#48#)) OR
 					(reg_q99 AND symb_decoder(16#d9#)) OR
 					(reg_q99 AND symb_decoder(16#51#)) OR
 					(reg_q99 AND symb_decoder(16#49#)) OR
 					(reg_q99 AND symb_decoder(16#01#)) OR
 					(reg_q99 AND symb_decoder(16#89#)) OR
 					(reg_q99 AND symb_decoder(16#76#)) OR
 					(reg_q99 AND symb_decoder(16#5a#)) OR
 					(reg_q99 AND symb_decoder(16#55#)) OR
 					(reg_q99 AND symb_decoder(16#66#)) OR
 					(reg_q99 AND symb_decoder(16#a6#)) OR
 					(reg_q99 AND symb_decoder(16#21#)) OR
 					(reg_q99 AND symb_decoder(16#38#)) OR
 					(reg_q99 AND symb_decoder(16#2c#)) OR
 					(reg_q99 AND symb_decoder(16#3f#)) OR
 					(reg_q99 AND symb_decoder(16#62#)) OR
 					(reg_q99 AND symb_decoder(16#97#)) OR
 					(reg_q99 AND symb_decoder(16#02#)) OR
 					(reg_q99 AND symb_decoder(16#46#)) OR
 					(reg_q99 AND symb_decoder(16#2d#)) OR
 					(reg_q99 AND symb_decoder(16#0d#)) OR
 					(reg_q99 AND symb_decoder(16#c9#)) OR
 					(reg_q99 AND symb_decoder(16#87#)) OR
 					(reg_q99 AND symb_decoder(16#20#)) OR
 					(reg_q99 AND symb_decoder(16#6c#)) OR
 					(reg_q99 AND symb_decoder(16#22#)) OR
 					(reg_q99 AND symb_decoder(16#c2#)) OR
 					(reg_q99 AND symb_decoder(16#08#)) OR
 					(reg_q99 AND symb_decoder(16#e3#)) OR
 					(reg_q99 AND symb_decoder(16#c4#)) OR
 					(reg_q99 AND symb_decoder(16#d2#)) OR
 					(reg_q99 AND symb_decoder(16#4b#)) OR
 					(reg_q99 AND symb_decoder(16#e6#)) OR
 					(reg_q99 AND symb_decoder(16#10#)) OR
 					(reg_q99 AND symb_decoder(16#f2#)) OR
 					(reg_q99 AND symb_decoder(16#83#)) OR
 					(reg_q99 AND symb_decoder(16#a7#)) OR
 					(reg_q99 AND symb_decoder(16#3e#)) OR
 					(reg_q99 AND symb_decoder(16#63#)) OR
 					(reg_q99 AND symb_decoder(16#44#)) OR
 					(reg_q99 AND symb_decoder(16#d3#)) OR
 					(reg_q99 AND symb_decoder(16#f9#)) OR
 					(reg_q99 AND symb_decoder(16#73#)) OR
 					(reg_q99 AND symb_decoder(16#0b#)) OR
 					(reg_q99 AND symb_decoder(16#7a#)) OR
 					(reg_q99 AND symb_decoder(16#fc#)) OR
 					(reg_q99 AND symb_decoder(16#aa#)) OR
 					(reg_q99 AND symb_decoder(16#80#)) OR
 					(reg_q99 AND symb_decoder(16#c6#)) OR
 					(reg_q99 AND symb_decoder(16#25#)) OR
 					(reg_q99 AND symb_decoder(16#ac#)) OR
 					(reg_q99 AND symb_decoder(16#40#)) OR
 					(reg_q99 AND symb_decoder(16#b6#)) OR
 					(reg_q99 AND symb_decoder(16#60#)) OR
 					(reg_q99 AND symb_decoder(16#fd#)) OR
 					(reg_q99 AND symb_decoder(16#f1#)) OR
 					(reg_q99 AND symb_decoder(16#b7#)) OR
 					(reg_q99 AND symb_decoder(16#36#)) OR
 					(reg_q99 AND symb_decoder(16#f0#)) OR
 					(reg_q99 AND symb_decoder(16#69#)) OR
 					(reg_q99 AND symb_decoder(16#bb#)) OR
 					(reg_q99 AND symb_decoder(16#2f#)) OR
 					(reg_q99 AND symb_decoder(16#96#)) OR
 					(reg_q99 AND symb_decoder(16#00#)) OR
 					(reg_q99 AND symb_decoder(16#b5#)) OR
 					(reg_q99 AND symb_decoder(16#ba#)) OR
 					(reg_q99 AND symb_decoder(16#ee#)) OR
 					(reg_q99 AND symb_decoder(16#95#)) OR
 					(reg_q99 AND symb_decoder(16#b4#)) OR
 					(reg_q99 AND symb_decoder(16#74#)) OR
 					(reg_q99 AND symb_decoder(16#17#)) OR
 					(reg_q99 AND symb_decoder(16#15#)) OR
 					(reg_q99 AND symb_decoder(16#52#)) OR
 					(reg_q99 AND symb_decoder(16#8e#)) OR
 					(reg_q99 AND symb_decoder(16#32#)) OR
 					(reg_q99 AND symb_decoder(16#09#)) OR
 					(reg_q99 AND symb_decoder(16#43#)) OR
 					(reg_q99 AND symb_decoder(16#e9#)) OR
 					(reg_q99 AND symb_decoder(16#04#)) OR
 					(reg_q99 AND symb_decoder(16#06#)) OR
 					(reg_q99 AND symb_decoder(16#b0#)) OR
 					(reg_q99 AND symb_decoder(16#e7#)) OR
 					(reg_q99 AND symb_decoder(16#b8#)) OR
 					(reg_q99 AND symb_decoder(16#cc#)) OR
 					(reg_q99 AND symb_decoder(16#07#)) OR
 					(reg_q99 AND symb_decoder(16#11#)) OR
 					(reg_q99 AND symb_decoder(16#f7#)) OR
 					(reg_q99 AND symb_decoder(16#c3#)) OR
 					(reg_q99 AND symb_decoder(16#bc#)) OR
 					(reg_q99 AND symb_decoder(16#d1#)) OR
 					(reg_q99 AND symb_decoder(16#bf#)) OR
 					(reg_q99 AND symb_decoder(16#5b#)) OR
 					(reg_q99 AND symb_decoder(16#8f#)) OR
 					(reg_q99 AND symb_decoder(16#ad#)) OR
 					(reg_q99 AND symb_decoder(16#da#)) OR
 					(reg_q99 AND symb_decoder(16#0a#)) OR
 					(reg_q99 AND symb_decoder(16#99#)) OR
 					(reg_q99 AND symb_decoder(16#4f#)) OR
 					(reg_q99 AND symb_decoder(16#e8#)) OR
 					(reg_q99 AND symb_decoder(16#9e#)) OR
 					(reg_q99 AND symb_decoder(16#5e#)) OR
 					(reg_q99 AND symb_decoder(16#1b#)) OR
 					(reg_q99 AND symb_decoder(16#ae#)) OR
 					(reg_q99 AND symb_decoder(16#d4#)) OR
 					(reg_q99 AND symb_decoder(16#65#)) OR
 					(reg_q99 AND symb_decoder(16#79#)) OR
 					(reg_q99 AND symb_decoder(16#e0#)) OR
 					(reg_q99 AND symb_decoder(16#e2#)) OR
 					(reg_q99 AND symb_decoder(16#1d#)) OR
 					(reg_q99 AND symb_decoder(16#64#)) OR
 					(reg_q99 AND symb_decoder(16#58#)) OR
 					(reg_q99 AND symb_decoder(16#cf#)) OR
 					(reg_q99 AND symb_decoder(16#ea#)) OR
 					(reg_q99 AND symb_decoder(16#81#)) OR
 					(reg_q99 AND symb_decoder(16#71#)) OR
 					(reg_q99 AND symb_decoder(16#9a#)) OR
 					(reg_q99 AND symb_decoder(16#85#)) OR
 					(reg_q99 AND symb_decoder(16#0e#)) OR
 					(reg_q99 AND symb_decoder(16#c0#)) OR
 					(reg_q99 AND symb_decoder(16#31#)) OR
 					(reg_q99 AND symb_decoder(16#57#)) OR
 					(reg_q99 AND symb_decoder(16#8b#)) OR
 					(reg_q99 AND symb_decoder(16#47#)) OR
 					(reg_q99 AND symb_decoder(16#a1#)) OR
 					(reg_q99 AND symb_decoder(16#94#)) OR
 					(reg_q99 AND symb_decoder(16#6d#)) OR
 					(reg_q99 AND symb_decoder(16#7d#)) OR
 					(reg_q99 AND symb_decoder(16#77#)) OR
 					(reg_q99 AND symb_decoder(16#5d#)) OR
 					(reg_q99 AND symb_decoder(16#93#)) OR
 					(reg_q99 AND symb_decoder(16#de#)) OR
 					(reg_q99 AND symb_decoder(16#90#)) OR
 					(reg_q99 AND symb_decoder(16#ab#)) OR
 					(reg_q99 AND symb_decoder(16#f8#)) OR
 					(reg_q99 AND symb_decoder(16#2e#)) OR
 					(reg_q99 AND symb_decoder(16#a5#)) OR
 					(reg_q99 AND symb_decoder(16#cd#)) OR
 					(reg_q99 AND symb_decoder(16#d7#)) OR
 					(reg_q99 AND symb_decoder(16#39#)) OR
 					(reg_q99 AND symb_decoder(16#ef#)) OR
 					(reg_q99 AND symb_decoder(16#86#)) OR
 					(reg_q99 AND symb_decoder(16#ff#)) OR
 					(reg_q99 AND symb_decoder(16#c5#)) OR
 					(reg_q99 AND symb_decoder(16#92#)) OR
 					(reg_q99 AND symb_decoder(16#dc#)) OR
 					(reg_q99 AND symb_decoder(16#1c#)) OR
 					(reg_q99 AND symb_decoder(16#0c#)) OR
 					(reg_q99 AND symb_decoder(16#df#)) OR
 					(reg_q99 AND symb_decoder(16#4c#)) OR
 					(reg_q99 AND symb_decoder(16#9b#)) OR
 					(reg_q99 AND symb_decoder(16#b3#)) OR
 					(reg_q99 AND symb_decoder(16#23#)) OR
 					(reg_q99 AND symb_decoder(16#3b#)) OR
 					(reg_q99 AND symb_decoder(16#5f#)) OR
 					(reg_q99 AND symb_decoder(16#1e#)) OR
 					(reg_q99 AND symb_decoder(16#13#)) OR
 					(reg_q99 AND symb_decoder(16#4a#)) OR
 					(reg_q99 AND symb_decoder(16#24#)) OR
 					(reg_q99 AND symb_decoder(16#12#)) OR
 					(reg_q99 AND symb_decoder(16#ca#)) OR
 					(reg_q99 AND symb_decoder(16#78#)) OR
 					(reg_q99 AND symb_decoder(16#ec#)) OR
 					(reg_q99 AND symb_decoder(16#61#)) OR
 					(reg_q99 AND symb_decoder(16#45#)) OR
 					(reg_q99 AND symb_decoder(16#41#)) OR
 					(reg_q99 AND symb_decoder(16#5c#)) OR
 					(reg_q99 AND symb_decoder(16#6b#)) OR
 					(reg_q99 AND symb_decoder(16#1a#)) OR
 					(reg_q99 AND symb_decoder(16#29#)) OR
 					(reg_q99 AND symb_decoder(16#2b#)) OR
 					(reg_q99 AND symb_decoder(16#c1#)) OR
 					(reg_q99 AND symb_decoder(16#8d#)) OR
 					(reg_q99 AND symb_decoder(16#e4#)) OR
 					(reg_q99 AND symb_decoder(16#b9#)) OR
 					(reg_q99 AND symb_decoder(16#82#)) OR
 					(reg_q99 AND symb_decoder(16#91#)) OR
 					(reg_q99 AND symb_decoder(16#a0#)) OR
 					(reg_q99 AND symb_decoder(16#4e#)) OR
 					(reg_q99 AND symb_decoder(16#3d#)) OR
 					(reg_q99 AND symb_decoder(16#b1#)) OR
 					(reg_q99 AND symb_decoder(16#72#)) OR
 					(reg_q99 AND symb_decoder(16#dd#)) OR
 					(reg_q99 AND symb_decoder(16#26#)) OR
 					(reg_q99 AND symb_decoder(16#6a#)) OR
 					(reg_q99 AND symb_decoder(16#a8#)) OR
 					(reg_q99 AND symb_decoder(16#7c#)) OR
 					(reg_q99 AND symb_decoder(16#fa#)) OR
 					(reg_q99 AND symb_decoder(16#70#)) OR
 					(reg_q99 AND symb_decoder(16#67#)) OR
 					(reg_q99 AND symb_decoder(16#a3#)) OR
 					(reg_q99 AND symb_decoder(16#35#)) OR
 					(reg_q99 AND symb_decoder(16#9f#)) OR
 					(reg_q99 AND symb_decoder(16#3a#)) OR
 					(reg_q99 AND symb_decoder(16#b2#)) OR
 					(reg_q99 AND symb_decoder(16#19#)) OR
 					(reg_q99 AND symb_decoder(16#d0#)) OR
 					(reg_q99 AND symb_decoder(16#14#)) OR
 					(reg_q99 AND symb_decoder(16#88#)) OR
 					(reg_q99 AND symb_decoder(16#d6#)) OR
 					(reg_q99 AND symb_decoder(16#53#)) OR
 					(reg_q99 AND symb_decoder(16#33#)) OR
 					(reg_q99 AND symb_decoder(16#37#));
reg_q99_init <= '0' ;
	p_reg_q99: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q99 <= reg_q99_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q99 <= reg_q99_init;
        else
          reg_q99 <= reg_q99_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph33

reg_q395_in <= (reg_q395 AND symb_decoder(16#6d#)) OR
 					(reg_q395 AND symb_decoder(16#cc#)) OR
 					(reg_q395 AND symb_decoder(16#95#)) OR
 					(reg_q395 AND symb_decoder(16#8d#)) OR
 					(reg_q395 AND symb_decoder(16#49#)) OR
 					(reg_q395 AND symb_decoder(16#c9#)) OR
 					(reg_q395 AND symb_decoder(16#af#)) OR
 					(reg_q395 AND symb_decoder(16#b3#)) OR
 					(reg_q395 AND symb_decoder(16#51#)) OR
 					(reg_q395 AND symb_decoder(16#47#)) OR
 					(reg_q395 AND symb_decoder(16#41#)) OR
 					(reg_q395 AND symb_decoder(16#88#)) OR
 					(reg_q395 AND symb_decoder(16#42#)) OR
 					(reg_q395 AND symb_decoder(16#d5#)) OR
 					(reg_q395 AND symb_decoder(16#fa#)) OR
 					(reg_q395 AND symb_decoder(16#6a#)) OR
 					(reg_q395 AND symb_decoder(16#33#)) OR
 					(reg_q395 AND symb_decoder(16#96#)) OR
 					(reg_q395 AND symb_decoder(16#38#)) OR
 					(reg_q395 AND symb_decoder(16#b8#)) OR
 					(reg_q395 AND symb_decoder(16#ae#)) OR
 					(reg_q395 AND symb_decoder(16#0f#)) OR
 					(reg_q395 AND symb_decoder(16#5c#)) OR
 					(reg_q395 AND symb_decoder(16#06#)) OR
 					(reg_q395 AND symb_decoder(16#c1#)) OR
 					(reg_q395 AND symb_decoder(16#36#)) OR
 					(reg_q395 AND symb_decoder(16#8c#)) OR
 					(reg_q395 AND symb_decoder(16#9d#)) OR
 					(reg_q395 AND symb_decoder(16#98#)) OR
 					(reg_q395 AND symb_decoder(16#b4#)) OR
 					(reg_q395 AND symb_decoder(16#ab#)) OR
 					(reg_q395 AND symb_decoder(16#3e#)) OR
 					(reg_q395 AND symb_decoder(16#83#)) OR
 					(reg_q395 AND symb_decoder(16#99#)) OR
 					(reg_q395 AND symb_decoder(16#a5#)) OR
 					(reg_q395 AND symb_decoder(16#60#)) OR
 					(reg_q395 AND symb_decoder(16#ca#)) OR
 					(reg_q395 AND symb_decoder(16#44#)) OR
 					(reg_q395 AND symb_decoder(16#64#)) OR
 					(reg_q395 AND symb_decoder(16#b5#)) OR
 					(reg_q395 AND symb_decoder(16#f0#)) OR
 					(reg_q395 AND symb_decoder(16#2c#)) OR
 					(reg_q395 AND symb_decoder(16#7e#)) OR
 					(reg_q395 AND symb_decoder(16#37#)) OR
 					(reg_q395 AND symb_decoder(16#f2#)) OR
 					(reg_q395 AND symb_decoder(16#d3#)) OR
 					(reg_q395 AND symb_decoder(16#3a#)) OR
 					(reg_q395 AND symb_decoder(16#63#)) OR
 					(reg_q395 AND symb_decoder(16#d4#)) OR
 					(reg_q395 AND symb_decoder(16#03#)) OR
 					(reg_q395 AND symb_decoder(16#4e#)) OR
 					(reg_q395 AND symb_decoder(16#a8#)) OR
 					(reg_q395 AND symb_decoder(16#a6#)) OR
 					(reg_q395 AND symb_decoder(16#ea#)) OR
 					(reg_q395 AND symb_decoder(16#e7#)) OR
 					(reg_q395 AND symb_decoder(16#1d#)) OR
 					(reg_q395 AND symb_decoder(16#69#)) OR
 					(reg_q395 AND symb_decoder(16#21#)) OR
 					(reg_q395 AND symb_decoder(16#cd#)) OR
 					(reg_q395 AND symb_decoder(16#02#)) OR
 					(reg_q395 AND symb_decoder(16#93#)) OR
 					(reg_q395 AND symb_decoder(16#68#)) OR
 					(reg_q395 AND symb_decoder(16#54#)) OR
 					(reg_q395 AND symb_decoder(16#58#)) OR
 					(reg_q395 AND symb_decoder(16#81#)) OR
 					(reg_q395 AND symb_decoder(16#bd#)) OR
 					(reg_q395 AND symb_decoder(16#01#)) OR
 					(reg_q395 AND symb_decoder(16#76#)) OR
 					(reg_q395 AND symb_decoder(16#2a#)) OR
 					(reg_q395 AND symb_decoder(16#cf#)) OR
 					(reg_q395 AND symb_decoder(16#e5#)) OR
 					(reg_q395 AND symb_decoder(16#ff#)) OR
 					(reg_q395 AND symb_decoder(16#62#)) OR
 					(reg_q395 AND symb_decoder(16#84#)) OR
 					(reg_q395 AND symb_decoder(16#9e#)) OR
 					(reg_q395 AND symb_decoder(16#50#)) OR
 					(reg_q395 AND symb_decoder(16#26#)) OR
 					(reg_q395 AND symb_decoder(16#15#)) OR
 					(reg_q395 AND symb_decoder(16#e8#)) OR
 					(reg_q395 AND symb_decoder(16#32#)) OR
 					(reg_q395 AND symb_decoder(16#91#)) OR
 					(reg_q395 AND symb_decoder(16#3b#)) OR
 					(reg_q395 AND symb_decoder(16#10#)) OR
 					(reg_q395 AND symb_decoder(16#0b#)) OR
 					(reg_q395 AND symb_decoder(16#39#)) OR
 					(reg_q395 AND symb_decoder(16#5b#)) OR
 					(reg_q395 AND symb_decoder(16#9f#)) OR
 					(reg_q395 AND symb_decoder(16#ee#)) OR
 					(reg_q395 AND symb_decoder(16#57#)) OR
 					(reg_q395 AND symb_decoder(16#ad#)) OR
 					(reg_q395 AND symb_decoder(16#f6#)) OR
 					(reg_q395 AND symb_decoder(16#2d#)) OR
 					(reg_q395 AND symb_decoder(16#a4#)) OR
 					(reg_q395 AND symb_decoder(16#09#)) OR
 					(reg_q395 AND symb_decoder(16#7f#)) OR
 					(reg_q395 AND symb_decoder(16#f9#)) OR
 					(reg_q395 AND symb_decoder(16#24#)) OR
 					(reg_q395 AND symb_decoder(16#c8#)) OR
 					(reg_q395 AND symb_decoder(16#25#)) OR
 					(reg_q395 AND symb_decoder(16#79#)) OR
 					(reg_q395 AND symb_decoder(16#0e#)) OR
 					(reg_q395 AND symb_decoder(16#d7#)) OR
 					(reg_q395 AND symb_decoder(16#b7#)) OR
 					(reg_q395 AND symb_decoder(16#b0#)) OR
 					(reg_q395 AND symb_decoder(16#04#)) OR
 					(reg_q395 AND symb_decoder(16#df#)) OR
 					(reg_q395 AND symb_decoder(16#d0#)) OR
 					(reg_q395 AND symb_decoder(16#18#)) OR
 					(reg_q395 AND symb_decoder(16#ba#)) OR
 					(reg_q395 AND symb_decoder(16#59#)) OR
 					(reg_q395 AND symb_decoder(16#e0#)) OR
 					(reg_q395 AND symb_decoder(16#97#)) OR
 					(reg_q395 AND symb_decoder(16#08#)) OR
 					(reg_q395 AND symb_decoder(16#8b#)) OR
 					(reg_q395 AND symb_decoder(16#4c#)) OR
 					(reg_q395 AND symb_decoder(16#ac#)) OR
 					(reg_q395 AND symb_decoder(16#31#)) OR
 					(reg_q395 AND symb_decoder(16#14#)) OR
 					(reg_q395 AND symb_decoder(16#13#)) OR
 					(reg_q395 AND symb_decoder(16#bb#)) OR
 					(reg_q395 AND symb_decoder(16#17#)) OR
 					(reg_q395 AND symb_decoder(16#fb#)) OR
 					(reg_q395 AND symb_decoder(16#16#)) OR
 					(reg_q395 AND symb_decoder(16#ce#)) OR
 					(reg_q395 AND symb_decoder(16#e6#)) OR
 					(reg_q395 AND symb_decoder(16#d9#)) OR
 					(reg_q395 AND symb_decoder(16#5d#)) OR
 					(reg_q395 AND symb_decoder(16#56#)) OR
 					(reg_q395 AND symb_decoder(16#65#)) OR
 					(reg_q395 AND symb_decoder(16#92#)) OR
 					(reg_q395 AND symb_decoder(16#85#)) OR
 					(reg_q395 AND symb_decoder(16#0c#)) OR
 					(reg_q395 AND symb_decoder(16#f3#)) OR
 					(reg_q395 AND symb_decoder(16#27#)) OR
 					(reg_q395 AND symb_decoder(16#89#)) OR
 					(reg_q395 AND symb_decoder(16#3d#)) OR
 					(reg_q395 AND symb_decoder(16#dd#)) OR
 					(reg_q395 AND symb_decoder(16#8e#)) OR
 					(reg_q395 AND symb_decoder(16#9a#)) OR
 					(reg_q395 AND symb_decoder(16#07#)) OR
 					(reg_q395 AND symb_decoder(16#19#)) OR
 					(reg_q395 AND symb_decoder(16#f1#)) OR
 					(reg_q395 AND symb_decoder(16#6c#)) OR
 					(reg_q395 AND symb_decoder(16#5e#)) OR
 					(reg_q395 AND symb_decoder(16#a3#)) OR
 					(reg_q395 AND symb_decoder(16#6f#)) OR
 					(reg_q395 AND symb_decoder(16#d1#)) OR
 					(reg_q395 AND symb_decoder(16#a7#)) OR
 					(reg_q395 AND symb_decoder(16#c5#)) OR
 					(reg_q395 AND symb_decoder(16#4b#)) OR
 					(reg_q395 AND symb_decoder(16#7c#)) OR
 					(reg_q395 AND symb_decoder(16#f7#)) OR
 					(reg_q395 AND symb_decoder(16#35#)) OR
 					(reg_q395 AND symb_decoder(16#9c#)) OR
 					(reg_q395 AND symb_decoder(16#2b#)) OR
 					(reg_q395 AND symb_decoder(16#1f#)) OR
 					(reg_q395 AND symb_decoder(16#6b#)) OR
 					(reg_q395 AND symb_decoder(16#bc#)) OR
 					(reg_q395 AND symb_decoder(16#7d#)) OR
 					(reg_q395 AND symb_decoder(16#1e#)) OR
 					(reg_q395 AND symb_decoder(16#94#)) OR
 					(reg_q395 AND symb_decoder(16#22#)) OR
 					(reg_q395 AND symb_decoder(16#30#)) OR
 					(reg_q395 AND symb_decoder(16#72#)) OR
 					(reg_q395 AND symb_decoder(16#29#)) OR
 					(reg_q395 AND symb_decoder(16#67#)) OR
 					(reg_q395 AND symb_decoder(16#74#)) OR
 					(reg_q395 AND symb_decoder(16#cb#)) OR
 					(reg_q395 AND symb_decoder(16#b6#)) OR
 					(reg_q395 AND symb_decoder(16#3f#)) OR
 					(reg_q395 AND symb_decoder(16#1b#)) OR
 					(reg_q395 AND symb_decoder(16#b9#)) OR
 					(reg_q395 AND symb_decoder(16#e9#)) OR
 					(reg_q395 AND symb_decoder(16#f8#)) OR
 					(reg_q395 AND symb_decoder(16#b1#)) OR
 					(reg_q395 AND symb_decoder(16#c4#)) OR
 					(reg_q395 AND symb_decoder(16#52#)) OR
 					(reg_q395 AND symb_decoder(16#de#)) OR
 					(reg_q395 AND symb_decoder(16#2f#)) OR
 					(reg_q395 AND symb_decoder(16#be#)) OR
 					(reg_q395 AND symb_decoder(16#9b#)) OR
 					(reg_q395 AND symb_decoder(16#43#)) OR
 					(reg_q395 AND symb_decoder(16#b2#)) OR
 					(reg_q395 AND symb_decoder(16#70#)) OR
 					(reg_q395 AND symb_decoder(16#75#)) OR
 					(reg_q395 AND symb_decoder(16#40#)) OR
 					(reg_q395 AND symb_decoder(16#a2#)) OR
 					(reg_q395 AND symb_decoder(16#71#)) OR
 					(reg_q395 AND symb_decoder(16#eb#)) OR
 					(reg_q395 AND symb_decoder(16#f5#)) OR
 					(reg_q395 AND symb_decoder(16#d2#)) OR
 					(reg_q395 AND symb_decoder(16#5a#)) OR
 					(reg_q395 AND symb_decoder(16#fe#)) OR
 					(reg_q395 AND symb_decoder(16#c3#)) OR
 					(reg_q395 AND symb_decoder(16#8f#)) OR
 					(reg_q395 AND symb_decoder(16#66#)) OR
 					(reg_q395 AND symb_decoder(16#aa#)) OR
 					(reg_q395 AND symb_decoder(16#7a#)) OR
 					(reg_q395 AND symb_decoder(16#87#)) OR
 					(reg_q395 AND symb_decoder(16#e4#)) OR
 					(reg_q395 AND symb_decoder(16#e1#)) OR
 					(reg_q395 AND symb_decoder(16#3c#)) OR
 					(reg_q395 AND symb_decoder(16#5f#)) OR
 					(reg_q395 AND symb_decoder(16#a0#)) OR
 					(reg_q395 AND symb_decoder(16#23#)) OR
 					(reg_q395 AND symb_decoder(16#1a#)) OR
 					(reg_q395 AND symb_decoder(16#4a#)) OR
 					(reg_q395 AND symb_decoder(16#46#)) OR
 					(reg_q395 AND symb_decoder(16#6e#)) OR
 					(reg_q395 AND symb_decoder(16#34#)) OR
 					(reg_q395 AND symb_decoder(16#48#)) OR
 					(reg_q395 AND symb_decoder(16#2e#)) OR
 					(reg_q395 AND symb_decoder(16#45#)) OR
 					(reg_q395 AND symb_decoder(16#fc#)) OR
 					(reg_q395 AND symb_decoder(16#73#)) OR
 					(reg_q395 AND symb_decoder(16#77#)) OR
 					(reg_q395 AND symb_decoder(16#ef#)) OR
 					(reg_q395 AND symb_decoder(16#12#)) OR
 					(reg_q395 AND symb_decoder(16#a1#)) OR
 					(reg_q395 AND symb_decoder(16#90#)) OR
 					(reg_q395 AND symb_decoder(16#28#)) OR
 					(reg_q395 AND symb_decoder(16#4d#)) OR
 					(reg_q395 AND symb_decoder(16#00#)) OR
 					(reg_q395 AND symb_decoder(16#e2#)) OR
 					(reg_q395 AND symb_decoder(16#c7#)) OR
 					(reg_q395 AND symb_decoder(16#a9#)) OR
 					(reg_q395 AND symb_decoder(16#da#)) OR
 					(reg_q395 AND symb_decoder(16#c0#)) OR
 					(reg_q395 AND symb_decoder(16#55#)) OR
 					(reg_q395 AND symb_decoder(16#bf#)) OR
 					(reg_q395 AND symb_decoder(16#f4#)) OR
 					(reg_q395 AND symb_decoder(16#c2#)) OR
 					(reg_q395 AND symb_decoder(16#7b#)) OR
 					(reg_q395 AND symb_decoder(16#86#)) OR
 					(reg_q395 AND symb_decoder(16#20#)) OR
 					(reg_q395 AND symb_decoder(16#05#)) OR
 					(reg_q395 AND symb_decoder(16#78#)) OR
 					(reg_q395 AND symb_decoder(16#c6#)) OR
 					(reg_q395 AND symb_decoder(16#d6#)) OR
 					(reg_q395 AND symb_decoder(16#db#)) OR
 					(reg_q395 AND symb_decoder(16#d8#)) OR
 					(reg_q395 AND symb_decoder(16#1c#)) OR
 					(reg_q395 AND symb_decoder(16#e3#)) OR
 					(reg_q395 AND symb_decoder(16#53#)) OR
 					(reg_q395 AND symb_decoder(16#61#)) OR
 					(reg_q395 AND symb_decoder(16#fd#)) OR
 					(reg_q395 AND symb_decoder(16#82#)) OR
 					(reg_q395 AND symb_decoder(16#dc#)) OR
 					(reg_q395 AND symb_decoder(16#ed#)) OR
 					(reg_q395 AND symb_decoder(16#8a#)) OR
 					(reg_q395 AND symb_decoder(16#4f#)) OR
 					(reg_q395 AND symb_decoder(16#ec#)) OR
 					(reg_q395 AND symb_decoder(16#80#)) OR
 					(reg_q395 AND symb_decoder(16#11#)) OR
 					(reg_q369 AND symb_decoder(16#d7#)) OR
 					(reg_q369 AND symb_decoder(16#c1#)) OR
 					(reg_q369 AND symb_decoder(16#a3#)) OR
 					(reg_q369 AND symb_decoder(16#91#)) OR
 					(reg_q369 AND symb_decoder(16#a8#)) OR
 					(reg_q369 AND symb_decoder(16#df#)) OR
 					(reg_q369 AND symb_decoder(16#1e#)) OR
 					(reg_q369 AND symb_decoder(16#69#)) OR
 					(reg_q369 AND symb_decoder(16#b4#)) OR
 					(reg_q369 AND symb_decoder(16#27#)) OR
 					(reg_q369 AND symb_decoder(16#33#)) OR
 					(reg_q369 AND symb_decoder(16#10#)) OR
 					(reg_q369 AND symb_decoder(16#19#)) OR
 					(reg_q369 AND symb_decoder(16#e3#)) OR
 					(reg_q369 AND symb_decoder(16#78#)) OR
 					(reg_q369 AND symb_decoder(16#5b#)) OR
 					(reg_q369 AND symb_decoder(16#75#)) OR
 					(reg_q369 AND symb_decoder(16#31#)) OR
 					(reg_q369 AND symb_decoder(16#4e#)) OR
 					(reg_q369 AND symb_decoder(16#39#)) OR
 					(reg_q369 AND symb_decoder(16#1c#)) OR
 					(reg_q369 AND symb_decoder(16#8f#)) OR
 					(reg_q369 AND symb_decoder(16#3e#)) OR
 					(reg_q369 AND symb_decoder(16#47#)) OR
 					(reg_q369 AND symb_decoder(16#77#)) OR
 					(reg_q369 AND symb_decoder(16#57#)) OR
 					(reg_q369 AND symb_decoder(16#9f#)) OR
 					(reg_q369 AND symb_decoder(16#96#)) OR
 					(reg_q369 AND symb_decoder(16#97#)) OR
 					(reg_q369 AND symb_decoder(16#06#)) OR
 					(reg_q369 AND symb_decoder(16#3c#)) OR
 					(reg_q369 AND symb_decoder(16#11#)) OR
 					(reg_q369 AND symb_decoder(16#62#)) OR
 					(reg_q369 AND symb_decoder(16#e0#)) OR
 					(reg_q369 AND symb_decoder(16#c7#)) OR
 					(reg_q369 AND symb_decoder(16#0e#)) OR
 					(reg_q369 AND symb_decoder(16#5c#)) OR
 					(reg_q369 AND symb_decoder(16#20#)) OR
 					(reg_q369 AND symb_decoder(16#24#)) OR
 					(reg_q369 AND symb_decoder(16#4d#)) OR
 					(reg_q369 AND symb_decoder(16#ea#)) OR
 					(reg_q369 AND symb_decoder(16#82#)) OR
 					(reg_q369 AND symb_decoder(16#e6#)) OR
 					(reg_q369 AND symb_decoder(16#db#)) OR
 					(reg_q369 AND symb_decoder(16#61#)) OR
 					(reg_q369 AND symb_decoder(16#e8#)) OR
 					(reg_q369 AND symb_decoder(16#dd#)) OR
 					(reg_q369 AND symb_decoder(16#a7#)) OR
 					(reg_q369 AND symb_decoder(16#50#)) OR
 					(reg_q369 AND symb_decoder(16#66#)) OR
 					(reg_q369 AND symb_decoder(16#41#)) OR
 					(reg_q369 AND symb_decoder(16#9a#)) OR
 					(reg_q369 AND symb_decoder(16#c3#)) OR
 					(reg_q369 AND symb_decoder(16#6c#)) OR
 					(reg_q369 AND symb_decoder(16#cd#)) OR
 					(reg_q369 AND symb_decoder(16#d8#)) OR
 					(reg_q369 AND symb_decoder(16#88#)) OR
 					(reg_q369 AND symb_decoder(16#5e#)) OR
 					(reg_q369 AND symb_decoder(16#3b#)) OR
 					(reg_q369 AND symb_decoder(16#f0#)) OR
 					(reg_q369 AND symb_decoder(16#2f#)) OR
 					(reg_q369 AND symb_decoder(16#b2#)) OR
 					(reg_q369 AND symb_decoder(16#b5#)) OR
 					(reg_q369 AND symb_decoder(16#a4#)) OR
 					(reg_q369 AND symb_decoder(16#23#)) OR
 					(reg_q369 AND symb_decoder(16#03#)) OR
 					(reg_q369 AND symb_decoder(16#29#)) OR
 					(reg_q369 AND symb_decoder(16#1b#)) OR
 					(reg_q369 AND symb_decoder(16#17#)) OR
 					(reg_q369 AND symb_decoder(16#ee#)) OR
 					(reg_q369 AND symb_decoder(16#08#)) OR
 					(reg_q369 AND symb_decoder(16#34#)) OR
 					(reg_q369 AND symb_decoder(16#af#)) OR
 					(reg_q369 AND symb_decoder(16#59#)) OR
 					(reg_q369 AND symb_decoder(16#e4#)) OR
 					(reg_q369 AND symb_decoder(16#49#)) OR
 					(reg_q369 AND symb_decoder(16#73#)) OR
 					(reg_q369 AND symb_decoder(16#bd#)) OR
 					(reg_q369 AND symb_decoder(16#0f#)) OR
 					(reg_q369 AND symb_decoder(16#6b#)) OR
 					(reg_q369 AND symb_decoder(16#63#)) OR
 					(reg_q369 AND symb_decoder(16#c0#)) OR
 					(reg_q369 AND symb_decoder(16#15#)) OR
 					(reg_q369 AND symb_decoder(16#18#)) OR
 					(reg_q369 AND symb_decoder(16#02#)) OR
 					(reg_q369 AND symb_decoder(16#f4#)) OR
 					(reg_q369 AND symb_decoder(16#a9#)) OR
 					(reg_q369 AND symb_decoder(16#12#)) OR
 					(reg_q369 AND symb_decoder(16#d1#)) OR
 					(reg_q369 AND symb_decoder(16#7f#)) OR
 					(reg_q369 AND symb_decoder(16#7d#)) OR
 					(reg_q369 AND symb_decoder(16#dc#)) OR
 					(reg_q369 AND symb_decoder(16#87#)) OR
 					(reg_q369 AND symb_decoder(16#ad#)) OR
 					(reg_q369 AND symb_decoder(16#16#)) OR
 					(reg_q369 AND symb_decoder(16#55#)) OR
 					(reg_q369 AND symb_decoder(16#8c#)) OR
 					(reg_q369 AND symb_decoder(16#ab#)) OR
 					(reg_q369 AND symb_decoder(16#2b#)) OR
 					(reg_q369 AND symb_decoder(16#8d#)) OR
 					(reg_q369 AND symb_decoder(16#00#)) OR
 					(reg_q369 AND symb_decoder(16#a5#)) OR
 					(reg_q369 AND symb_decoder(16#0b#)) OR
 					(reg_q369 AND symb_decoder(16#e5#)) OR
 					(reg_q369 AND symb_decoder(16#bc#)) OR
 					(reg_q369 AND symb_decoder(16#37#)) OR
 					(reg_q369 AND symb_decoder(16#76#)) OR
 					(reg_q369 AND symb_decoder(16#ef#)) OR
 					(reg_q369 AND symb_decoder(16#c2#)) OR
 					(reg_q369 AND symb_decoder(16#f9#)) OR
 					(reg_q369 AND symb_decoder(16#74#)) OR
 					(reg_q369 AND symb_decoder(16#53#)) OR
 					(reg_q369 AND symb_decoder(16#7e#)) OR
 					(reg_q369 AND symb_decoder(16#b6#)) OR
 					(reg_q369 AND symb_decoder(16#5f#)) OR
 					(reg_q369 AND symb_decoder(16#eb#)) OR
 					(reg_q369 AND symb_decoder(16#86#)) OR
 					(reg_q369 AND symb_decoder(16#42#)) OR
 					(reg_q369 AND symb_decoder(16#13#)) OR
 					(reg_q369 AND symb_decoder(16#71#)) OR
 					(reg_q369 AND symb_decoder(16#1f#)) OR
 					(reg_q369 AND symb_decoder(16#a1#)) OR
 					(reg_q369 AND symb_decoder(16#4f#)) OR
 					(reg_q369 AND symb_decoder(16#0c#)) OR
 					(reg_q369 AND symb_decoder(16#85#)) OR
 					(reg_q369 AND symb_decoder(16#38#)) OR
 					(reg_q369 AND symb_decoder(16#56#)) OR
 					(reg_q369 AND symb_decoder(16#92#)) OR
 					(reg_q369 AND symb_decoder(16#4a#)) OR
 					(reg_q369 AND symb_decoder(16#52#)) OR
 					(reg_q369 AND symb_decoder(16#28#)) OR
 					(reg_q369 AND symb_decoder(16#c8#)) OR
 					(reg_q369 AND symb_decoder(16#35#)) OR
 					(reg_q369 AND symb_decoder(16#04#)) OR
 					(reg_q369 AND symb_decoder(16#83#)) OR
 					(reg_q369 AND symb_decoder(16#4c#)) OR
 					(reg_q369 AND symb_decoder(16#26#)) OR
 					(reg_q369 AND symb_decoder(16#f3#)) OR
 					(reg_q369 AND symb_decoder(16#9b#)) OR
 					(reg_q369 AND symb_decoder(16#84#)) OR
 					(reg_q369 AND symb_decoder(16#22#)) OR
 					(reg_q369 AND symb_decoder(16#21#)) OR
 					(reg_q369 AND symb_decoder(16#3f#)) OR
 					(reg_q369 AND symb_decoder(16#ba#)) OR
 					(reg_q369 AND symb_decoder(16#43#)) OR
 					(reg_q369 AND symb_decoder(16#07#)) OR
 					(reg_q369 AND symb_decoder(16#a2#)) OR
 					(reg_q369 AND symb_decoder(16#95#)) OR
 					(reg_q369 AND symb_decoder(16#b8#)) OR
 					(reg_q369 AND symb_decoder(16#d3#)) OR
 					(reg_q369 AND symb_decoder(16#d5#)) OR
 					(reg_q369 AND symb_decoder(16#bb#)) OR
 					(reg_q369 AND symb_decoder(16#f6#)) OR
 					(reg_q369 AND symb_decoder(16#f1#)) OR
 					(reg_q369 AND symb_decoder(16#5d#)) OR
 					(reg_q369 AND symb_decoder(16#79#)) OR
 					(reg_q369 AND symb_decoder(16#81#)) OR
 					(reg_q369 AND symb_decoder(16#01#)) OR
 					(reg_q369 AND symb_decoder(16#c5#)) OR
 					(reg_q369 AND symb_decoder(16#fa#)) OR
 					(reg_q369 AND symb_decoder(16#36#)) OR
 					(reg_q369 AND symb_decoder(16#9c#)) OR
 					(reg_q369 AND symb_decoder(16#98#)) OR
 					(reg_q369 AND symb_decoder(16#70#)) OR
 					(reg_q369 AND symb_decoder(16#89#)) OR
 					(reg_q369 AND symb_decoder(16#9e#)) OR
 					(reg_q369 AND symb_decoder(16#80#)) OR
 					(reg_q369 AND symb_decoder(16#c4#)) OR
 					(reg_q369 AND symb_decoder(16#67#)) OR
 					(reg_q369 AND symb_decoder(16#7b#)) OR
 					(reg_q369 AND symb_decoder(16#65#)) OR
 					(reg_q369 AND symb_decoder(16#c9#)) OR
 					(reg_q369 AND symb_decoder(16#cc#)) OR
 					(reg_q369 AND symb_decoder(16#4b#)) OR
 					(reg_q369 AND symb_decoder(16#9d#)) OR
 					(reg_q369 AND symb_decoder(16#ae#)) OR
 					(reg_q369 AND symb_decoder(16#c6#)) OR
 					(reg_q369 AND symb_decoder(16#3d#)) OR
 					(reg_q369 AND symb_decoder(16#90#)) OR
 					(reg_q369 AND symb_decoder(16#54#)) OR
 					(reg_q369 AND symb_decoder(16#cb#)) OR
 					(reg_q369 AND symb_decoder(16#7c#)) OR
 					(reg_q369 AND symb_decoder(16#2e#)) OR
 					(reg_q369 AND symb_decoder(16#2c#)) OR
 					(reg_q369 AND symb_decoder(16#a6#)) OR
 					(reg_q369 AND symb_decoder(16#ff#)) OR
 					(reg_q369 AND symb_decoder(16#46#)) OR
 					(reg_q369 AND symb_decoder(16#fb#)) OR
 					(reg_q369 AND symb_decoder(16#a0#)) OR
 					(reg_q369 AND symb_decoder(16#8e#)) OR
 					(reg_q369 AND symb_decoder(16#68#)) OR
 					(reg_q369 AND symb_decoder(16#44#)) OR
 					(reg_q369 AND symb_decoder(16#7a#)) OR
 					(reg_q369 AND symb_decoder(16#e1#)) OR
 					(reg_q369 AND symb_decoder(16#ac#)) OR
 					(reg_q369 AND symb_decoder(16#1a#)) OR
 					(reg_q369 AND symb_decoder(16#e7#)) OR
 					(reg_q369 AND symb_decoder(16#48#)) OR
 					(reg_q369 AND symb_decoder(16#8b#)) OR
 					(reg_q369 AND symb_decoder(16#be#)) OR
 					(reg_q369 AND symb_decoder(16#b1#)) OR
 					(reg_q369 AND symb_decoder(16#45#)) OR
 					(reg_q369 AND symb_decoder(16#f5#)) OR
 					(reg_q369 AND symb_decoder(16#93#)) OR
 					(reg_q369 AND symb_decoder(16#e9#)) OR
 					(reg_q369 AND symb_decoder(16#8a#)) OR
 					(reg_q369 AND symb_decoder(16#72#)) OR
 					(reg_q369 AND symb_decoder(16#aa#)) OR
 					(reg_q369 AND symb_decoder(16#b7#)) OR
 					(reg_q369 AND symb_decoder(16#5a#)) OR
 					(reg_q369 AND symb_decoder(16#58#)) OR
 					(reg_q369 AND symb_decoder(16#60#)) OR
 					(reg_q369 AND symb_decoder(16#fc#)) OR
 					(reg_q369 AND symb_decoder(16#d2#)) OR
 					(reg_q369 AND symb_decoder(16#f2#)) OR
 					(reg_q369 AND symb_decoder(16#14#)) OR
 					(reg_q369 AND symb_decoder(16#6a#)) OR
 					(reg_q369 AND symb_decoder(16#b3#)) OR
 					(reg_q369 AND symb_decoder(16#ec#)) OR
 					(reg_q369 AND symb_decoder(16#05#)) OR
 					(reg_q369 AND symb_decoder(16#1d#)) OR
 					(reg_q369 AND symb_decoder(16#ed#)) OR
 					(reg_q369 AND symb_decoder(16#bf#)) OR
 					(reg_q369 AND symb_decoder(16#fd#)) OR
 					(reg_q369 AND symb_decoder(16#f8#)) OR
 					(reg_q369 AND symb_decoder(16#e2#)) OR
 					(reg_q369 AND symb_decoder(16#25#)) OR
 					(reg_q369 AND symb_decoder(16#51#)) OR
 					(reg_q369 AND symb_decoder(16#64#)) OR
 					(reg_q369 AND symb_decoder(16#3a#)) OR
 					(reg_q369 AND symb_decoder(16#94#)) OR
 					(reg_q369 AND symb_decoder(16#b0#)) OR
 					(reg_q369 AND symb_decoder(16#09#)) OR
 					(reg_q369 AND symb_decoder(16#cf#)) OR
 					(reg_q369 AND symb_decoder(16#da#)) OR
 					(reg_q369 AND symb_decoder(16#32#)) OR
 					(reg_q369 AND symb_decoder(16#de#)) OR
 					(reg_q369 AND symb_decoder(16#d9#)) OR
 					(reg_q369 AND symb_decoder(16#6f#)) OR
 					(reg_q369 AND symb_decoder(16#d0#)) OR
 					(reg_q369 AND symb_decoder(16#d4#)) OR
 					(reg_q369 AND symb_decoder(16#6e#)) OR
 					(reg_q369 AND symb_decoder(16#b9#)) OR
 					(reg_q369 AND symb_decoder(16#fe#)) OR
 					(reg_q369 AND symb_decoder(16#2a#)) OR
 					(reg_q369 AND symb_decoder(16#d6#)) OR
 					(reg_q369 AND symb_decoder(16#ce#)) OR
 					(reg_q369 AND symb_decoder(16#6d#)) OR
 					(reg_q369 AND symb_decoder(16#ca#)) OR
 					(reg_q369 AND symb_decoder(16#40#)) OR
 					(reg_q369 AND symb_decoder(16#2d#)) OR
 					(reg_q369 AND symb_decoder(16#30#)) OR
 					(reg_q369 AND symb_decoder(16#99#)) OR
 					(reg_q369 AND symb_decoder(16#f7#));
reg_q526_in <= (reg_q522 AND symb_decoder(16#2f#)) OR
 					(reg_q542 AND symb_decoder(16#2f#));
reg_q800_in <= (reg_q788 AND symb_decoder(16#bf#)) OR
 					(reg_q788 AND symb_decoder(16#be#)) OR
 					(reg_q788 AND symb_decoder(16#5f#)) OR
 					(reg_q788 AND symb_decoder(16#db#)) OR
 					(reg_q788 AND symb_decoder(16#26#)) OR
 					(reg_q788 AND symb_decoder(16#76#)) OR
 					(reg_q788 AND symb_decoder(16#01#)) OR
 					(reg_q788 AND symb_decoder(16#8b#)) OR
 					(reg_q788 AND symb_decoder(16#21#)) OR
 					(reg_q788 AND symb_decoder(16#2a#)) OR
 					(reg_q788 AND symb_decoder(16#c5#)) OR
 					(reg_q788 AND symb_decoder(16#58#)) OR
 					(reg_q788 AND symb_decoder(16#59#)) OR
 					(reg_q788 AND symb_decoder(16#a8#)) OR
 					(reg_q788 AND symb_decoder(16#70#)) OR
 					(reg_q788 AND symb_decoder(16#9d#)) OR
 					(reg_q788 AND symb_decoder(16#60#)) OR
 					(reg_q788 AND symb_decoder(16#2c#)) OR
 					(reg_q788 AND symb_decoder(16#51#)) OR
 					(reg_q788 AND symb_decoder(16#62#)) OR
 					(reg_q788 AND symb_decoder(16#eb#)) OR
 					(reg_q788 AND symb_decoder(16#84#)) OR
 					(reg_q788 AND symb_decoder(16#0e#)) OR
 					(reg_q788 AND symb_decoder(16#32#)) OR
 					(reg_q788 AND symb_decoder(16#9a#)) OR
 					(reg_q788 AND symb_decoder(16#1d#)) OR
 					(reg_q788 AND symb_decoder(16#1c#)) OR
 					(reg_q788 AND symb_decoder(16#6d#)) OR
 					(reg_q788 AND symb_decoder(16#e8#)) OR
 					(reg_q788 AND symb_decoder(16#0b#)) OR
 					(reg_q788 AND symb_decoder(16#40#)) OR
 					(reg_q788 AND symb_decoder(16#5d#)) OR
 					(reg_q788 AND symb_decoder(16#fd#)) OR
 					(reg_q788 AND symb_decoder(16#39#)) OR
 					(reg_q788 AND symb_decoder(16#13#)) OR
 					(reg_q788 AND symb_decoder(16#03#)) OR
 					(reg_q788 AND symb_decoder(16#ff#)) OR
 					(reg_q788 AND symb_decoder(16#2e#)) OR
 					(reg_q788 AND symb_decoder(16#48#)) OR
 					(reg_q788 AND symb_decoder(16#fc#)) OR
 					(reg_q788 AND symb_decoder(16#e2#)) OR
 					(reg_q788 AND symb_decoder(16#b9#)) OR
 					(reg_q788 AND symb_decoder(16#6f#)) OR
 					(reg_q788 AND symb_decoder(16#74#)) OR
 					(reg_q788 AND symb_decoder(16#02#)) OR
 					(reg_q788 AND symb_decoder(16#97#)) OR
 					(reg_q788 AND symb_decoder(16#e4#)) OR
 					(reg_q788 AND symb_decoder(16#8a#)) OR
 					(reg_q788 AND symb_decoder(16#aa#)) OR
 					(reg_q788 AND symb_decoder(16#07#)) OR
 					(reg_q788 AND symb_decoder(16#f7#)) OR
 					(reg_q788 AND symb_decoder(16#25#)) OR
 					(reg_q788 AND symb_decoder(16#b4#)) OR
 					(reg_q788 AND symb_decoder(16#29#)) OR
 					(reg_q788 AND symb_decoder(16#f3#)) OR
 					(reg_q788 AND symb_decoder(16#52#)) OR
 					(reg_q788 AND symb_decoder(16#4e#)) OR
 					(reg_q788 AND symb_decoder(16#5e#)) OR
 					(reg_q788 AND symb_decoder(16#b2#)) OR
 					(reg_q788 AND symb_decoder(16#90#)) OR
 					(reg_q788 AND symb_decoder(16#b0#)) OR
 					(reg_q788 AND symb_decoder(16#cf#)) OR
 					(reg_q788 AND symb_decoder(16#69#)) OR
 					(reg_q788 AND symb_decoder(16#e0#)) OR
 					(reg_q788 AND symb_decoder(16#53#)) OR
 					(reg_q788 AND symb_decoder(16#82#)) OR
 					(reg_q788 AND symb_decoder(16#1b#)) OR
 					(reg_q788 AND symb_decoder(16#20#)) OR
 					(reg_q788 AND symb_decoder(16#dc#)) OR
 					(reg_q788 AND symb_decoder(16#24#)) OR
 					(reg_q788 AND symb_decoder(16#c7#)) OR
 					(reg_q788 AND symb_decoder(16#4d#)) OR
 					(reg_q788 AND symb_decoder(16#5a#)) OR
 					(reg_q788 AND symb_decoder(16#22#)) OR
 					(reg_q788 AND symb_decoder(16#a5#)) OR
 					(reg_q788 AND symb_decoder(16#67#)) OR
 					(reg_q788 AND symb_decoder(16#3c#)) OR
 					(reg_q788 AND symb_decoder(16#e9#)) OR
 					(reg_q788 AND symb_decoder(16#79#)) OR
 					(reg_q788 AND symb_decoder(16#78#)) OR
 					(reg_q788 AND symb_decoder(16#6c#)) OR
 					(reg_q788 AND symb_decoder(16#68#)) OR
 					(reg_q788 AND symb_decoder(16#86#)) OR
 					(reg_q788 AND symb_decoder(16#10#)) OR
 					(reg_q788 AND symb_decoder(16#31#)) OR
 					(reg_q788 AND symb_decoder(16#38#)) OR
 					(reg_q788 AND symb_decoder(16#23#)) OR
 					(reg_q788 AND symb_decoder(16#ad#)) OR
 					(reg_q788 AND symb_decoder(16#11#)) OR
 					(reg_q788 AND symb_decoder(16#80#)) OR
 					(reg_q788 AND symb_decoder(16#f8#)) OR
 					(reg_q788 AND symb_decoder(16#45#)) OR
 					(reg_q788 AND symb_decoder(16#15#)) OR
 					(reg_q788 AND symb_decoder(16#d2#)) OR
 					(reg_q788 AND symb_decoder(16#5b#)) OR
 					(reg_q788 AND symb_decoder(16#3b#)) OR
 					(reg_q788 AND symb_decoder(16#a1#)) OR
 					(reg_q788 AND symb_decoder(16#b8#)) OR
 					(reg_q788 AND symb_decoder(16#d4#)) OR
 					(reg_q788 AND symb_decoder(16#8e#)) OR
 					(reg_q788 AND symb_decoder(16#99#)) OR
 					(reg_q788 AND symb_decoder(16#c2#)) OR
 					(reg_q788 AND symb_decoder(16#7f#)) OR
 					(reg_q788 AND symb_decoder(16#cb#)) OR
 					(reg_q788 AND symb_decoder(16#63#)) OR
 					(reg_q788 AND symb_decoder(16#b5#)) OR
 					(reg_q788 AND symb_decoder(16#4b#)) OR
 					(reg_q788 AND symb_decoder(16#2d#)) OR
 					(reg_q788 AND symb_decoder(16#30#)) OR
 					(reg_q788 AND symb_decoder(16#61#)) OR
 					(reg_q788 AND symb_decoder(16#a0#)) OR
 					(reg_q788 AND symb_decoder(16#f6#)) OR
 					(reg_q788 AND symb_decoder(16#c3#)) OR
 					(reg_q788 AND symb_decoder(16#5c#)) OR
 					(reg_q788 AND symb_decoder(16#d5#)) OR
 					(reg_q788 AND symb_decoder(16#7b#)) OR
 					(reg_q788 AND symb_decoder(16#fe#)) OR
 					(reg_q788 AND symb_decoder(16#cd#)) OR
 					(reg_q788 AND symb_decoder(16#6e#)) OR
 					(reg_q788 AND symb_decoder(16#72#)) OR
 					(reg_q788 AND symb_decoder(16#e7#)) OR
 					(reg_q788 AND symb_decoder(16#c4#)) OR
 					(reg_q788 AND symb_decoder(16#2b#)) OR
 					(reg_q788 AND symb_decoder(16#f0#)) OR
 					(reg_q788 AND symb_decoder(16#14#)) OR
 					(reg_q788 AND symb_decoder(16#df#)) OR
 					(reg_q788 AND symb_decoder(16#3f#)) OR
 					(reg_q788 AND symb_decoder(16#00#)) OR
 					(reg_q788 AND symb_decoder(16#08#)) OR
 					(reg_q788 AND symb_decoder(16#d7#)) OR
 					(reg_q788 AND symb_decoder(16#c9#)) OR
 					(reg_q788 AND symb_decoder(16#a6#)) OR
 					(reg_q788 AND symb_decoder(16#64#)) OR
 					(reg_q788 AND symb_decoder(16#a7#)) OR
 					(reg_q788 AND symb_decoder(16#d3#)) OR
 					(reg_q788 AND symb_decoder(16#44#)) OR
 					(reg_q788 AND symb_decoder(16#8f#)) OR
 					(reg_q788 AND symb_decoder(16#c1#)) OR
 					(reg_q788 AND symb_decoder(16#d8#)) OR
 					(reg_q788 AND symb_decoder(16#54#)) OR
 					(reg_q788 AND symb_decoder(16#34#)) OR
 					(reg_q788 AND symb_decoder(16#e6#)) OR
 					(reg_q788 AND symb_decoder(16#bb#)) OR
 					(reg_q788 AND symb_decoder(16#b6#)) OR
 					(reg_q788 AND symb_decoder(16#65#)) OR
 					(reg_q788 AND symb_decoder(16#3d#)) OR
 					(reg_q788 AND symb_decoder(16#f5#)) OR
 					(reg_q788 AND symb_decoder(16#b7#)) OR
 					(reg_q788 AND symb_decoder(16#f1#)) OR
 					(reg_q788 AND symb_decoder(16#9f#)) OR
 					(reg_q788 AND symb_decoder(16#4c#)) OR
 					(reg_q788 AND symb_decoder(16#af#)) OR
 					(reg_q788 AND symb_decoder(16#cc#)) OR
 					(reg_q788 AND symb_decoder(16#92#)) OR
 					(reg_q788 AND symb_decoder(16#09#)) OR
 					(reg_q788 AND symb_decoder(16#9e#)) OR
 					(reg_q788 AND symb_decoder(16#e1#)) OR
 					(reg_q788 AND symb_decoder(16#ca#)) OR
 					(reg_q788 AND symb_decoder(16#ce#)) OR
 					(reg_q788 AND symb_decoder(16#3e#)) OR
 					(reg_q788 AND symb_decoder(16#e5#)) OR
 					(reg_q788 AND symb_decoder(16#19#)) OR
 					(reg_q788 AND symb_decoder(16#94#)) OR
 					(reg_q788 AND symb_decoder(16#83#)) OR
 					(reg_q788 AND symb_decoder(16#87#)) OR
 					(reg_q788 AND symb_decoder(16#56#)) OR
 					(reg_q788 AND symb_decoder(16#81#)) OR
 					(reg_q788 AND symb_decoder(16#1f#)) OR
 					(reg_q788 AND symb_decoder(16#6a#)) OR
 					(reg_q788 AND symb_decoder(16#06#)) OR
 					(reg_q788 AND symb_decoder(16#c6#)) OR
 					(reg_q788 AND symb_decoder(16#75#)) OR
 					(reg_q788 AND symb_decoder(16#9c#)) OR
 					(reg_q788 AND symb_decoder(16#ba#)) OR
 					(reg_q788 AND symb_decoder(16#12#)) OR
 					(reg_q788 AND symb_decoder(16#dd#)) OR
 					(reg_q788 AND symb_decoder(16#8d#)) OR
 					(reg_q788 AND symb_decoder(16#73#)) OR
 					(reg_q788 AND symb_decoder(16#2f#)) OR
 					(reg_q788 AND symb_decoder(16#0f#)) OR
 					(reg_q788 AND symb_decoder(16#1e#)) OR
 					(reg_q788 AND symb_decoder(16#77#)) OR
 					(reg_q788 AND symb_decoder(16#91#)) OR
 					(reg_q788 AND symb_decoder(16#93#)) OR
 					(reg_q788 AND symb_decoder(16#1a#)) OR
 					(reg_q788 AND symb_decoder(16#ef#)) OR
 					(reg_q788 AND symb_decoder(16#37#)) OR
 					(reg_q788 AND symb_decoder(16#8c#)) OR
 					(reg_q788 AND symb_decoder(16#a9#)) OR
 					(reg_q788 AND symb_decoder(16#d6#)) OR
 					(reg_q788 AND symb_decoder(16#ea#)) OR
 					(reg_q788 AND symb_decoder(16#16#)) OR
 					(reg_q788 AND symb_decoder(16#98#)) OR
 					(reg_q788 AND symb_decoder(16#46#)) OR
 					(reg_q788 AND symb_decoder(16#43#)) OR
 					(reg_q788 AND symb_decoder(16#ae#)) OR
 					(reg_q788 AND symb_decoder(16#28#)) OR
 					(reg_q788 AND symb_decoder(16#ec#)) OR
 					(reg_q788 AND symb_decoder(16#95#)) OR
 					(reg_q788 AND symb_decoder(16#3a#)) OR
 					(reg_q788 AND symb_decoder(16#88#)) OR
 					(reg_q788 AND symb_decoder(16#c8#)) OR
 					(reg_q788 AND symb_decoder(16#04#)) OR
 					(reg_q788 AND symb_decoder(16#a4#)) OR
 					(reg_q788 AND symb_decoder(16#66#)) OR
 					(reg_q788 AND symb_decoder(16#de#)) OR
 					(reg_q788 AND symb_decoder(16#b1#)) OR
 					(reg_q788 AND symb_decoder(16#42#)) OR
 					(reg_q788 AND symb_decoder(16#f2#)) OR
 					(reg_q788 AND symb_decoder(16#e3#)) OR
 					(reg_q788 AND symb_decoder(16#7a#)) OR
 					(reg_q788 AND symb_decoder(16#d9#)) OR
 					(reg_q788 AND symb_decoder(16#c0#)) OR
 					(reg_q788 AND symb_decoder(16#33#)) OR
 					(reg_q788 AND symb_decoder(16#a2#)) OR
 					(reg_q788 AND symb_decoder(16#ac#)) OR
 					(reg_q788 AND symb_decoder(16#36#)) OR
 					(reg_q788 AND symb_decoder(16#27#)) OR
 					(reg_q788 AND symb_decoder(16#d1#)) OR
 					(reg_q788 AND symb_decoder(16#55#)) OR
 					(reg_q788 AND symb_decoder(16#9b#)) OR
 					(reg_q788 AND symb_decoder(16#35#)) OR
 					(reg_q788 AND symb_decoder(16#49#)) OR
 					(reg_q788 AND symb_decoder(16#bd#)) OR
 					(reg_q788 AND symb_decoder(16#a3#)) OR
 					(reg_q788 AND symb_decoder(16#f4#)) OR
 					(reg_q788 AND symb_decoder(16#ee#)) OR
 					(reg_q788 AND symb_decoder(16#85#)) OR
 					(reg_q788 AND symb_decoder(16#0c#)) OR
 					(reg_q788 AND symb_decoder(16#71#)) OR
 					(reg_q788 AND symb_decoder(16#57#)) OR
 					(reg_q788 AND symb_decoder(16#bc#)) OR
 					(reg_q788 AND symb_decoder(16#96#)) OR
 					(reg_q788 AND symb_decoder(16#7e#)) OR
 					(reg_q788 AND symb_decoder(16#6b#)) OR
 					(reg_q788 AND symb_decoder(16#ab#)) OR
 					(reg_q788 AND symb_decoder(16#18#)) OR
 					(reg_q788 AND symb_decoder(16#50#)) OR
 					(reg_q788 AND symb_decoder(16#ed#)) OR
 					(reg_q788 AND symb_decoder(16#47#)) OR
 					(reg_q788 AND symb_decoder(16#d0#)) OR
 					(reg_q788 AND symb_decoder(16#b3#)) OR
 					(reg_q788 AND symb_decoder(16#f9#)) OR
 					(reg_q788 AND symb_decoder(16#fa#)) OR
 					(reg_q788 AND symb_decoder(16#4f#)) OR
 					(reg_q788 AND symb_decoder(16#da#)) OR
 					(reg_q788 AND symb_decoder(16#05#)) OR
 					(reg_q788 AND symb_decoder(16#7c#)) OR
 					(reg_q788 AND symb_decoder(16#89#)) OR
 					(reg_q788 AND symb_decoder(16#fb#)) OR
 					(reg_q788 AND symb_decoder(16#17#)) OR
 					(reg_q788 AND symb_decoder(16#4a#)) OR
 					(reg_q788 AND symb_decoder(16#41#)) OR
 					(reg_q788 AND symb_decoder(16#7d#)) OR
 					(reg_q800 AND symb_decoder(16#04#)) OR
 					(reg_q800 AND symb_decoder(16#bd#)) OR
 					(reg_q800 AND symb_decoder(16#f5#)) OR
 					(reg_q800 AND symb_decoder(16#90#)) OR
 					(reg_q800 AND symb_decoder(16#41#)) OR
 					(reg_q800 AND symb_decoder(16#b1#)) OR
 					(reg_q800 AND symb_decoder(16#b2#)) OR
 					(reg_q800 AND symb_decoder(16#8a#)) OR
 					(reg_q800 AND symb_decoder(16#d4#)) OR
 					(reg_q800 AND symb_decoder(16#de#)) OR
 					(reg_q800 AND symb_decoder(16#f7#)) OR
 					(reg_q800 AND symb_decoder(16#5d#)) OR
 					(reg_q800 AND symb_decoder(16#cd#)) OR
 					(reg_q800 AND symb_decoder(16#c9#)) OR
 					(reg_q800 AND symb_decoder(16#92#)) OR
 					(reg_q800 AND symb_decoder(16#4b#)) OR
 					(reg_q800 AND symb_decoder(16#35#)) OR
 					(reg_q800 AND symb_decoder(16#91#)) OR
 					(reg_q800 AND symb_decoder(16#eb#)) OR
 					(reg_q800 AND symb_decoder(16#ad#)) OR
 					(reg_q800 AND symb_decoder(16#a8#)) OR
 					(reg_q800 AND symb_decoder(16#54#)) OR
 					(reg_q800 AND symb_decoder(16#57#)) OR
 					(reg_q800 AND symb_decoder(16#79#)) OR
 					(reg_q800 AND symb_decoder(16#09#)) OR
 					(reg_q800 AND symb_decoder(16#6d#)) OR
 					(reg_q800 AND symb_decoder(16#e6#)) OR
 					(reg_q800 AND symb_decoder(16#7c#)) OR
 					(reg_q800 AND symb_decoder(16#d5#)) OR
 					(reg_q800 AND symb_decoder(16#bb#)) OR
 					(reg_q800 AND symb_decoder(16#a5#)) OR
 					(reg_q800 AND symb_decoder(16#e2#)) OR
 					(reg_q800 AND symb_decoder(16#6e#)) OR
 					(reg_q800 AND symb_decoder(16#d8#)) OR
 					(reg_q800 AND symb_decoder(16#11#)) OR
 					(reg_q800 AND symb_decoder(16#4a#)) OR
 					(reg_q800 AND symb_decoder(16#26#)) OR
 					(reg_q800 AND symb_decoder(16#0f#)) OR
 					(reg_q800 AND symb_decoder(16#77#)) OR
 					(reg_q800 AND symb_decoder(16#14#)) OR
 					(reg_q800 AND symb_decoder(16#6f#)) OR
 					(reg_q800 AND symb_decoder(16#05#)) OR
 					(reg_q800 AND symb_decoder(16#c8#)) OR
 					(reg_q800 AND symb_decoder(16#16#)) OR
 					(reg_q800 AND symb_decoder(16#4f#)) OR
 					(reg_q800 AND symb_decoder(16#17#)) OR
 					(reg_q800 AND symb_decoder(16#95#)) OR
 					(reg_q800 AND symb_decoder(16#fc#)) OR
 					(reg_q800 AND symb_decoder(16#4e#)) OR
 					(reg_q800 AND symb_decoder(16#7a#)) OR
 					(reg_q800 AND symb_decoder(16#d6#)) OR
 					(reg_q800 AND symb_decoder(16#66#)) OR
 					(reg_q800 AND symb_decoder(16#4c#)) OR
 					(reg_q800 AND symb_decoder(16#d0#)) OR
 					(reg_q800 AND symb_decoder(16#33#)) OR
 					(reg_q800 AND symb_decoder(16#fe#)) OR
 					(reg_q800 AND symb_decoder(16#d2#)) OR
 					(reg_q800 AND symb_decoder(16#bf#)) OR
 					(reg_q800 AND symb_decoder(16#96#)) OR
 					(reg_q800 AND symb_decoder(16#fd#)) OR
 					(reg_q800 AND symb_decoder(16#86#)) OR
 					(reg_q800 AND symb_decoder(16#98#)) OR
 					(reg_q800 AND symb_decoder(16#9f#)) OR
 					(reg_q800 AND symb_decoder(16#6b#)) OR
 					(reg_q800 AND symb_decoder(16#df#)) OR
 					(reg_q800 AND symb_decoder(16#da#)) OR
 					(reg_q800 AND symb_decoder(16#d3#)) OR
 					(reg_q800 AND symb_decoder(16#08#)) OR
 					(reg_q800 AND symb_decoder(16#23#)) OR
 					(reg_q800 AND symb_decoder(16#5e#)) OR
 					(reg_q800 AND symb_decoder(16#07#)) OR
 					(reg_q800 AND symb_decoder(16#9d#)) OR
 					(reg_q800 AND symb_decoder(16#ce#)) OR
 					(reg_q800 AND symb_decoder(16#81#)) OR
 					(reg_q800 AND symb_decoder(16#ec#)) OR
 					(reg_q800 AND symb_decoder(16#12#)) OR
 					(reg_q800 AND symb_decoder(16#d9#)) OR
 					(reg_q800 AND symb_decoder(16#27#)) OR
 					(reg_q800 AND symb_decoder(16#75#)) OR
 					(reg_q800 AND symb_decoder(16#03#)) OR
 					(reg_q800 AND symb_decoder(16#ab#)) OR
 					(reg_q800 AND symb_decoder(16#c5#)) OR
 					(reg_q800 AND symb_decoder(16#f0#)) OR
 					(reg_q800 AND symb_decoder(16#13#)) OR
 					(reg_q800 AND symb_decoder(16#69#)) OR
 					(reg_q800 AND symb_decoder(16#e5#)) OR
 					(reg_q800 AND symb_decoder(16#55#)) OR
 					(reg_q800 AND symb_decoder(16#30#)) OR
 					(reg_q800 AND symb_decoder(16#b4#)) OR
 					(reg_q800 AND symb_decoder(16#ed#)) OR
 					(reg_q800 AND symb_decoder(16#1a#)) OR
 					(reg_q800 AND symb_decoder(16#53#)) OR
 					(reg_q800 AND symb_decoder(16#25#)) OR
 					(reg_q800 AND symb_decoder(16#15#)) OR
 					(reg_q800 AND symb_decoder(16#b6#)) OR
 					(reg_q800 AND symb_decoder(16#2a#)) OR
 					(reg_q800 AND symb_decoder(16#9a#)) OR
 					(reg_q800 AND symb_decoder(16#e1#)) OR
 					(reg_q800 AND symb_decoder(16#34#)) OR
 					(reg_q800 AND symb_decoder(16#a2#)) OR
 					(reg_q800 AND symb_decoder(16#1b#)) OR
 					(reg_q800 AND symb_decoder(16#63#)) OR
 					(reg_q800 AND symb_decoder(16#29#)) OR
 					(reg_q800 AND symb_decoder(16#af#)) OR
 					(reg_q800 AND symb_decoder(16#1c#)) OR
 					(reg_q800 AND symb_decoder(16#94#)) OR
 					(reg_q800 AND symb_decoder(16#42#)) OR
 					(reg_q800 AND symb_decoder(16#36#)) OR
 					(reg_q800 AND symb_decoder(16#b7#)) OR
 					(reg_q800 AND symb_decoder(16#3d#)) OR
 					(reg_q800 AND symb_decoder(16#32#)) OR
 					(reg_q800 AND symb_decoder(16#78#)) OR
 					(reg_q800 AND symb_decoder(16#e3#)) OR
 					(reg_q800 AND symb_decoder(16#3a#)) OR
 					(reg_q800 AND symb_decoder(16#c7#)) OR
 					(reg_q800 AND symb_decoder(16#d1#)) OR
 					(reg_q800 AND symb_decoder(16#1d#)) OR
 					(reg_q800 AND symb_decoder(16#28#)) OR
 					(reg_q800 AND symb_decoder(16#83#)) OR
 					(reg_q800 AND symb_decoder(16#00#)) OR
 					(reg_q800 AND symb_decoder(16#71#)) OR
 					(reg_q800 AND symb_decoder(16#49#)) OR
 					(reg_q800 AND symb_decoder(16#ff#)) OR
 					(reg_q800 AND symb_decoder(16#a9#)) OR
 					(reg_q800 AND symb_decoder(16#a4#)) OR
 					(reg_q800 AND symb_decoder(16#2e#)) OR
 					(reg_q800 AND symb_decoder(16#87#)) OR
 					(reg_q800 AND symb_decoder(16#1f#)) OR
 					(reg_q800 AND symb_decoder(16#68#)) OR
 					(reg_q800 AND symb_decoder(16#a7#)) OR
 					(reg_q800 AND symb_decoder(16#8b#)) OR
 					(reg_q800 AND symb_decoder(16#f1#)) OR
 					(reg_q800 AND symb_decoder(16#bc#)) OR
 					(reg_q800 AND symb_decoder(16#b0#)) OR
 					(reg_q800 AND symb_decoder(16#6a#)) OR
 					(reg_q800 AND symb_decoder(16#be#)) OR
 					(reg_q800 AND symb_decoder(16#24#)) OR
 					(reg_q800 AND symb_decoder(16#70#)) OR
 					(reg_q800 AND symb_decoder(16#7d#)) OR
 					(reg_q800 AND symb_decoder(16#48#)) OR
 					(reg_q800 AND symb_decoder(16#aa#)) OR
 					(reg_q800 AND symb_decoder(16#85#)) OR
 					(reg_q800 AND symb_decoder(16#47#)) OR
 					(reg_q800 AND symb_decoder(16#02#)) OR
 					(reg_q800 AND symb_decoder(16#c1#)) OR
 					(reg_q800 AND symb_decoder(16#1e#)) OR
 					(reg_q800 AND symb_decoder(16#06#)) OR
 					(reg_q800 AND symb_decoder(16#e0#)) OR
 					(reg_q800 AND symb_decoder(16#99#)) OR
 					(reg_q800 AND symb_decoder(16#45#)) OR
 					(reg_q800 AND symb_decoder(16#0c#)) OR
 					(reg_q800 AND symb_decoder(16#e4#)) OR
 					(reg_q800 AND symb_decoder(16#c0#)) OR
 					(reg_q800 AND symb_decoder(16#b9#)) OR
 					(reg_q800 AND symb_decoder(16#5c#)) OR
 					(reg_q800 AND symb_decoder(16#67#)) OR
 					(reg_q800 AND symb_decoder(16#f3#)) OR
 					(reg_q800 AND symb_decoder(16#6c#)) OR
 					(reg_q800 AND symb_decoder(16#5f#)) OR
 					(reg_q800 AND symb_decoder(16#97#)) OR
 					(reg_q800 AND symb_decoder(16#8e#)) OR
 					(reg_q800 AND symb_decoder(16#46#)) OR
 					(reg_q800 AND symb_decoder(16#52#)) OR
 					(reg_q800 AND symb_decoder(16#93#)) OR
 					(reg_q800 AND symb_decoder(16#a0#)) OR
 					(reg_q800 AND symb_decoder(16#f2#)) OR
 					(reg_q800 AND symb_decoder(16#dd#)) OR
 					(reg_q800 AND symb_decoder(16#f4#)) OR
 					(reg_q800 AND symb_decoder(16#7b#)) OR
 					(reg_q800 AND symb_decoder(16#84#)) OR
 					(reg_q800 AND symb_decoder(16#20#)) OR
 					(reg_q800 AND symb_decoder(16#a1#)) OR
 					(reg_q800 AND symb_decoder(16#21#)) OR
 					(reg_q800 AND symb_decoder(16#b8#)) OR
 					(reg_q800 AND symb_decoder(16#fb#)) OR
 					(reg_q800 AND symb_decoder(16#72#)) OR
 					(reg_q800 AND symb_decoder(16#d7#)) OR
 					(reg_q800 AND symb_decoder(16#e7#)) OR
 					(reg_q800 AND symb_decoder(16#db#)) OR
 					(reg_q800 AND symb_decoder(16#3f#)) OR
 					(reg_q800 AND symb_decoder(16#19#)) OR
 					(reg_q800 AND symb_decoder(16#7e#)) OR
 					(reg_q800 AND symb_decoder(16#5a#)) OR
 					(reg_q800 AND symb_decoder(16#9c#)) OR
 					(reg_q800 AND symb_decoder(16#39#)) OR
 					(reg_q800 AND symb_decoder(16#9e#)) OR
 					(reg_q800 AND symb_decoder(16#62#)) OR
 					(reg_q800 AND symb_decoder(16#31#)) OR
 					(reg_q800 AND symb_decoder(16#80#)) OR
 					(reg_q800 AND symb_decoder(16#a3#)) OR
 					(reg_q800 AND symb_decoder(16#ac#)) OR
 					(reg_q800 AND symb_decoder(16#43#)) OR
 					(reg_q800 AND symb_decoder(16#f6#)) OR
 					(reg_q800 AND symb_decoder(16#89#)) OR
 					(reg_q800 AND symb_decoder(16#5b#)) OR
 					(reg_q800 AND symb_decoder(16#ba#)) OR
 					(reg_q800 AND symb_decoder(16#64#)) OR
 					(reg_q800 AND symb_decoder(16#74#)) OR
 					(reg_q800 AND symb_decoder(16#01#)) OR
 					(reg_q800 AND symb_decoder(16#3e#)) OR
 					(reg_q800 AND symb_decoder(16#cf#)) OR
 					(reg_q800 AND symb_decoder(16#f8#)) OR
 					(reg_q800 AND symb_decoder(16#65#)) OR
 					(reg_q800 AND symb_decoder(16#50#)) OR
 					(reg_q800 AND symb_decoder(16#c4#)) OR
 					(reg_q800 AND symb_decoder(16#3b#)) OR
 					(reg_q800 AND symb_decoder(16#ca#)) OR
 					(reg_q800 AND symb_decoder(16#cc#)) OR
 					(reg_q800 AND symb_decoder(16#b5#)) OR
 					(reg_q800 AND symb_decoder(16#2b#)) OR
 					(reg_q800 AND symb_decoder(16#82#)) OR
 					(reg_q800 AND symb_decoder(16#37#)) OR
 					(reg_q800 AND symb_decoder(16#fa#)) OR
 					(reg_q800 AND symb_decoder(16#c3#)) OR
 					(reg_q800 AND symb_decoder(16#60#)) OR
 					(reg_q800 AND symb_decoder(16#4d#)) OR
 					(reg_q800 AND symb_decoder(16#88#)) OR
 					(reg_q800 AND symb_decoder(16#ea#)) OR
 					(reg_q800 AND symb_decoder(16#51#)) OR
 					(reg_q800 AND symb_decoder(16#dc#)) OR
 					(reg_q800 AND symb_decoder(16#f9#)) OR
 					(reg_q800 AND symb_decoder(16#10#)) OR
 					(reg_q800 AND symb_decoder(16#76#)) OR
 					(reg_q800 AND symb_decoder(16#61#)) OR
 					(reg_q800 AND symb_decoder(16#cb#)) OR
 					(reg_q800 AND symb_decoder(16#ae#)) OR
 					(reg_q800 AND symb_decoder(16#ee#)) OR
 					(reg_q800 AND symb_decoder(16#2c#)) OR
 					(reg_q800 AND symb_decoder(16#2d#)) OR
 					(reg_q800 AND symb_decoder(16#0e#)) OR
 					(reg_q800 AND symb_decoder(16#ef#)) OR
 					(reg_q800 AND symb_decoder(16#0b#)) OR
 					(reg_q800 AND symb_decoder(16#9b#)) OR
 					(reg_q800 AND symb_decoder(16#2f#)) OR
 					(reg_q800 AND symb_decoder(16#a6#)) OR
 					(reg_q800 AND symb_decoder(16#e8#)) OR
 					(reg_q800 AND symb_decoder(16#8f#)) OR
 					(reg_q800 AND symb_decoder(16#40#)) OR
 					(reg_q800 AND symb_decoder(16#8d#)) OR
 					(reg_q800 AND symb_decoder(16#c6#)) OR
 					(reg_q800 AND symb_decoder(16#7f#)) OR
 					(reg_q800 AND symb_decoder(16#22#)) OR
 					(reg_q800 AND symb_decoder(16#58#)) OR
 					(reg_q800 AND symb_decoder(16#44#)) OR
 					(reg_q800 AND symb_decoder(16#18#)) OR
 					(reg_q800 AND symb_decoder(16#b3#)) OR
 					(reg_q800 AND symb_decoder(16#c2#)) OR
 					(reg_q800 AND symb_decoder(16#8c#)) OR
 					(reg_q800 AND symb_decoder(16#59#)) OR
 					(reg_q800 AND symb_decoder(16#e9#)) OR
 					(reg_q800 AND symb_decoder(16#73#)) OR
 					(reg_q800 AND symb_decoder(16#3c#)) OR
 					(reg_q800 AND symb_decoder(16#38#)) OR
 					(reg_q800 AND symb_decoder(16#56#));
reg_q486_in <= (reg_q486 AND symb_decoder(16#39#)) OR
 					(reg_q486 AND symb_decoder(16#37#)) OR
 					(reg_q486 AND symb_decoder(16#38#)) OR
 					(reg_q486 AND symb_decoder(16#33#)) OR
 					(reg_q486 AND symb_decoder(16#34#)) OR
 					(reg_q486 AND symb_decoder(16#31#)) OR
 					(reg_q486 AND symb_decoder(16#35#)) OR
 					(reg_q486 AND symb_decoder(16#32#)) OR
 					(reg_q486 AND symb_decoder(16#30#)) OR
 					(reg_q486 AND symb_decoder(16#36#)) OR
 					(reg_q484 AND symb_decoder(16#32#)) OR
 					(reg_q484 AND symb_decoder(16#33#)) OR
 					(reg_q484 AND symb_decoder(16#30#)) OR
 					(reg_q484 AND symb_decoder(16#34#)) OR
 					(reg_q484 AND symb_decoder(16#36#)) OR
 					(reg_q484 AND symb_decoder(16#37#)) OR
 					(reg_q484 AND symb_decoder(16#31#)) OR
 					(reg_q484 AND symb_decoder(16#39#)) OR
 					(reg_q484 AND symb_decoder(16#38#)) OR
 					(reg_q484 AND symb_decoder(16#35#));
reg_q1757_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q1756 AND symb_decoder(16#0d#)) OR
 					(reg_q1756 AND symb_decoder(16#0a#));
reg_q484_in <= (reg_q494 AND symb_decoder(16#3a#)) OR
 					(reg_q480 AND symb_decoder(16#3a#));
reg_q774_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q773 AND symb_decoder(16#73#)) OR
 					(reg_q773 AND symb_decoder(16#53#));
reg_fullgraph33_init <= "000";

reg_fullgraph33_sel <= "0" & reg_q774_in & reg_q484_in & reg_q1757_in & reg_q486_in & reg_q800_in & reg_q526_in & reg_q395_in;

	--coder fullgraph33
with reg_fullgraph33_sel select
reg_fullgraph33_in <=
	"001" when "00000001",
	"010" when "00000010",
	"011" when "00000100",
	"100" when "00001000",
	"101" when "00010000",
	"110" when "00100000",
	"111" when "01000000",
	"000" when others;
 --end coder

	p_reg_fullgraph33: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph33 <= reg_fullgraph33_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph33 <= reg_fullgraph33_init;
        else
          reg_fullgraph33 <= reg_fullgraph33_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph33

		reg_q395 <= '1' when reg_fullgraph33 = "001" else '0'; 
		reg_q526 <= '1' when reg_fullgraph33 = "010" else '0'; 
		reg_q800 <= '1' when reg_fullgraph33 = "011" else '0'; 
		reg_q486 <= '1' when reg_fullgraph33 = "100" else '0'; 
		reg_q1757 <= '1' when reg_fullgraph33 = "101" else '0'; 
		reg_q484 <= '1' when reg_fullgraph33 = "110" else '0'; 
		reg_q774 <= '1' when reg_fullgraph33 = "111" else '0'; 
--end decoder 

reg_q2677_in <= (reg_q2651 AND symb_decoder(16#dc#)) OR
 					(reg_q2651 AND symb_decoder(16#a6#)) OR
 					(reg_q2651 AND symb_decoder(16#79#)) OR
 					(reg_q2651 AND symb_decoder(16#80#)) OR
 					(reg_q2651 AND symb_decoder(16#a3#)) OR
 					(reg_q2651 AND symb_decoder(16#70#)) OR
 					(reg_q2651 AND symb_decoder(16#26#)) OR
 					(reg_q2651 AND symb_decoder(16#06#)) OR
 					(reg_q2651 AND symb_decoder(16#54#)) OR
 					(reg_q2651 AND symb_decoder(16#86#)) OR
 					(reg_q2651 AND symb_decoder(16#5c#)) OR
 					(reg_q2651 AND symb_decoder(16#0a#)) OR
 					(reg_q2651 AND symb_decoder(16#13#)) OR
 					(reg_q2651 AND symb_decoder(16#66#)) OR
 					(reg_q2651 AND symb_decoder(16#91#)) OR
 					(reg_q2651 AND symb_decoder(16#ac#)) OR
 					(reg_q2651 AND symb_decoder(16#1f#)) OR
 					(reg_q2651 AND symb_decoder(16#a5#)) OR
 					(reg_q2651 AND symb_decoder(16#a2#)) OR
 					(reg_q2651 AND symb_decoder(16#2c#)) OR
 					(reg_q2651 AND symb_decoder(16#3a#)) OR
 					(reg_q2651 AND symb_decoder(16#42#)) OR
 					(reg_q2651 AND symb_decoder(16#9b#)) OR
 					(reg_q2651 AND symb_decoder(16#9d#)) OR
 					(reg_q2651 AND symb_decoder(16#f2#)) OR
 					(reg_q2651 AND symb_decoder(16#5a#)) OR
 					(reg_q2651 AND symb_decoder(16#32#)) OR
 					(reg_q2651 AND symb_decoder(16#76#)) OR
 					(reg_q2651 AND symb_decoder(16#74#)) OR
 					(reg_q2651 AND symb_decoder(16#37#)) OR
 					(reg_q2651 AND symb_decoder(16#f9#)) OR
 					(reg_q2651 AND symb_decoder(16#27#)) OR
 					(reg_q2651 AND symb_decoder(16#3f#)) OR
 					(reg_q2651 AND symb_decoder(16#0b#)) OR
 					(reg_q2651 AND symb_decoder(16#24#)) OR
 					(reg_q2651 AND symb_decoder(16#07#)) OR
 					(reg_q2651 AND symb_decoder(16#fd#)) OR
 					(reg_q2651 AND symb_decoder(16#2f#)) OR
 					(reg_q2651 AND symb_decoder(16#d0#)) OR
 					(reg_q2651 AND symb_decoder(16#c0#)) OR
 					(reg_q2651 AND symb_decoder(16#a4#)) OR
 					(reg_q2651 AND symb_decoder(16#b7#)) OR
 					(reg_q2651 AND symb_decoder(16#a9#)) OR
 					(reg_q2651 AND symb_decoder(16#fc#)) OR
 					(reg_q2651 AND symb_decoder(16#38#)) OR
 					(reg_q2651 AND symb_decoder(16#50#)) OR
 					(reg_q2651 AND symb_decoder(16#5b#)) OR
 					(reg_q2651 AND symb_decoder(16#78#)) OR
 					(reg_q2651 AND symb_decoder(16#8a#)) OR
 					(reg_q2651 AND symb_decoder(16#b4#)) OR
 					(reg_q2651 AND symb_decoder(16#be#)) OR
 					(reg_q2651 AND symb_decoder(16#f1#)) OR
 					(reg_q2651 AND symb_decoder(16#4d#)) OR
 					(reg_q2651 AND symb_decoder(16#11#)) OR
 					(reg_q2651 AND symb_decoder(16#c7#)) OR
 					(reg_q2651 AND symb_decoder(16#12#)) OR
 					(reg_q2651 AND symb_decoder(16#d9#)) OR
 					(reg_q2651 AND symb_decoder(16#a8#)) OR
 					(reg_q2651 AND symb_decoder(16#9f#)) OR
 					(reg_q2651 AND symb_decoder(16#6c#)) OR
 					(reg_q2651 AND symb_decoder(16#41#)) OR
 					(reg_q2651 AND symb_decoder(16#90#)) OR
 					(reg_q2651 AND symb_decoder(16#6d#)) OR
 					(reg_q2651 AND symb_decoder(16#00#)) OR
 					(reg_q2651 AND symb_decoder(16#fa#)) OR
 					(reg_q2651 AND symb_decoder(16#3e#)) OR
 					(reg_q2651 AND symb_decoder(16#89#)) OR
 					(reg_q2651 AND symb_decoder(16#36#)) OR
 					(reg_q2651 AND symb_decoder(16#cd#)) OR
 					(reg_q2651 AND symb_decoder(16#fb#)) OR
 					(reg_q2651 AND symb_decoder(16#eb#)) OR
 					(reg_q2651 AND symb_decoder(16#e9#)) OR
 					(reg_q2651 AND symb_decoder(16#4f#)) OR
 					(reg_q2651 AND symb_decoder(16#cc#)) OR
 					(reg_q2651 AND symb_decoder(16#e5#)) OR
 					(reg_q2651 AND symb_decoder(16#40#)) OR
 					(reg_q2651 AND symb_decoder(16#f4#)) OR
 					(reg_q2651 AND symb_decoder(16#92#)) OR
 					(reg_q2651 AND symb_decoder(16#45#)) OR
 					(reg_q2651 AND symb_decoder(16#96#)) OR
 					(reg_q2651 AND symb_decoder(16#1b#)) OR
 					(reg_q2651 AND symb_decoder(16#01#)) OR
 					(reg_q2651 AND symb_decoder(16#4c#)) OR
 					(reg_q2651 AND symb_decoder(16#4e#)) OR
 					(reg_q2651 AND symb_decoder(16#6e#)) OR
 					(reg_q2651 AND symb_decoder(16#21#)) OR
 					(reg_q2651 AND symb_decoder(16#14#)) OR
 					(reg_q2651 AND symb_decoder(16#87#)) OR
 					(reg_q2651 AND symb_decoder(16#6f#)) OR
 					(reg_q2651 AND symb_decoder(16#71#)) OR
 					(reg_q2651 AND symb_decoder(16#62#)) OR
 					(reg_q2651 AND symb_decoder(16#e3#)) OR
 					(reg_q2651 AND symb_decoder(16#b5#)) OR
 					(reg_q2651 AND symb_decoder(16#49#)) OR
 					(reg_q2651 AND symb_decoder(16#65#)) OR
 					(reg_q2651 AND symb_decoder(16#2e#)) OR
 					(reg_q2651 AND symb_decoder(16#99#)) OR
 					(reg_q2651 AND symb_decoder(16#4b#)) OR
 					(reg_q2651 AND symb_decoder(16#bc#)) OR
 					(reg_q2651 AND symb_decoder(16#48#)) OR
 					(reg_q2651 AND symb_decoder(16#f6#)) OR
 					(reg_q2651 AND symb_decoder(16#e2#)) OR
 					(reg_q2651 AND symb_decoder(16#3c#)) OR
 					(reg_q2651 AND symb_decoder(16#6b#)) OR
 					(reg_q2651 AND symb_decoder(16#db#)) OR
 					(reg_q2651 AND symb_decoder(16#25#)) OR
 					(reg_q2651 AND symb_decoder(16#d4#)) OR
 					(reg_q2651 AND symb_decoder(16#17#)) OR
 					(reg_q2651 AND symb_decoder(16#2d#)) OR
 					(reg_q2651 AND symb_decoder(16#29#)) OR
 					(reg_q2651 AND symb_decoder(16#16#)) OR
 					(reg_q2651 AND symb_decoder(16#08#)) OR
 					(reg_q2651 AND symb_decoder(16#44#)) OR
 					(reg_q2651 AND symb_decoder(16#e8#)) OR
 					(reg_q2651 AND symb_decoder(16#5f#)) OR
 					(reg_q2651 AND symb_decoder(16#c1#)) OR
 					(reg_q2651 AND symb_decoder(16#02#)) OR
 					(reg_q2651 AND symb_decoder(16#7e#)) OR
 					(reg_q2651 AND symb_decoder(16#58#)) OR
 					(reg_q2651 AND symb_decoder(16#7c#)) OR
 					(reg_q2651 AND symb_decoder(16#1e#)) OR
 					(reg_q2651 AND symb_decoder(16#dd#)) OR
 					(reg_q2651 AND symb_decoder(16#f5#)) OR
 					(reg_q2651 AND symb_decoder(16#ee#)) OR
 					(reg_q2651 AND symb_decoder(16#9c#)) OR
 					(reg_q2651 AND symb_decoder(16#04#)) OR
 					(reg_q2651 AND symb_decoder(16#52#)) OR
 					(reg_q2651 AND symb_decoder(16#d5#)) OR
 					(reg_q2651 AND symb_decoder(16#47#)) OR
 					(reg_q2651 AND symb_decoder(16#5e#)) OR
 					(reg_q2651 AND symb_decoder(16#69#)) OR
 					(reg_q2651 AND symb_decoder(16#ba#)) OR
 					(reg_q2651 AND symb_decoder(16#57#)) OR
 					(reg_q2651 AND symb_decoder(16#a1#)) OR
 					(reg_q2651 AND symb_decoder(16#33#)) OR
 					(reg_q2651 AND symb_decoder(16#df#)) OR
 					(reg_q2651 AND symb_decoder(16#18#)) OR
 					(reg_q2651 AND symb_decoder(16#e7#)) OR
 					(reg_q2651 AND symb_decoder(16#d8#)) OR
 					(reg_q2651 AND symb_decoder(16#b8#)) OR
 					(reg_q2651 AND symb_decoder(16#c5#)) OR
 					(reg_q2651 AND symb_decoder(16#c8#)) OR
 					(reg_q2651 AND symb_decoder(16#d2#)) OR
 					(reg_q2651 AND symb_decoder(16#9e#)) OR
 					(reg_q2651 AND symb_decoder(16#ef#)) OR
 					(reg_q2651 AND symb_decoder(16#ce#)) OR
 					(reg_q2651 AND symb_decoder(16#0e#)) OR
 					(reg_q2651 AND symb_decoder(16#56#)) OR
 					(reg_q2651 AND symb_decoder(16#30#)) OR
 					(reg_q2651 AND symb_decoder(16#19#)) OR
 					(reg_q2651 AND symb_decoder(16#ad#)) OR
 					(reg_q2651 AND symb_decoder(16#a7#)) OR
 					(reg_q2651 AND symb_decoder(16#f7#)) OR
 					(reg_q2651 AND symb_decoder(16#b6#)) OR
 					(reg_q2651 AND symb_decoder(16#b0#)) OR
 					(reg_q2651 AND symb_decoder(16#cf#)) OR
 					(reg_q2651 AND symb_decoder(16#f0#)) OR
 					(reg_q2651 AND symb_decoder(16#d6#)) OR
 					(reg_q2651 AND symb_decoder(16#67#)) OR
 					(reg_q2651 AND symb_decoder(16#60#)) OR
 					(reg_q2651 AND symb_decoder(16#15#)) OR
 					(reg_q2651 AND symb_decoder(16#39#)) OR
 					(reg_q2651 AND symb_decoder(16#8e#)) OR
 					(reg_q2651 AND symb_decoder(16#8f#)) OR
 					(reg_q2651 AND symb_decoder(16#ae#)) OR
 					(reg_q2651 AND symb_decoder(16#2b#)) OR
 					(reg_q2651 AND symb_decoder(16#6a#)) OR
 					(reg_q2651 AND symb_decoder(16#a0#)) OR
 					(reg_q2651 AND symb_decoder(16#53#)) OR
 					(reg_q2651 AND symb_decoder(16#e1#)) OR
 					(reg_q2651 AND symb_decoder(16#ff#)) OR
 					(reg_q2651 AND symb_decoder(16#35#)) OR
 					(reg_q2651 AND symb_decoder(16#e6#)) OR
 					(reg_q2651 AND symb_decoder(16#64#)) OR
 					(reg_q2651 AND symb_decoder(16#46#)) OR
 					(reg_q2651 AND symb_decoder(16#8d#)) OR
 					(reg_q2651 AND symb_decoder(16#b9#)) OR
 					(reg_q2651 AND symb_decoder(16#43#)) OR
 					(reg_q2651 AND symb_decoder(16#34#)) OR
 					(reg_q2651 AND symb_decoder(16#23#)) OR
 					(reg_q2651 AND symb_decoder(16#85#)) OR
 					(reg_q2651 AND symb_decoder(16#98#)) OR
 					(reg_q2651 AND symb_decoder(16#97#)) OR
 					(reg_q2651 AND symb_decoder(16#05#)) OR
 					(reg_q2651 AND symb_decoder(16#83#)) OR
 					(reg_q2651 AND symb_decoder(16#81#)) OR
 					(reg_q2651 AND symb_decoder(16#59#)) OR
 					(reg_q2651 AND symb_decoder(16#de#)) OR
 					(reg_q2651 AND symb_decoder(16#4a#)) OR
 					(reg_q2651 AND symb_decoder(16#8c#)) OR
 					(reg_q2651 AND symb_decoder(16#94#)) OR
 					(reg_q2651 AND symb_decoder(16#77#)) OR
 					(reg_q2651 AND symb_decoder(16#3d#)) OR
 					(reg_q2651 AND symb_decoder(16#b2#)) OR
 					(reg_q2651 AND symb_decoder(16#ca#)) OR
 					(reg_q2651 AND symb_decoder(16#61#)) OR
 					(reg_q2651 AND symb_decoder(16#e4#)) OR
 					(reg_q2651 AND symb_decoder(16#d1#)) OR
 					(reg_q2651 AND symb_decoder(16#10#)) OR
 					(reg_q2651 AND symb_decoder(16#ec#)) OR
 					(reg_q2651 AND symb_decoder(16#7a#)) OR
 					(reg_q2651 AND symb_decoder(16#fe#)) OR
 					(reg_q2651 AND symb_decoder(16#cb#)) OR
 					(reg_q2651 AND symb_decoder(16#0d#)) OR
 					(reg_q2651 AND symb_decoder(16#da#)) OR
 					(reg_q2651 AND symb_decoder(16#22#)) OR
 					(reg_q2651 AND symb_decoder(16#51#)) OR
 					(reg_q2651 AND symb_decoder(16#9a#)) OR
 					(reg_q2651 AND symb_decoder(16#09#)) OR
 					(reg_q2651 AND symb_decoder(16#c4#)) OR
 					(reg_q2651 AND symb_decoder(16#ed#)) OR
 					(reg_q2651 AND symb_decoder(16#b3#)) OR
 					(reg_q2651 AND symb_decoder(16#1c#)) OR
 					(reg_q2651 AND symb_decoder(16#95#)) OR
 					(reg_q2651 AND symb_decoder(16#84#)) OR
 					(reg_q2651 AND symb_decoder(16#f8#)) OR
 					(reg_q2651 AND symb_decoder(16#bd#)) OR
 					(reg_q2651 AND symb_decoder(16#88#)) OR
 					(reg_q2651 AND symb_decoder(16#bb#)) OR
 					(reg_q2651 AND symb_decoder(16#bf#)) OR
 					(reg_q2651 AND symb_decoder(16#73#)) OR
 					(reg_q2651 AND symb_decoder(16#c2#)) OR
 					(reg_q2651 AND symb_decoder(16#d7#)) OR
 					(reg_q2651 AND symb_decoder(16#7f#)) OR
 					(reg_q2651 AND symb_decoder(16#c3#)) OR
 					(reg_q2651 AND symb_decoder(16#aa#)) OR
 					(reg_q2651 AND symb_decoder(16#0f#)) OR
 					(reg_q2651 AND symb_decoder(16#20#)) OR
 					(reg_q2651 AND symb_decoder(16#1a#)) OR
 					(reg_q2651 AND symb_decoder(16#68#)) OR
 					(reg_q2651 AND symb_decoder(16#55#)) OR
 					(reg_q2651 AND symb_decoder(16#7d#)) OR
 					(reg_q2651 AND symb_decoder(16#31#)) OR
 					(reg_q2651 AND symb_decoder(16#03#)) OR
 					(reg_q2651 AND symb_decoder(16#f3#)) OR
 					(reg_q2651 AND symb_decoder(16#3b#)) OR
 					(reg_q2651 AND symb_decoder(16#93#)) OR
 					(reg_q2651 AND symb_decoder(16#72#)) OR
 					(reg_q2651 AND symb_decoder(16#ea#)) OR
 					(reg_q2651 AND symb_decoder(16#ab#)) OR
 					(reg_q2651 AND symb_decoder(16#5d#)) OR
 					(reg_q2651 AND symb_decoder(16#c6#)) OR
 					(reg_q2651 AND symb_decoder(16#63#)) OR
 					(reg_q2651 AND symb_decoder(16#1d#)) OR
 					(reg_q2651 AND symb_decoder(16#e0#)) OR
 					(reg_q2651 AND symb_decoder(16#0c#)) OR
 					(reg_q2651 AND symb_decoder(16#75#)) OR
 					(reg_q2651 AND symb_decoder(16#d3#)) OR
 					(reg_q2651 AND symb_decoder(16#8b#)) OR
 					(reg_q2651 AND symb_decoder(16#2a#)) OR
 					(reg_q2651 AND symb_decoder(16#28#)) OR
 					(reg_q2651 AND symb_decoder(16#c9#)) OR
 					(reg_q2651 AND symb_decoder(16#b1#)) OR
 					(reg_q2651 AND symb_decoder(16#7b#)) OR
 					(reg_q2651 AND symb_decoder(16#af#)) OR
 					(reg_q2651 AND symb_decoder(16#82#)) OR
 					(reg_q2677 AND symb_decoder(16#a5#)) OR
 					(reg_q2677 AND symb_decoder(16#79#)) OR
 					(reg_q2677 AND symb_decoder(16#8f#)) OR
 					(reg_q2677 AND symb_decoder(16#13#)) OR
 					(reg_q2677 AND symb_decoder(16#10#)) OR
 					(reg_q2677 AND symb_decoder(16#4f#)) OR
 					(reg_q2677 AND symb_decoder(16#5a#)) OR
 					(reg_q2677 AND symb_decoder(16#1a#)) OR
 					(reg_q2677 AND symb_decoder(16#83#)) OR
 					(reg_q2677 AND symb_decoder(16#7f#)) OR
 					(reg_q2677 AND symb_decoder(16#e3#)) OR
 					(reg_q2677 AND symb_decoder(16#64#)) OR
 					(reg_q2677 AND symb_decoder(16#c8#)) OR
 					(reg_q2677 AND symb_decoder(16#94#)) OR
 					(reg_q2677 AND symb_decoder(16#d2#)) OR
 					(reg_q2677 AND symb_decoder(16#80#)) OR
 					(reg_q2677 AND symb_decoder(16#38#)) OR
 					(reg_q2677 AND symb_decoder(16#f7#)) OR
 					(reg_q2677 AND symb_decoder(16#ad#)) OR
 					(reg_q2677 AND symb_decoder(16#54#)) OR
 					(reg_q2677 AND symb_decoder(16#d8#)) OR
 					(reg_q2677 AND symb_decoder(16#15#)) OR
 					(reg_q2677 AND symb_decoder(16#43#)) OR
 					(reg_q2677 AND symb_decoder(16#3d#)) OR
 					(reg_q2677 AND symb_decoder(16#9a#)) OR
 					(reg_q2677 AND symb_decoder(16#6b#)) OR
 					(reg_q2677 AND symb_decoder(16#01#)) OR
 					(reg_q2677 AND symb_decoder(16#e0#)) OR
 					(reg_q2677 AND symb_decoder(16#bf#)) OR
 					(reg_q2677 AND symb_decoder(16#08#)) OR
 					(reg_q2677 AND symb_decoder(16#cb#)) OR
 					(reg_q2677 AND symb_decoder(16#2d#)) OR
 					(reg_q2677 AND symb_decoder(16#c7#)) OR
 					(reg_q2677 AND symb_decoder(16#41#)) OR
 					(reg_q2677 AND symb_decoder(16#74#)) OR
 					(reg_q2677 AND symb_decoder(16#02#)) OR
 					(reg_q2677 AND symb_decoder(16#1c#)) OR
 					(reg_q2677 AND symb_decoder(16#c5#)) OR
 					(reg_q2677 AND symb_decoder(16#20#)) OR
 					(reg_q2677 AND symb_decoder(16#5d#)) OR
 					(reg_q2677 AND symb_decoder(16#cf#)) OR
 					(reg_q2677 AND symb_decoder(16#89#)) OR
 					(reg_q2677 AND symb_decoder(16#0f#)) OR
 					(reg_q2677 AND symb_decoder(16#b0#)) OR
 					(reg_q2677 AND symb_decoder(16#a9#)) OR
 					(reg_q2677 AND symb_decoder(16#d0#)) OR
 					(reg_q2677 AND symb_decoder(16#29#)) OR
 					(reg_q2677 AND symb_decoder(16#0a#)) OR
 					(reg_q2677 AND symb_decoder(16#b5#)) OR
 					(reg_q2677 AND symb_decoder(16#44#)) OR
 					(reg_q2677 AND symb_decoder(16#d9#)) OR
 					(reg_q2677 AND symb_decoder(16#ed#)) OR
 					(reg_q2677 AND symb_decoder(16#9b#)) OR
 					(reg_q2677 AND symb_decoder(16#d1#)) OR
 					(reg_q2677 AND symb_decoder(16#5b#)) OR
 					(reg_q2677 AND symb_decoder(16#46#)) OR
 					(reg_q2677 AND symb_decoder(16#50#)) OR
 					(reg_q2677 AND symb_decoder(16#d6#)) OR
 					(reg_q2677 AND symb_decoder(16#3a#)) OR
 					(reg_q2677 AND symb_decoder(16#28#)) OR
 					(reg_q2677 AND symb_decoder(16#66#)) OR
 					(reg_q2677 AND symb_decoder(16#f6#)) OR
 					(reg_q2677 AND symb_decoder(16#55#)) OR
 					(reg_q2677 AND symb_decoder(16#26#)) OR
 					(reg_q2677 AND symb_decoder(16#bc#)) OR
 					(reg_q2677 AND symb_decoder(16#e7#)) OR
 					(reg_q2677 AND symb_decoder(16#95#)) OR
 					(reg_q2677 AND symb_decoder(16#9f#)) OR
 					(reg_q2677 AND symb_decoder(16#47#)) OR
 					(reg_q2677 AND symb_decoder(16#b3#)) OR
 					(reg_q2677 AND symb_decoder(16#33#)) OR
 					(reg_q2677 AND symb_decoder(16#c3#)) OR
 					(reg_q2677 AND symb_decoder(16#05#)) OR
 					(reg_q2677 AND symb_decoder(16#3f#)) OR
 					(reg_q2677 AND symb_decoder(16#00#)) OR
 					(reg_q2677 AND symb_decoder(16#60#)) OR
 					(reg_q2677 AND symb_decoder(16#7b#)) OR
 					(reg_q2677 AND symb_decoder(16#8b#)) OR
 					(reg_q2677 AND symb_decoder(16#45#)) OR
 					(reg_q2677 AND symb_decoder(16#9c#)) OR
 					(reg_q2677 AND symb_decoder(16#04#)) OR
 					(reg_q2677 AND symb_decoder(16#75#)) OR
 					(reg_q2677 AND symb_decoder(16#63#)) OR
 					(reg_q2677 AND symb_decoder(16#49#)) OR
 					(reg_q2677 AND symb_decoder(16#6e#)) OR
 					(reg_q2677 AND symb_decoder(16#51#)) OR
 					(reg_q2677 AND symb_decoder(16#4e#)) OR
 					(reg_q2677 AND symb_decoder(16#f1#)) OR
 					(reg_q2677 AND symb_decoder(16#fb#)) OR
 					(reg_q2677 AND symb_decoder(16#be#)) OR
 					(reg_q2677 AND symb_decoder(16#57#)) OR
 					(reg_q2677 AND symb_decoder(16#71#)) OR
 					(reg_q2677 AND symb_decoder(16#2a#)) OR
 					(reg_q2677 AND symb_decoder(16#ee#)) OR
 					(reg_q2677 AND symb_decoder(16#96#)) OR
 					(reg_q2677 AND symb_decoder(16#48#)) OR
 					(reg_q2677 AND symb_decoder(16#69#)) OR
 					(reg_q2677 AND symb_decoder(16#30#)) OR
 					(reg_q2677 AND symb_decoder(16#81#)) OR
 					(reg_q2677 AND symb_decoder(16#12#)) OR
 					(reg_q2677 AND symb_decoder(16#c6#)) OR
 					(reg_q2677 AND symb_decoder(16#85#)) OR
 					(reg_q2677 AND symb_decoder(16#03#)) OR
 					(reg_q2677 AND symb_decoder(16#70#)) OR
 					(reg_q2677 AND symb_decoder(16#a8#)) OR
 					(reg_q2677 AND symb_decoder(16#24#)) OR
 					(reg_q2677 AND symb_decoder(16#a4#)) OR
 					(reg_q2677 AND symb_decoder(16#21#)) OR
 					(reg_q2677 AND symb_decoder(16#aa#)) OR
 					(reg_q2677 AND symb_decoder(16#e8#)) OR
 					(reg_q2677 AND symb_decoder(16#0d#)) OR
 					(reg_q2677 AND symb_decoder(16#cd#)) OR
 					(reg_q2677 AND symb_decoder(16#ab#)) OR
 					(reg_q2677 AND symb_decoder(16#23#)) OR
 					(reg_q2677 AND symb_decoder(16#58#)) OR
 					(reg_q2677 AND symb_decoder(16#f3#)) OR
 					(reg_q2677 AND symb_decoder(16#35#)) OR
 					(reg_q2677 AND symb_decoder(16#82#)) OR
 					(reg_q2677 AND symb_decoder(16#93#)) OR
 					(reg_q2677 AND symb_decoder(16#d4#)) OR
 					(reg_q2677 AND symb_decoder(16#76#)) OR
 					(reg_q2677 AND symb_decoder(16#67#)) OR
 					(reg_q2677 AND symb_decoder(16#53#)) OR
 					(reg_q2677 AND symb_decoder(16#1d#)) OR
 					(reg_q2677 AND symb_decoder(16#bb#)) OR
 					(reg_q2677 AND symb_decoder(16#7d#)) OR
 					(reg_q2677 AND symb_decoder(16#73#)) OR
 					(reg_q2677 AND symb_decoder(16#17#)) OR
 					(reg_q2677 AND symb_decoder(16#32#)) OR
 					(reg_q2677 AND symb_decoder(16#b6#)) OR
 					(reg_q2677 AND symb_decoder(16#fd#)) OR
 					(reg_q2677 AND symb_decoder(16#91#)) OR
 					(reg_q2677 AND symb_decoder(16#b7#)) OR
 					(reg_q2677 AND symb_decoder(16#39#)) OR
 					(reg_q2677 AND symb_decoder(16#ba#)) OR
 					(reg_q2677 AND symb_decoder(16#34#)) OR
 					(reg_q2677 AND symb_decoder(16#98#)) OR
 					(reg_q2677 AND symb_decoder(16#2e#)) OR
 					(reg_q2677 AND symb_decoder(16#df#)) OR
 					(reg_q2677 AND symb_decoder(16#87#)) OR
 					(reg_q2677 AND symb_decoder(16#2b#)) OR
 					(reg_q2677 AND symb_decoder(16#d7#)) OR
 					(reg_q2677 AND symb_decoder(16#ce#)) OR
 					(reg_q2677 AND symb_decoder(16#90#)) OR
 					(reg_q2677 AND symb_decoder(16#7a#)) OR
 					(reg_q2677 AND symb_decoder(16#14#)) OR
 					(reg_q2677 AND symb_decoder(16#6d#)) OR
 					(reg_q2677 AND symb_decoder(16#f2#)) OR
 					(reg_q2677 AND symb_decoder(16#2c#)) OR
 					(reg_q2677 AND symb_decoder(16#16#)) OR
 					(reg_q2677 AND symb_decoder(16#dd#)) OR
 					(reg_q2677 AND symb_decoder(16#0c#)) OR
 					(reg_q2677 AND symb_decoder(16#52#)) OR
 					(reg_q2677 AND symb_decoder(16#3e#)) OR
 					(reg_q2677 AND symb_decoder(16#40#)) OR
 					(reg_q2677 AND symb_decoder(16#b1#)) OR
 					(reg_q2677 AND symb_decoder(16#fc#)) OR
 					(reg_q2677 AND symb_decoder(16#e5#)) OR
 					(reg_q2677 AND symb_decoder(16#b9#)) OR
 					(reg_q2677 AND symb_decoder(16#42#)) OR
 					(reg_q2677 AND symb_decoder(16#e2#)) OR
 					(reg_q2677 AND symb_decoder(16#1f#)) OR
 					(reg_q2677 AND symb_decoder(16#d5#)) OR
 					(reg_q2677 AND symb_decoder(16#f0#)) OR
 					(reg_q2677 AND symb_decoder(16#4a#)) OR
 					(reg_q2677 AND symb_decoder(16#8a#)) OR
 					(reg_q2677 AND symb_decoder(16#07#)) OR
 					(reg_q2677 AND symb_decoder(16#6c#)) OR
 					(reg_q2677 AND symb_decoder(16#7c#)) OR
 					(reg_q2677 AND symb_decoder(16#86#)) OR
 					(reg_q2677 AND symb_decoder(16#c4#)) OR
 					(reg_q2677 AND symb_decoder(16#37#)) OR
 					(reg_q2677 AND symb_decoder(16#4d#)) OR
 					(reg_q2677 AND symb_decoder(16#25#)) OR
 					(reg_q2677 AND symb_decoder(16#0b#)) OR
 					(reg_q2677 AND symb_decoder(16#8e#)) OR
 					(reg_q2677 AND symb_decoder(16#68#)) OR
 					(reg_q2677 AND symb_decoder(16#ca#)) OR
 					(reg_q2677 AND symb_decoder(16#a2#)) OR
 					(reg_q2677 AND symb_decoder(16#5c#)) OR
 					(reg_q2677 AND symb_decoder(16#3c#)) OR
 					(reg_q2677 AND symb_decoder(16#36#)) OR
 					(reg_q2677 AND symb_decoder(16#e4#)) OR
 					(reg_q2677 AND symb_decoder(16#56#)) OR
 					(reg_q2677 AND symb_decoder(16#b2#)) OR
 					(reg_q2677 AND symb_decoder(16#f4#)) OR
 					(reg_q2677 AND symb_decoder(16#b8#)) OR
 					(reg_q2677 AND symb_decoder(16#97#)) OR
 					(reg_q2677 AND symb_decoder(16#ea#)) OR
 					(reg_q2677 AND symb_decoder(16#4c#)) OR
 					(reg_q2677 AND symb_decoder(16#f9#)) OR
 					(reg_q2677 AND symb_decoder(16#a3#)) OR
 					(reg_q2677 AND symb_decoder(16#65#)) OR
 					(reg_q2677 AND symb_decoder(16#62#)) OR
 					(reg_q2677 AND symb_decoder(16#72#)) OR
 					(reg_q2677 AND symb_decoder(16#c1#)) OR
 					(reg_q2677 AND symb_decoder(16#fe#)) OR
 					(reg_q2677 AND symb_decoder(16#31#)) OR
 					(reg_q2677 AND symb_decoder(16#99#)) OR
 					(reg_q2677 AND symb_decoder(16#de#)) OR
 					(reg_q2677 AND symb_decoder(16#88#)) OR
 					(reg_q2677 AND symb_decoder(16#ef#)) OR
 					(reg_q2677 AND symb_decoder(16#ac#)) OR
 					(reg_q2677 AND symb_decoder(16#b4#)) OR
 					(reg_q2677 AND symb_decoder(16#5f#)) OR
 					(reg_q2677 AND symb_decoder(16#06#)) OR
 					(reg_q2677 AND symb_decoder(16#fa#)) OR
 					(reg_q2677 AND symb_decoder(16#9d#)) OR
 					(reg_q2677 AND symb_decoder(16#61#)) OR
 					(reg_q2677 AND symb_decoder(16#8c#)) OR
 					(reg_q2677 AND symb_decoder(16#09#)) OR
 					(reg_q2677 AND symb_decoder(16#1e#)) OR
 					(reg_q2677 AND symb_decoder(16#e1#)) OR
 					(reg_q2677 AND symb_decoder(16#a7#)) OR
 					(reg_q2677 AND symb_decoder(16#a6#)) OR
 					(reg_q2677 AND symb_decoder(16#2f#)) OR
 					(reg_q2677 AND symb_decoder(16#6a#)) OR
 					(reg_q2677 AND symb_decoder(16#d3#)) OR
 					(reg_q2677 AND symb_decoder(16#ec#)) OR
 					(reg_q2677 AND symb_decoder(16#cc#)) OR
 					(reg_q2677 AND symb_decoder(16#22#)) OR
 					(reg_q2677 AND symb_decoder(16#9e#)) OR
 					(reg_q2677 AND symb_decoder(16#18#)) OR
 					(reg_q2677 AND symb_decoder(16#11#)) OR
 					(reg_q2677 AND symb_decoder(16#af#)) OR
 					(reg_q2677 AND symb_decoder(16#a0#)) OR
 					(reg_q2677 AND symb_decoder(16#a1#)) OR
 					(reg_q2677 AND symb_decoder(16#78#)) OR
 					(reg_q2677 AND symb_decoder(16#5e#)) OR
 					(reg_q2677 AND symb_decoder(16#7e#)) OR
 					(reg_q2677 AND symb_decoder(16#f8#)) OR
 					(reg_q2677 AND symb_decoder(16#8d#)) OR
 					(reg_q2677 AND symb_decoder(16#bd#)) OR
 					(reg_q2677 AND symb_decoder(16#3b#)) OR
 					(reg_q2677 AND symb_decoder(16#59#)) OR
 					(reg_q2677 AND symb_decoder(16#da#)) OR
 					(reg_q2677 AND symb_decoder(16#ae#)) OR
 					(reg_q2677 AND symb_decoder(16#e9#)) OR
 					(reg_q2677 AND symb_decoder(16#c9#)) OR
 					(reg_q2677 AND symb_decoder(16#f5#)) OR
 					(reg_q2677 AND symb_decoder(16#77#)) OR
 					(reg_q2677 AND symb_decoder(16#c2#)) OR
 					(reg_q2677 AND symb_decoder(16#db#)) OR
 					(reg_q2677 AND symb_decoder(16#e6#)) OR
 					(reg_q2677 AND symb_decoder(16#1b#)) OR
 					(reg_q2677 AND symb_decoder(16#dc#)) OR
 					(reg_q2677 AND symb_decoder(16#c0#)) OR
 					(reg_q2677 AND symb_decoder(16#eb#)) OR
 					(reg_q2677 AND symb_decoder(16#6f#)) OR
 					(reg_q2677 AND symb_decoder(16#27#)) OR
 					(reg_q2677 AND symb_decoder(16#4b#)) OR
 					(reg_q2677 AND symb_decoder(16#84#)) OR
 					(reg_q2677 AND symb_decoder(16#19#)) OR
 					(reg_q2677 AND symb_decoder(16#0e#)) OR
 					(reg_q2677 AND symb_decoder(16#ff#)) OR
 					(reg_q2677 AND symb_decoder(16#92#));
reg_q2677_init <= '0' ;
	p_reg_q2677: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2677 <= reg_q2677_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2677 <= reg_q2677_init;
        else
          reg_q2677 <= reg_q2677_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1145_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1145 AND symb_decoder(16#ba#)) OR
 					(reg_q1145 AND symb_decoder(16#c3#)) OR
 					(reg_q1145 AND symb_decoder(16#73#)) OR
 					(reg_q1145 AND symb_decoder(16#2a#)) OR
 					(reg_q1145 AND symb_decoder(16#cd#)) OR
 					(reg_q1145 AND symb_decoder(16#da#)) OR
 					(reg_q1145 AND symb_decoder(16#31#)) OR
 					(reg_q1145 AND symb_decoder(16#f8#)) OR
 					(reg_q1145 AND symb_decoder(16#b7#)) OR
 					(reg_q1145 AND symb_decoder(16#ef#)) OR
 					(reg_q1145 AND symb_decoder(16#63#)) OR
 					(reg_q1145 AND symb_decoder(16#3b#)) OR
 					(reg_q1145 AND symb_decoder(16#aa#)) OR
 					(reg_q1145 AND symb_decoder(16#0a#)) OR
 					(reg_q1145 AND symb_decoder(16#48#)) OR
 					(reg_q1145 AND symb_decoder(16#03#)) OR
 					(reg_q1145 AND symb_decoder(16#25#)) OR
 					(reg_q1145 AND symb_decoder(16#b1#)) OR
 					(reg_q1145 AND symb_decoder(16#4e#)) OR
 					(reg_q1145 AND symb_decoder(16#4a#)) OR
 					(reg_q1145 AND symb_decoder(16#72#)) OR
 					(reg_q1145 AND symb_decoder(16#93#)) OR
 					(reg_q1145 AND symb_decoder(16#0d#)) OR
 					(reg_q1145 AND symb_decoder(16#ae#)) OR
 					(reg_q1145 AND symb_decoder(16#05#)) OR
 					(reg_q1145 AND symb_decoder(16#d0#)) OR
 					(reg_q1145 AND symb_decoder(16#54#)) OR
 					(reg_q1145 AND symb_decoder(16#1c#)) OR
 					(reg_q1145 AND symb_decoder(16#ea#)) OR
 					(reg_q1145 AND symb_decoder(16#b9#)) OR
 					(reg_q1145 AND symb_decoder(16#a3#)) OR
 					(reg_q1145 AND symb_decoder(16#e0#)) OR
 					(reg_q1145 AND symb_decoder(16#b2#)) OR
 					(reg_q1145 AND symb_decoder(16#49#)) OR
 					(reg_q1145 AND symb_decoder(16#0b#)) OR
 					(reg_q1145 AND symb_decoder(16#1e#)) OR
 					(reg_q1145 AND symb_decoder(16#74#)) OR
 					(reg_q1145 AND symb_decoder(16#83#)) OR
 					(reg_q1145 AND symb_decoder(16#b8#)) OR
 					(reg_q1145 AND symb_decoder(16#0e#)) OR
 					(reg_q1145 AND symb_decoder(16#f9#)) OR
 					(reg_q1145 AND symb_decoder(16#90#)) OR
 					(reg_q1145 AND symb_decoder(16#bb#)) OR
 					(reg_q1145 AND symb_decoder(16#61#)) OR
 					(reg_q1145 AND symb_decoder(16#4f#)) OR
 					(reg_q1145 AND symb_decoder(16#08#)) OR
 					(reg_q1145 AND symb_decoder(16#fd#)) OR
 					(reg_q1145 AND symb_decoder(16#b3#)) OR
 					(reg_q1145 AND symb_decoder(16#f1#)) OR
 					(reg_q1145 AND symb_decoder(16#bf#)) OR
 					(reg_q1145 AND symb_decoder(16#29#)) OR
 					(reg_q1145 AND symb_decoder(16#43#)) OR
 					(reg_q1145 AND symb_decoder(16#e9#)) OR
 					(reg_q1145 AND symb_decoder(16#38#)) OR
 					(reg_q1145 AND symb_decoder(16#c6#)) OR
 					(reg_q1145 AND symb_decoder(16#23#)) OR
 					(reg_q1145 AND symb_decoder(16#6c#)) OR
 					(reg_q1145 AND symb_decoder(16#32#)) OR
 					(reg_q1145 AND symb_decoder(16#1a#)) OR
 					(reg_q1145 AND symb_decoder(16#e1#)) OR
 					(reg_q1145 AND symb_decoder(16#7d#)) OR
 					(reg_q1145 AND symb_decoder(16#9d#)) OR
 					(reg_q1145 AND symb_decoder(16#9c#)) OR
 					(reg_q1145 AND symb_decoder(16#55#)) OR
 					(reg_q1145 AND symb_decoder(16#5f#)) OR
 					(reg_q1145 AND symb_decoder(16#dc#)) OR
 					(reg_q1145 AND symb_decoder(16#01#)) OR
 					(reg_q1145 AND symb_decoder(16#3a#)) OR
 					(reg_q1145 AND symb_decoder(16#d3#)) OR
 					(reg_q1145 AND symb_decoder(16#ee#)) OR
 					(reg_q1145 AND symb_decoder(16#db#)) OR
 					(reg_q1145 AND symb_decoder(16#84#)) OR
 					(reg_q1145 AND symb_decoder(16#8e#)) OR
 					(reg_q1145 AND symb_decoder(16#9a#)) OR
 					(reg_q1145 AND symb_decoder(16#1f#)) OR
 					(reg_q1145 AND symb_decoder(16#d9#)) OR
 					(reg_q1145 AND symb_decoder(16#fb#)) OR
 					(reg_q1145 AND symb_decoder(16#a6#)) OR
 					(reg_q1145 AND symb_decoder(16#24#)) OR
 					(reg_q1145 AND symb_decoder(16#ce#)) OR
 					(reg_q1145 AND symb_decoder(16#7a#)) OR
 					(reg_q1145 AND symb_decoder(16#47#)) OR
 					(reg_q1145 AND symb_decoder(16#91#)) OR
 					(reg_q1145 AND symb_decoder(16#ec#)) OR
 					(reg_q1145 AND symb_decoder(16#16#)) OR
 					(reg_q1145 AND symb_decoder(16#6a#)) OR
 					(reg_q1145 AND symb_decoder(16#a2#)) OR
 					(reg_q1145 AND symb_decoder(16#66#)) OR
 					(reg_q1145 AND symb_decoder(16#6f#)) OR
 					(reg_q1145 AND symb_decoder(16#6b#)) OR
 					(reg_q1145 AND symb_decoder(16#36#)) OR
 					(reg_q1145 AND symb_decoder(16#8c#)) OR
 					(reg_q1145 AND symb_decoder(16#79#)) OR
 					(reg_q1145 AND symb_decoder(16#cc#)) OR
 					(reg_q1145 AND symb_decoder(16#57#)) OR
 					(reg_q1145 AND symb_decoder(16#a9#)) OR
 					(reg_q1145 AND symb_decoder(16#69#)) OR
 					(reg_q1145 AND symb_decoder(16#e8#)) OR
 					(reg_q1145 AND symb_decoder(16#c8#)) OR
 					(reg_q1145 AND symb_decoder(16#d1#)) OR
 					(reg_q1145 AND symb_decoder(16#33#)) OR
 					(reg_q1145 AND symb_decoder(16#bd#)) OR
 					(reg_q1145 AND symb_decoder(16#c9#)) OR
 					(reg_q1145 AND symb_decoder(16#0f#)) OR
 					(reg_q1145 AND symb_decoder(16#71#)) OR
 					(reg_q1145 AND symb_decoder(16#60#)) OR
 					(reg_q1145 AND symb_decoder(16#9b#)) OR
 					(reg_q1145 AND symb_decoder(16#dd#)) OR
 					(reg_q1145 AND symb_decoder(16#a0#)) OR
 					(reg_q1145 AND symb_decoder(16#e5#)) OR
 					(reg_q1145 AND symb_decoder(16#2c#)) OR
 					(reg_q1145 AND symb_decoder(16#67#)) OR
 					(reg_q1145 AND symb_decoder(16#5a#)) OR
 					(reg_q1145 AND symb_decoder(16#78#)) OR
 					(reg_q1145 AND symb_decoder(16#3c#)) OR
 					(reg_q1145 AND symb_decoder(16#56#)) OR
 					(reg_q1145 AND symb_decoder(16#40#)) OR
 					(reg_q1145 AND symb_decoder(16#51#)) OR
 					(reg_q1145 AND symb_decoder(16#15#)) OR
 					(reg_q1145 AND symb_decoder(16#e6#)) OR
 					(reg_q1145 AND symb_decoder(16#19#)) OR
 					(reg_q1145 AND symb_decoder(16#6d#)) OR
 					(reg_q1145 AND symb_decoder(16#42#)) OR
 					(reg_q1145 AND symb_decoder(16#e4#)) OR
 					(reg_q1145 AND symb_decoder(16#50#)) OR
 					(reg_q1145 AND symb_decoder(16#22#)) OR
 					(reg_q1145 AND symb_decoder(16#2f#)) OR
 					(reg_q1145 AND symb_decoder(16#52#)) OR
 					(reg_q1145 AND symb_decoder(16#30#)) OR
 					(reg_q1145 AND symb_decoder(16#04#)) OR
 					(reg_q1145 AND symb_decoder(16#2d#)) OR
 					(reg_q1145 AND symb_decoder(16#70#)) OR
 					(reg_q1145 AND symb_decoder(16#e3#)) OR
 					(reg_q1145 AND symb_decoder(16#7b#)) OR
 					(reg_q1145 AND symb_decoder(16#d8#)) OR
 					(reg_q1145 AND symb_decoder(16#df#)) OR
 					(reg_q1145 AND symb_decoder(16#28#)) OR
 					(reg_q1145 AND symb_decoder(16#a7#)) OR
 					(reg_q1145 AND symb_decoder(16#a8#)) OR
 					(reg_q1145 AND symb_decoder(16#f3#)) OR
 					(reg_q1145 AND symb_decoder(16#81#)) OR
 					(reg_q1145 AND symb_decoder(16#9e#)) OR
 					(reg_q1145 AND symb_decoder(16#5e#)) OR
 					(reg_q1145 AND symb_decoder(16#86#)) OR
 					(reg_q1145 AND symb_decoder(16#76#)) OR
 					(reg_q1145 AND symb_decoder(16#27#)) OR
 					(reg_q1145 AND symb_decoder(16#37#)) OR
 					(reg_q1145 AND symb_decoder(16#c4#)) OR
 					(reg_q1145 AND symb_decoder(16#f6#)) OR
 					(reg_q1145 AND symb_decoder(16#d4#)) OR
 					(reg_q1145 AND symb_decoder(16#88#)) OR
 					(reg_q1145 AND symb_decoder(16#8b#)) OR
 					(reg_q1145 AND symb_decoder(16#ff#)) OR
 					(reg_q1145 AND symb_decoder(16#f0#)) OR
 					(reg_q1145 AND symb_decoder(16#2b#)) OR
 					(reg_q1145 AND symb_decoder(16#b5#)) OR
 					(reg_q1145 AND symb_decoder(16#a4#)) OR
 					(reg_q1145 AND symb_decoder(16#80#)) OR
 					(reg_q1145 AND symb_decoder(16#09#)) OR
 					(reg_q1145 AND symb_decoder(16#b0#)) OR
 					(reg_q1145 AND symb_decoder(16#2e#)) OR
 					(reg_q1145 AND symb_decoder(16#c7#)) OR
 					(reg_q1145 AND symb_decoder(16#34#)) OR
 					(reg_q1145 AND symb_decoder(16#d5#)) OR
 					(reg_q1145 AND symb_decoder(16#8a#)) OR
 					(reg_q1145 AND symb_decoder(16#4c#)) OR
 					(reg_q1145 AND symb_decoder(16#82#)) OR
 					(reg_q1145 AND symb_decoder(16#53#)) OR
 					(reg_q1145 AND symb_decoder(16#1d#)) OR
 					(reg_q1145 AND symb_decoder(16#bc#)) OR
 					(reg_q1145 AND symb_decoder(16#44#)) OR
 					(reg_q1145 AND symb_decoder(16#c2#)) OR
 					(reg_q1145 AND symb_decoder(16#45#)) OR
 					(reg_q1145 AND symb_decoder(16#fc#)) OR
 					(reg_q1145 AND symb_decoder(16#c1#)) OR
 					(reg_q1145 AND symb_decoder(16#c0#)) OR
 					(reg_q1145 AND symb_decoder(16#12#)) OR
 					(reg_q1145 AND symb_decoder(16#5d#)) OR
 					(reg_q1145 AND symb_decoder(16#4d#)) OR
 					(reg_q1145 AND symb_decoder(16#68#)) OR
 					(reg_q1145 AND symb_decoder(16#9f#)) OR
 					(reg_q1145 AND symb_decoder(16#26#)) OR
 					(reg_q1145 AND symb_decoder(16#b6#)) OR
 					(reg_q1145 AND symb_decoder(16#99#)) OR
 					(reg_q1145 AND symb_decoder(16#07#)) OR
 					(reg_q1145 AND symb_decoder(16#fa#)) OR
 					(reg_q1145 AND symb_decoder(16#8f#)) OR
 					(reg_q1145 AND symb_decoder(16#ac#)) OR
 					(reg_q1145 AND symb_decoder(16#97#)) OR
 					(reg_q1145 AND symb_decoder(16#ca#)) OR
 					(reg_q1145 AND symb_decoder(16#21#)) OR
 					(reg_q1145 AND symb_decoder(16#1b#)) OR
 					(reg_q1145 AND symb_decoder(16#00#)) OR
 					(reg_q1145 AND symb_decoder(16#cb#)) OR
 					(reg_q1145 AND symb_decoder(16#13#)) OR
 					(reg_q1145 AND symb_decoder(16#85#)) OR
 					(reg_q1145 AND symb_decoder(16#87#)) OR
 					(reg_q1145 AND symb_decoder(16#59#)) OR
 					(reg_q1145 AND symb_decoder(16#62#)) OR
 					(reg_q1145 AND symb_decoder(16#ab#)) OR
 					(reg_q1145 AND symb_decoder(16#92#)) OR
 					(reg_q1145 AND symb_decoder(16#3f#)) OR
 					(reg_q1145 AND symb_decoder(16#5c#)) OR
 					(reg_q1145 AND symb_decoder(16#3e#)) OR
 					(reg_q1145 AND symb_decoder(16#06#)) OR
 					(reg_q1145 AND symb_decoder(16#f7#)) OR
 					(reg_q1145 AND symb_decoder(16#96#)) OR
 					(reg_q1145 AND symb_decoder(16#e2#)) OR
 					(reg_q1145 AND symb_decoder(16#d2#)) OR
 					(reg_q1145 AND symb_decoder(16#7e#)) OR
 					(reg_q1145 AND symb_decoder(16#7f#)) OR
 					(reg_q1145 AND symb_decoder(16#a1#)) OR
 					(reg_q1145 AND symb_decoder(16#20#)) OR
 					(reg_q1145 AND symb_decoder(16#f4#)) OR
 					(reg_q1145 AND symb_decoder(16#0c#)) OR
 					(reg_q1145 AND symb_decoder(16#de#)) OR
 					(reg_q1145 AND symb_decoder(16#c5#)) OR
 					(reg_q1145 AND symb_decoder(16#ad#)) OR
 					(reg_q1145 AND symb_decoder(16#64#)) OR
 					(reg_q1145 AND symb_decoder(16#eb#)) OR
 					(reg_q1145 AND symb_decoder(16#10#)) OR
 					(reg_q1145 AND symb_decoder(16#02#)) OR
 					(reg_q1145 AND symb_decoder(16#95#)) OR
 					(reg_q1145 AND symb_decoder(16#fe#)) OR
 					(reg_q1145 AND symb_decoder(16#17#)) OR
 					(reg_q1145 AND symb_decoder(16#3d#)) OR
 					(reg_q1145 AND symb_decoder(16#75#)) OR
 					(reg_q1145 AND symb_decoder(16#39#)) OR
 					(reg_q1145 AND symb_decoder(16#18#)) OR
 					(reg_q1145 AND symb_decoder(16#6e#)) OR
 					(reg_q1145 AND symb_decoder(16#ed#)) OR
 					(reg_q1145 AND symb_decoder(16#5b#)) OR
 					(reg_q1145 AND symb_decoder(16#af#)) OR
 					(reg_q1145 AND symb_decoder(16#f2#)) OR
 					(reg_q1145 AND symb_decoder(16#be#)) OR
 					(reg_q1145 AND symb_decoder(16#77#)) OR
 					(reg_q1145 AND symb_decoder(16#35#)) OR
 					(reg_q1145 AND symb_decoder(16#e7#)) OR
 					(reg_q1145 AND symb_decoder(16#a5#)) OR
 					(reg_q1145 AND symb_decoder(16#89#)) OR
 					(reg_q1145 AND symb_decoder(16#58#)) OR
 					(reg_q1145 AND symb_decoder(16#11#)) OR
 					(reg_q1145 AND symb_decoder(16#8d#)) OR
 					(reg_q1145 AND symb_decoder(16#41#)) OR
 					(reg_q1145 AND symb_decoder(16#f5#)) OR
 					(reg_q1145 AND symb_decoder(16#d6#)) OR
 					(reg_q1145 AND symb_decoder(16#14#)) OR
 					(reg_q1145 AND symb_decoder(16#65#)) OR
 					(reg_q1145 AND symb_decoder(16#98#)) OR
 					(reg_q1145 AND symb_decoder(16#cf#)) OR
 					(reg_q1145 AND symb_decoder(16#4b#)) OR
 					(reg_q1145 AND symb_decoder(16#94#)) OR
 					(reg_q1145 AND symb_decoder(16#7c#)) OR
 					(reg_q1145 AND symb_decoder(16#d7#)) OR
 					(reg_q1145 AND symb_decoder(16#b4#)) OR
 					(reg_q1145 AND symb_decoder(16#46#));
reg_q1145_init <= '0' ;
	p_reg_q1145: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1145 <= reg_q1145_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1145 <= reg_q1145_init;
        else
          reg_q1145 <= reg_q1145_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q133_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q133 AND symb_decoder(16#0e#)) OR
 					(reg_q133 AND symb_decoder(16#11#)) OR
 					(reg_q133 AND symb_decoder(16#f6#)) OR
 					(reg_q133 AND symb_decoder(16#bb#)) OR
 					(reg_q133 AND symb_decoder(16#ca#)) OR
 					(reg_q133 AND symb_decoder(16#25#)) OR
 					(reg_q133 AND symb_decoder(16#c2#)) OR
 					(reg_q133 AND symb_decoder(16#4e#)) OR
 					(reg_q133 AND symb_decoder(16#96#)) OR
 					(reg_q133 AND symb_decoder(16#b7#)) OR
 					(reg_q133 AND symb_decoder(16#22#)) OR
 					(reg_q133 AND symb_decoder(16#81#)) OR
 					(reg_q133 AND symb_decoder(16#86#)) OR
 					(reg_q133 AND symb_decoder(16#18#)) OR
 					(reg_q133 AND symb_decoder(16#b5#)) OR
 					(reg_q133 AND symb_decoder(16#1b#)) OR
 					(reg_q133 AND symb_decoder(16#63#)) OR
 					(reg_q133 AND symb_decoder(16#b4#)) OR
 					(reg_q133 AND symb_decoder(16#62#)) OR
 					(reg_q133 AND symb_decoder(16#8d#)) OR
 					(reg_q133 AND symb_decoder(16#09#)) OR
 					(reg_q133 AND symb_decoder(16#c8#)) OR
 					(reg_q133 AND symb_decoder(16#5c#)) OR
 					(reg_q133 AND symb_decoder(16#c4#)) OR
 					(reg_q133 AND symb_decoder(16#75#)) OR
 					(reg_q133 AND symb_decoder(16#b1#)) OR
 					(reg_q133 AND symb_decoder(16#ad#)) OR
 					(reg_q133 AND symb_decoder(16#d0#)) OR
 					(reg_q133 AND symb_decoder(16#c5#)) OR
 					(reg_q133 AND symb_decoder(16#05#)) OR
 					(reg_q133 AND symb_decoder(16#f0#)) OR
 					(reg_q133 AND symb_decoder(16#ae#)) OR
 					(reg_q133 AND symb_decoder(16#a8#)) OR
 					(reg_q133 AND symb_decoder(16#c0#)) OR
 					(reg_q133 AND symb_decoder(16#08#)) OR
 					(reg_q133 AND symb_decoder(16#78#)) OR
 					(reg_q133 AND symb_decoder(16#0d#)) OR
 					(reg_q133 AND symb_decoder(16#85#)) OR
 					(reg_q133 AND symb_decoder(16#15#)) OR
 					(reg_q133 AND symb_decoder(16#2c#)) OR
 					(reg_q133 AND symb_decoder(16#64#)) OR
 					(reg_q133 AND symb_decoder(16#8f#)) OR
 					(reg_q133 AND symb_decoder(16#cd#)) OR
 					(reg_q133 AND symb_decoder(16#e7#)) OR
 					(reg_q133 AND symb_decoder(16#c1#)) OR
 					(reg_q133 AND symb_decoder(16#e8#)) OR
 					(reg_q133 AND symb_decoder(16#5d#)) OR
 					(reg_q133 AND symb_decoder(16#4d#)) OR
 					(reg_q133 AND symb_decoder(16#35#)) OR
 					(reg_q133 AND symb_decoder(16#51#)) OR
 					(reg_q133 AND symb_decoder(16#ac#)) OR
 					(reg_q133 AND symb_decoder(16#f9#)) OR
 					(reg_q133 AND symb_decoder(16#1e#)) OR
 					(reg_q133 AND symb_decoder(16#db#)) OR
 					(reg_q133 AND symb_decoder(16#52#)) OR
 					(reg_q133 AND symb_decoder(16#ba#)) OR
 					(reg_q133 AND symb_decoder(16#6b#)) OR
 					(reg_q133 AND symb_decoder(16#32#)) OR
 					(reg_q133 AND symb_decoder(16#e3#)) OR
 					(reg_q133 AND symb_decoder(16#89#)) OR
 					(reg_q133 AND symb_decoder(16#83#)) OR
 					(reg_q133 AND symb_decoder(16#53#)) OR
 					(reg_q133 AND symb_decoder(16#3a#)) OR
 					(reg_q133 AND symb_decoder(16#fd#)) OR
 					(reg_q133 AND symb_decoder(16#37#)) OR
 					(reg_q133 AND symb_decoder(16#61#)) OR
 					(reg_q133 AND symb_decoder(16#bc#)) OR
 					(reg_q133 AND symb_decoder(16#fa#)) OR
 					(reg_q133 AND symb_decoder(16#2b#)) OR
 					(reg_q133 AND symb_decoder(16#70#)) OR
 					(reg_q133 AND symb_decoder(16#54#)) OR
 					(reg_q133 AND symb_decoder(16#b2#)) OR
 					(reg_q133 AND symb_decoder(16#07#)) OR
 					(reg_q133 AND symb_decoder(16#da#)) OR
 					(reg_q133 AND symb_decoder(16#1c#)) OR
 					(reg_q133 AND symb_decoder(16#a3#)) OR
 					(reg_q133 AND symb_decoder(16#0b#)) OR
 					(reg_q133 AND symb_decoder(16#b0#)) OR
 					(reg_q133 AND symb_decoder(16#5e#)) OR
 					(reg_q133 AND symb_decoder(16#34#)) OR
 					(reg_q133 AND symb_decoder(16#45#)) OR
 					(reg_q133 AND symb_decoder(16#80#)) OR
 					(reg_q133 AND symb_decoder(16#47#)) OR
 					(reg_q133 AND symb_decoder(16#74#)) OR
 					(reg_q133 AND symb_decoder(16#0a#)) OR
 					(reg_q133 AND symb_decoder(16#24#)) OR
 					(reg_q133 AND symb_decoder(16#de#)) OR
 					(reg_q133 AND symb_decoder(16#66#)) OR
 					(reg_q133 AND symb_decoder(16#21#)) OR
 					(reg_q133 AND symb_decoder(16#c6#)) OR
 					(reg_q133 AND symb_decoder(16#f3#)) OR
 					(reg_q133 AND symb_decoder(16#50#)) OR
 					(reg_q133 AND symb_decoder(16#9d#)) OR
 					(reg_q133 AND symb_decoder(16#7f#)) OR
 					(reg_q133 AND symb_decoder(16#ee#)) OR
 					(reg_q133 AND symb_decoder(16#7e#)) OR
 					(reg_q133 AND symb_decoder(16#16#)) OR
 					(reg_q133 AND symb_decoder(16#87#)) OR
 					(reg_q133 AND symb_decoder(16#cf#)) OR
 					(reg_q133 AND symb_decoder(16#d6#)) OR
 					(reg_q133 AND symb_decoder(16#a0#)) OR
 					(reg_q133 AND symb_decoder(16#49#)) OR
 					(reg_q133 AND symb_decoder(16#6d#)) OR
 					(reg_q133 AND symb_decoder(16#20#)) OR
 					(reg_q133 AND symb_decoder(16#d5#)) OR
 					(reg_q133 AND symb_decoder(16#73#)) OR
 					(reg_q133 AND symb_decoder(16#91#)) OR
 					(reg_q133 AND symb_decoder(16#c3#)) OR
 					(reg_q133 AND symb_decoder(16#42#)) OR
 					(reg_q133 AND symb_decoder(16#9f#)) OR
 					(reg_q133 AND symb_decoder(16#7a#)) OR
 					(reg_q133 AND symb_decoder(16#1f#)) OR
 					(reg_q133 AND symb_decoder(16#01#)) OR
 					(reg_q133 AND symb_decoder(16#5b#)) OR
 					(reg_q133 AND symb_decoder(16#dd#)) OR
 					(reg_q133 AND symb_decoder(16#55#)) OR
 					(reg_q133 AND symb_decoder(16#3e#)) OR
 					(reg_q133 AND symb_decoder(16#a5#)) OR
 					(reg_q133 AND symb_decoder(16#2a#)) OR
 					(reg_q133 AND symb_decoder(16#ea#)) OR
 					(reg_q133 AND symb_decoder(16#7d#)) OR
 					(reg_q133 AND symb_decoder(16#3f#)) OR
 					(reg_q133 AND symb_decoder(16#8b#)) OR
 					(reg_q133 AND symb_decoder(16#f8#)) OR
 					(reg_q133 AND symb_decoder(16#68#)) OR
 					(reg_q133 AND symb_decoder(16#41#)) OR
 					(reg_q133 AND symb_decoder(16#71#)) OR
 					(reg_q133 AND symb_decoder(16#23#)) OR
 					(reg_q133 AND symb_decoder(16#82#)) OR
 					(reg_q133 AND symb_decoder(16#36#)) OR
 					(reg_q133 AND symb_decoder(16#aa#)) OR
 					(reg_q133 AND symb_decoder(16#3d#)) OR
 					(reg_q133 AND symb_decoder(16#27#)) OR
 					(reg_q133 AND symb_decoder(16#a7#)) OR
 					(reg_q133 AND symb_decoder(16#90#)) OR
 					(reg_q133 AND symb_decoder(16#9b#)) OR
 					(reg_q133 AND symb_decoder(16#a9#)) OR
 					(reg_q133 AND symb_decoder(16#06#)) OR
 					(reg_q133 AND symb_decoder(16#0f#)) OR
 					(reg_q133 AND symb_decoder(16#5a#)) OR
 					(reg_q133 AND symb_decoder(16#ce#)) OR
 					(reg_q133 AND symb_decoder(16#03#)) OR
 					(reg_q133 AND symb_decoder(16#26#)) OR
 					(reg_q133 AND symb_decoder(16#00#)) OR
 					(reg_q133 AND symb_decoder(16#d9#)) OR
 					(reg_q133 AND symb_decoder(16#fe#)) OR
 					(reg_q133 AND symb_decoder(16#a6#)) OR
 					(reg_q133 AND symb_decoder(16#b9#)) OR
 					(reg_q133 AND symb_decoder(16#d8#)) OR
 					(reg_q133 AND symb_decoder(16#79#)) OR
 					(reg_q133 AND symb_decoder(16#48#)) OR
 					(reg_q133 AND symb_decoder(16#8c#)) OR
 					(reg_q133 AND symb_decoder(16#be#)) OR
 					(reg_q133 AND symb_decoder(16#f4#)) OR
 					(reg_q133 AND symb_decoder(16#88#)) OR
 					(reg_q133 AND symb_decoder(16#d3#)) OR
 					(reg_q133 AND symb_decoder(16#92#)) OR
 					(reg_q133 AND symb_decoder(16#4c#)) OR
 					(reg_q133 AND symb_decoder(16#c7#)) OR
 					(reg_q133 AND symb_decoder(16#94#)) OR
 					(reg_q133 AND symb_decoder(16#6c#)) OR
 					(reg_q133 AND symb_decoder(16#7b#)) OR
 					(reg_q133 AND symb_decoder(16#ef#)) OR
 					(reg_q133 AND symb_decoder(16#ff#)) OR
 					(reg_q133 AND symb_decoder(16#60#)) OR
 					(reg_q133 AND symb_decoder(16#28#)) OR
 					(reg_q133 AND symb_decoder(16#44#)) OR
 					(reg_q133 AND symb_decoder(16#f5#)) OR
 					(reg_q133 AND symb_decoder(16#cb#)) OR
 					(reg_q133 AND symb_decoder(16#5f#)) OR
 					(reg_q133 AND symb_decoder(16#38#)) OR
 					(reg_q133 AND symb_decoder(16#af#)) OR
 					(reg_q133 AND symb_decoder(16#72#)) OR
 					(reg_q133 AND symb_decoder(16#77#)) OR
 					(reg_q133 AND symb_decoder(16#bd#)) OR
 					(reg_q133 AND symb_decoder(16#17#)) OR
 					(reg_q133 AND symb_decoder(16#4f#)) OR
 					(reg_q133 AND symb_decoder(16#e2#)) OR
 					(reg_q133 AND symb_decoder(16#2e#)) OR
 					(reg_q133 AND symb_decoder(16#9c#)) OR
 					(reg_q133 AND symb_decoder(16#fb#)) OR
 					(reg_q133 AND symb_decoder(16#40#)) OR
 					(reg_q133 AND symb_decoder(16#13#)) OR
 					(reg_q133 AND symb_decoder(16#3c#)) OR
 					(reg_q133 AND symb_decoder(16#57#)) OR
 					(reg_q133 AND symb_decoder(16#4a#)) OR
 					(reg_q133 AND symb_decoder(16#a2#)) OR
 					(reg_q133 AND symb_decoder(16#98#)) OR
 					(reg_q133 AND symb_decoder(16#4b#)) OR
 					(reg_q133 AND symb_decoder(16#a4#)) OR
 					(reg_q133 AND symb_decoder(16#93#)) OR
 					(reg_q133 AND symb_decoder(16#04#)) OR
 					(reg_q133 AND symb_decoder(16#58#)) OR
 					(reg_q133 AND symb_decoder(16#2d#)) OR
 					(reg_q133 AND symb_decoder(16#1a#)) OR
 					(reg_q133 AND symb_decoder(16#dc#)) OR
 					(reg_q133 AND symb_decoder(16#33#)) OR
 					(reg_q133 AND symb_decoder(16#f2#)) OR
 					(reg_q133 AND symb_decoder(16#69#)) OR
 					(reg_q133 AND symb_decoder(16#b6#)) OR
 					(reg_q133 AND symb_decoder(16#30#)) OR
 					(reg_q133 AND symb_decoder(16#56#)) OR
 					(reg_q133 AND symb_decoder(16#e6#)) OR
 					(reg_q133 AND symb_decoder(16#ab#)) OR
 					(reg_q133 AND symb_decoder(16#6a#)) OR
 					(reg_q133 AND symb_decoder(16#43#)) OR
 					(reg_q133 AND symb_decoder(16#e1#)) OR
 					(reg_q133 AND symb_decoder(16#b8#)) OR
 					(reg_q133 AND symb_decoder(16#e4#)) OR
 					(reg_q133 AND symb_decoder(16#e0#)) OR
 					(reg_q133 AND symb_decoder(16#76#)) OR
 					(reg_q133 AND symb_decoder(16#a1#)) OR
 					(reg_q133 AND symb_decoder(16#d1#)) OR
 					(reg_q133 AND symb_decoder(16#6f#)) OR
 					(reg_q133 AND symb_decoder(16#31#)) OR
 					(reg_q133 AND symb_decoder(16#fc#)) OR
 					(reg_q133 AND symb_decoder(16#46#)) OR
 					(reg_q133 AND symb_decoder(16#d4#)) OR
 					(reg_q133 AND symb_decoder(16#3b#)) OR
 					(reg_q133 AND symb_decoder(16#8a#)) OR
 					(reg_q133 AND symb_decoder(16#2f#)) OR
 					(reg_q133 AND symb_decoder(16#95#)) OR
 					(reg_q133 AND symb_decoder(16#97#)) OR
 					(reg_q133 AND symb_decoder(16#59#)) OR
 					(reg_q133 AND symb_decoder(16#c9#)) OR
 					(reg_q133 AND symb_decoder(16#b3#)) OR
 					(reg_q133 AND symb_decoder(16#f7#)) OR
 					(reg_q133 AND symb_decoder(16#19#)) OR
 					(reg_q133 AND symb_decoder(16#9e#)) OR
 					(reg_q133 AND symb_decoder(16#ed#)) OR
 					(reg_q133 AND symb_decoder(16#7c#)) OR
 					(reg_q133 AND symb_decoder(16#d7#)) OR
 					(reg_q133 AND symb_decoder(16#e5#)) OR
 					(reg_q133 AND symb_decoder(16#e9#)) OR
 					(reg_q133 AND symb_decoder(16#f1#)) OR
 					(reg_q133 AND symb_decoder(16#6e#)) OR
 					(reg_q133 AND symb_decoder(16#0c#)) OR
 					(reg_q133 AND symb_decoder(16#df#)) OR
 					(reg_q133 AND symb_decoder(16#12#)) OR
 					(reg_q133 AND symb_decoder(16#ec#)) OR
 					(reg_q133 AND symb_decoder(16#29#)) OR
 					(reg_q133 AND symb_decoder(16#10#)) OR
 					(reg_q133 AND symb_decoder(16#9a#)) OR
 					(reg_q133 AND symb_decoder(16#cc#)) OR
 					(reg_q133 AND symb_decoder(16#d2#)) OR
 					(reg_q133 AND symb_decoder(16#02#)) OR
 					(reg_q133 AND symb_decoder(16#1d#)) OR
 					(reg_q133 AND symb_decoder(16#65#)) OR
 					(reg_q133 AND symb_decoder(16#bf#)) OR
 					(reg_q133 AND symb_decoder(16#99#)) OR
 					(reg_q133 AND symb_decoder(16#14#)) OR
 					(reg_q133 AND symb_decoder(16#67#)) OR
 					(reg_q133 AND symb_decoder(16#84#)) OR
 					(reg_q133 AND symb_decoder(16#eb#)) OR
 					(reg_q133 AND symb_decoder(16#8e#)) OR
 					(reg_q133 AND symb_decoder(16#39#));
reg_q133_init <= '0' ;
	p_reg_q133: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q133 <= reg_q133_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q133 <= reg_q133_init;
        else
          reg_q133 <= reg_q133_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1204_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1204 AND symb_decoder(16#33#)) OR
 					(reg_q1204 AND symb_decoder(16#f9#)) OR
 					(reg_q1204 AND symb_decoder(16#1f#)) OR
 					(reg_q1204 AND symb_decoder(16#d3#)) OR
 					(reg_q1204 AND symb_decoder(16#7a#)) OR
 					(reg_q1204 AND symb_decoder(16#bf#)) OR
 					(reg_q1204 AND symb_decoder(16#80#)) OR
 					(reg_q1204 AND symb_decoder(16#b1#)) OR
 					(reg_q1204 AND symb_decoder(16#f7#)) OR
 					(reg_q1204 AND symb_decoder(16#b7#)) OR
 					(reg_q1204 AND symb_decoder(16#a3#)) OR
 					(reg_q1204 AND symb_decoder(16#d1#)) OR
 					(reg_q1204 AND symb_decoder(16#8c#)) OR
 					(reg_q1204 AND symb_decoder(16#24#)) OR
 					(reg_q1204 AND symb_decoder(16#0e#)) OR
 					(reg_q1204 AND symb_decoder(16#b8#)) OR
 					(reg_q1204 AND symb_decoder(16#0a#)) OR
 					(reg_q1204 AND symb_decoder(16#6b#)) OR
 					(reg_q1204 AND symb_decoder(16#ee#)) OR
 					(reg_q1204 AND symb_decoder(16#2e#)) OR
 					(reg_q1204 AND symb_decoder(16#da#)) OR
 					(reg_q1204 AND symb_decoder(16#db#)) OR
 					(reg_q1204 AND symb_decoder(16#b4#)) OR
 					(reg_q1204 AND symb_decoder(16#50#)) OR
 					(reg_q1204 AND symb_decoder(16#97#)) OR
 					(reg_q1204 AND symb_decoder(16#89#)) OR
 					(reg_q1204 AND symb_decoder(16#aa#)) OR
 					(reg_q1204 AND symb_decoder(16#a0#)) OR
 					(reg_q1204 AND symb_decoder(16#12#)) OR
 					(reg_q1204 AND symb_decoder(16#63#)) OR
 					(reg_q1204 AND symb_decoder(16#9d#)) OR
 					(reg_q1204 AND symb_decoder(16#e0#)) OR
 					(reg_q1204 AND symb_decoder(16#ac#)) OR
 					(reg_q1204 AND symb_decoder(16#6c#)) OR
 					(reg_q1204 AND symb_decoder(16#e7#)) OR
 					(reg_q1204 AND symb_decoder(16#20#)) OR
 					(reg_q1204 AND symb_decoder(16#b2#)) OR
 					(reg_q1204 AND symb_decoder(16#3a#)) OR
 					(reg_q1204 AND symb_decoder(16#cf#)) OR
 					(reg_q1204 AND symb_decoder(16#66#)) OR
 					(reg_q1204 AND symb_decoder(16#cc#)) OR
 					(reg_q1204 AND symb_decoder(16#22#)) OR
 					(reg_q1204 AND symb_decoder(16#37#)) OR
 					(reg_q1204 AND symb_decoder(16#ef#)) OR
 					(reg_q1204 AND symb_decoder(16#32#)) OR
 					(reg_q1204 AND symb_decoder(16#46#)) OR
 					(reg_q1204 AND symb_decoder(16#76#)) OR
 					(reg_q1204 AND symb_decoder(16#a4#)) OR
 					(reg_q1204 AND symb_decoder(16#a7#)) OR
 					(reg_q1204 AND symb_decoder(16#93#)) OR
 					(reg_q1204 AND symb_decoder(16#df#)) OR
 					(reg_q1204 AND symb_decoder(16#c3#)) OR
 					(reg_q1204 AND symb_decoder(16#7b#)) OR
 					(reg_q1204 AND symb_decoder(16#6d#)) OR
 					(reg_q1204 AND symb_decoder(16#7c#)) OR
 					(reg_q1204 AND symb_decoder(16#ff#)) OR
 					(reg_q1204 AND symb_decoder(16#f2#)) OR
 					(reg_q1204 AND symb_decoder(16#42#)) OR
 					(reg_q1204 AND symb_decoder(16#57#)) OR
 					(reg_q1204 AND symb_decoder(16#60#)) OR
 					(reg_q1204 AND symb_decoder(16#9a#)) OR
 					(reg_q1204 AND symb_decoder(16#6f#)) OR
 					(reg_q1204 AND symb_decoder(16#ce#)) OR
 					(reg_q1204 AND symb_decoder(16#c2#)) OR
 					(reg_q1204 AND symb_decoder(16#61#)) OR
 					(reg_q1204 AND symb_decoder(16#0c#)) OR
 					(reg_q1204 AND symb_decoder(16#26#)) OR
 					(reg_q1204 AND symb_decoder(16#45#)) OR
 					(reg_q1204 AND symb_decoder(16#5f#)) OR
 					(reg_q1204 AND symb_decoder(16#28#)) OR
 					(reg_q1204 AND symb_decoder(16#51#)) OR
 					(reg_q1204 AND symb_decoder(16#73#)) OR
 					(reg_q1204 AND symb_decoder(16#75#)) OR
 					(reg_q1204 AND symb_decoder(16#d8#)) OR
 					(reg_q1204 AND symb_decoder(16#43#)) OR
 					(reg_q1204 AND symb_decoder(16#a8#)) OR
 					(reg_q1204 AND symb_decoder(16#8b#)) OR
 					(reg_q1204 AND symb_decoder(16#af#)) OR
 					(reg_q1204 AND symb_decoder(16#71#)) OR
 					(reg_q1204 AND symb_decoder(16#9e#)) OR
 					(reg_q1204 AND symb_decoder(16#16#)) OR
 					(reg_q1204 AND symb_decoder(16#ad#)) OR
 					(reg_q1204 AND symb_decoder(16#ea#)) OR
 					(reg_q1204 AND symb_decoder(16#dc#)) OR
 					(reg_q1204 AND symb_decoder(16#07#)) OR
 					(reg_q1204 AND symb_decoder(16#87#)) OR
 					(reg_q1204 AND symb_decoder(16#d0#)) OR
 					(reg_q1204 AND symb_decoder(16#15#)) OR
 					(reg_q1204 AND symb_decoder(16#a6#)) OR
 					(reg_q1204 AND symb_decoder(16#74#)) OR
 					(reg_q1204 AND symb_decoder(16#38#)) OR
 					(reg_q1204 AND symb_decoder(16#0d#)) OR
 					(reg_q1204 AND symb_decoder(16#94#)) OR
 					(reg_q1204 AND symb_decoder(16#5a#)) OR
 					(reg_q1204 AND symb_decoder(16#91#)) OR
 					(reg_q1204 AND symb_decoder(16#dd#)) OR
 					(reg_q1204 AND symb_decoder(16#cd#)) OR
 					(reg_q1204 AND symb_decoder(16#be#)) OR
 					(reg_q1204 AND symb_decoder(16#36#)) OR
 					(reg_q1204 AND symb_decoder(16#72#)) OR
 					(reg_q1204 AND symb_decoder(16#1d#)) OR
 					(reg_q1204 AND symb_decoder(16#c6#)) OR
 					(reg_q1204 AND symb_decoder(16#5d#)) OR
 					(reg_q1204 AND symb_decoder(16#4f#)) OR
 					(reg_q1204 AND symb_decoder(16#a2#)) OR
 					(reg_q1204 AND symb_decoder(16#f5#)) OR
 					(reg_q1204 AND symb_decoder(16#8f#)) OR
 					(reg_q1204 AND symb_decoder(16#cb#)) OR
 					(reg_q1204 AND symb_decoder(16#39#)) OR
 					(reg_q1204 AND symb_decoder(16#98#)) OR
 					(reg_q1204 AND symb_decoder(16#2a#)) OR
 					(reg_q1204 AND symb_decoder(16#e8#)) OR
 					(reg_q1204 AND symb_decoder(16#0b#)) OR
 					(reg_q1204 AND symb_decoder(16#f4#)) OR
 					(reg_q1204 AND symb_decoder(16#4c#)) OR
 					(reg_q1204 AND symb_decoder(16#ae#)) OR
 					(reg_q1204 AND symb_decoder(16#19#)) OR
 					(reg_q1204 AND symb_decoder(16#1c#)) OR
 					(reg_q1204 AND symb_decoder(16#f1#)) OR
 					(reg_q1204 AND symb_decoder(16#e5#)) OR
 					(reg_q1204 AND symb_decoder(16#54#)) OR
 					(reg_q1204 AND symb_decoder(16#f6#)) OR
 					(reg_q1204 AND symb_decoder(16#d7#)) OR
 					(reg_q1204 AND symb_decoder(16#17#)) OR
 					(reg_q1204 AND symb_decoder(16#95#)) OR
 					(reg_q1204 AND symb_decoder(16#64#)) OR
 					(reg_q1204 AND symb_decoder(16#96#)) OR
 					(reg_q1204 AND symb_decoder(16#53#)) OR
 					(reg_q1204 AND symb_decoder(16#d2#)) OR
 					(reg_q1204 AND symb_decoder(16#e6#)) OR
 					(reg_q1204 AND symb_decoder(16#55#)) OR
 					(reg_q1204 AND symb_decoder(16#b5#)) OR
 					(reg_q1204 AND symb_decoder(16#2b#)) OR
 					(reg_q1204 AND symb_decoder(16#fb#)) OR
 					(reg_q1204 AND symb_decoder(16#79#)) OR
 					(reg_q1204 AND symb_decoder(16#f3#)) OR
 					(reg_q1204 AND symb_decoder(16#fe#)) OR
 					(reg_q1204 AND symb_decoder(16#d4#)) OR
 					(reg_q1204 AND symb_decoder(16#4b#)) OR
 					(reg_q1204 AND symb_decoder(16#62#)) OR
 					(reg_q1204 AND symb_decoder(16#09#)) OR
 					(reg_q1204 AND symb_decoder(16#7e#)) OR
 					(reg_q1204 AND symb_decoder(16#27#)) OR
 					(reg_q1204 AND symb_decoder(16#18#)) OR
 					(reg_q1204 AND symb_decoder(16#21#)) OR
 					(reg_q1204 AND symb_decoder(16#c1#)) OR
 					(reg_q1204 AND symb_decoder(16#fd#)) OR
 					(reg_q1204 AND symb_decoder(16#59#)) OR
 					(reg_q1204 AND symb_decoder(16#e2#)) OR
 					(reg_q1204 AND symb_decoder(16#b9#)) OR
 					(reg_q1204 AND symb_decoder(16#29#)) OR
 					(reg_q1204 AND symb_decoder(16#8a#)) OR
 					(reg_q1204 AND symb_decoder(16#3b#)) OR
 					(reg_q1204 AND symb_decoder(16#30#)) OR
 					(reg_q1204 AND symb_decoder(16#3e#)) OR
 					(reg_q1204 AND symb_decoder(16#02#)) OR
 					(reg_q1204 AND symb_decoder(16#86#)) OR
 					(reg_q1204 AND symb_decoder(16#eb#)) OR
 					(reg_q1204 AND symb_decoder(16#e4#)) OR
 					(reg_q1204 AND symb_decoder(16#11#)) OR
 					(reg_q1204 AND symb_decoder(16#bd#)) OR
 					(reg_q1204 AND symb_decoder(16#a9#)) OR
 					(reg_q1204 AND symb_decoder(16#06#)) OR
 					(reg_q1204 AND symb_decoder(16#99#)) OR
 					(reg_q1204 AND symb_decoder(16#e9#)) OR
 					(reg_q1204 AND symb_decoder(16#c4#)) OR
 					(reg_q1204 AND symb_decoder(16#1e#)) OR
 					(reg_q1204 AND symb_decoder(16#3f#)) OR
 					(reg_q1204 AND symb_decoder(16#5b#)) OR
 					(reg_q1204 AND symb_decoder(16#49#)) OR
 					(reg_q1204 AND symb_decoder(16#fa#)) OR
 					(reg_q1204 AND symb_decoder(16#9b#)) OR
 					(reg_q1204 AND symb_decoder(16#d9#)) OR
 					(reg_q1204 AND symb_decoder(16#bc#)) OR
 					(reg_q1204 AND symb_decoder(16#e3#)) OR
 					(reg_q1204 AND symb_decoder(16#4a#)) OR
 					(reg_q1204 AND symb_decoder(16#10#)) OR
 					(reg_q1204 AND symb_decoder(16#84#)) OR
 					(reg_q1204 AND symb_decoder(16#d5#)) OR
 					(reg_q1204 AND symb_decoder(16#68#)) OR
 					(reg_q1204 AND symb_decoder(16#6e#)) OR
 					(reg_q1204 AND symb_decoder(16#de#)) OR
 					(reg_q1204 AND symb_decoder(16#78#)) OR
 					(reg_q1204 AND symb_decoder(16#13#)) OR
 					(reg_q1204 AND symb_decoder(16#8e#)) OR
 					(reg_q1204 AND symb_decoder(16#47#)) OR
 					(reg_q1204 AND symb_decoder(16#3d#)) OR
 					(reg_q1204 AND symb_decoder(16#f0#)) OR
 					(reg_q1204 AND symb_decoder(16#88#)) OR
 					(reg_q1204 AND symb_decoder(16#c8#)) OR
 					(reg_q1204 AND symb_decoder(16#b3#)) OR
 					(reg_q1204 AND symb_decoder(16#05#)) OR
 					(reg_q1204 AND symb_decoder(16#2f#)) OR
 					(reg_q1204 AND symb_decoder(16#e1#)) OR
 					(reg_q1204 AND symb_decoder(16#ca#)) OR
 					(reg_q1204 AND symb_decoder(16#2c#)) OR
 					(reg_q1204 AND symb_decoder(16#81#)) OR
 					(reg_q1204 AND symb_decoder(16#4e#)) OR
 					(reg_q1204 AND symb_decoder(16#25#)) OR
 					(reg_q1204 AND symb_decoder(16#77#)) OR
 					(reg_q1204 AND symb_decoder(16#8d#)) OR
 					(reg_q1204 AND symb_decoder(16#0f#)) OR
 					(reg_q1204 AND symb_decoder(16#14#)) OR
 					(reg_q1204 AND symb_decoder(16#40#)) OR
 					(reg_q1204 AND symb_decoder(16#58#)) OR
 					(reg_q1204 AND symb_decoder(16#c0#)) OR
 					(reg_q1204 AND symb_decoder(16#23#)) OR
 					(reg_q1204 AND symb_decoder(16#35#)) OR
 					(reg_q1204 AND symb_decoder(16#4d#)) OR
 					(reg_q1204 AND symb_decoder(16#bb#)) OR
 					(reg_q1204 AND symb_decoder(16#5e#)) OR
 					(reg_q1204 AND symb_decoder(16#08#)) OR
 					(reg_q1204 AND symb_decoder(16#03#)) OR
 					(reg_q1204 AND symb_decoder(16#a1#)) OR
 					(reg_q1204 AND symb_decoder(16#c7#)) OR
 					(reg_q1204 AND symb_decoder(16#85#)) OR
 					(reg_q1204 AND symb_decoder(16#c9#)) OR
 					(reg_q1204 AND symb_decoder(16#5c#)) OR
 					(reg_q1204 AND symb_decoder(16#a5#)) OR
 					(reg_q1204 AND symb_decoder(16#ab#)) OR
 					(reg_q1204 AND symb_decoder(16#ba#)) OR
 					(reg_q1204 AND symb_decoder(16#1a#)) OR
 					(reg_q1204 AND symb_decoder(16#48#)) OR
 					(reg_q1204 AND symb_decoder(16#65#)) OR
 					(reg_q1204 AND symb_decoder(16#56#)) OR
 					(reg_q1204 AND symb_decoder(16#ed#)) OR
 					(reg_q1204 AND symb_decoder(16#c5#)) OR
 					(reg_q1204 AND symb_decoder(16#69#)) OR
 					(reg_q1204 AND symb_decoder(16#67#)) OR
 					(reg_q1204 AND symb_decoder(16#9f#)) OR
 					(reg_q1204 AND symb_decoder(16#7d#)) OR
 					(reg_q1204 AND symb_decoder(16#9c#)) OR
 					(reg_q1204 AND symb_decoder(16#04#)) OR
 					(reg_q1204 AND symb_decoder(16#83#)) OR
 					(reg_q1204 AND symb_decoder(16#3c#)) OR
 					(reg_q1204 AND symb_decoder(16#92#)) OR
 					(reg_q1204 AND symb_decoder(16#b0#)) OR
 					(reg_q1204 AND symb_decoder(16#7f#)) OR
 					(reg_q1204 AND symb_decoder(16#fc#)) OR
 					(reg_q1204 AND symb_decoder(16#6a#)) OR
 					(reg_q1204 AND symb_decoder(16#31#)) OR
 					(reg_q1204 AND symb_decoder(16#f8#)) OR
 					(reg_q1204 AND symb_decoder(16#70#)) OR
 					(reg_q1204 AND symb_decoder(16#44#)) OR
 					(reg_q1204 AND symb_decoder(16#00#)) OR
 					(reg_q1204 AND symb_decoder(16#90#)) OR
 					(reg_q1204 AND symb_decoder(16#b6#)) OR
 					(reg_q1204 AND symb_decoder(16#d6#)) OR
 					(reg_q1204 AND symb_decoder(16#82#)) OR
 					(reg_q1204 AND symb_decoder(16#ec#)) OR
 					(reg_q1204 AND symb_decoder(16#34#)) OR
 					(reg_q1204 AND symb_decoder(16#41#)) OR
 					(reg_q1204 AND symb_decoder(16#52#)) OR
 					(reg_q1204 AND symb_decoder(16#01#)) OR
 					(reg_q1204 AND symb_decoder(16#1b#)) OR
 					(reg_q1204 AND symb_decoder(16#2d#));
reg_q1204_init <= '0' ;
	p_reg_q1204: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1204 <= reg_q1204_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1204 <= reg_q1204_init;
        else
          reg_q1204 <= reg_q1204_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph38

reg_q2216_in <= (reg_q2216 AND symb_decoder(16#31#)) OR
 					(reg_q2216 AND symb_decoder(16#82#)) OR
 					(reg_q2216 AND symb_decoder(16#ae#)) OR
 					(reg_q2216 AND symb_decoder(16#ca#)) OR
 					(reg_q2216 AND symb_decoder(16#87#)) OR
 					(reg_q2216 AND symb_decoder(16#8c#)) OR
 					(reg_q2216 AND symb_decoder(16#be#)) OR
 					(reg_q2216 AND symb_decoder(16#6c#)) OR
 					(reg_q2216 AND symb_decoder(16#9e#)) OR
 					(reg_q2216 AND symb_decoder(16#90#)) OR
 					(reg_q2216 AND symb_decoder(16#f3#)) OR
 					(reg_q2216 AND symb_decoder(16#41#)) OR
 					(reg_q2216 AND symb_decoder(16#d7#)) OR
 					(reg_q2216 AND symb_decoder(16#b1#)) OR
 					(reg_q2216 AND symb_decoder(16#77#)) OR
 					(reg_q2216 AND symb_decoder(16#de#)) OR
 					(reg_q2216 AND symb_decoder(16#18#)) OR
 					(reg_q2216 AND symb_decoder(16#56#)) OR
 					(reg_q2216 AND symb_decoder(16#36#)) OR
 					(reg_q2216 AND symb_decoder(16#cd#)) OR
 					(reg_q2216 AND symb_decoder(16#ff#)) OR
 					(reg_q2216 AND symb_decoder(16#da#)) OR
 					(reg_q2216 AND symb_decoder(16#54#)) OR
 					(reg_q2216 AND symb_decoder(16#38#)) OR
 					(reg_q2216 AND symb_decoder(16#3b#)) OR
 					(reg_q2216 AND symb_decoder(16#07#)) OR
 					(reg_q2216 AND symb_decoder(16#a7#)) OR
 					(reg_q2216 AND symb_decoder(16#2f#)) OR
 					(reg_q2216 AND symb_decoder(16#bf#)) OR
 					(reg_q2216 AND symb_decoder(16#9b#)) OR
 					(reg_q2216 AND symb_decoder(16#63#)) OR
 					(reg_q2216 AND symb_decoder(16#37#)) OR
 					(reg_q2216 AND symb_decoder(16#fb#)) OR
 					(reg_q2216 AND symb_decoder(16#cb#)) OR
 					(reg_q2216 AND symb_decoder(16#ef#)) OR
 					(reg_q2216 AND symb_decoder(16#58#)) OR
 					(reg_q2216 AND symb_decoder(16#a3#)) OR
 					(reg_q2216 AND symb_decoder(16#75#)) OR
 					(reg_q2216 AND symb_decoder(16#4e#)) OR
 					(reg_q2216 AND symb_decoder(16#f4#)) OR
 					(reg_q2216 AND symb_decoder(16#7a#)) OR
 					(reg_q2216 AND symb_decoder(16#93#)) OR
 					(reg_q2216 AND symb_decoder(16#4a#)) OR
 					(reg_q2216 AND symb_decoder(16#14#)) OR
 					(reg_q2216 AND symb_decoder(16#3c#)) OR
 					(reg_q2216 AND symb_decoder(16#ee#)) OR
 					(reg_q2216 AND symb_decoder(16#69#)) OR
 					(reg_q2216 AND symb_decoder(16#1d#)) OR
 					(reg_q2216 AND symb_decoder(16#83#)) OR
 					(reg_q2216 AND symb_decoder(16#76#)) OR
 					(reg_q2216 AND symb_decoder(16#00#)) OR
 					(reg_q2216 AND symb_decoder(16#c0#)) OR
 					(reg_q2216 AND symb_decoder(16#04#)) OR
 					(reg_q2216 AND symb_decoder(16#5a#)) OR
 					(reg_q2216 AND symb_decoder(16#65#)) OR
 					(reg_q2216 AND symb_decoder(16#4f#)) OR
 					(reg_q2216 AND symb_decoder(16#29#)) OR
 					(reg_q2216 AND symb_decoder(16#b3#)) OR
 					(reg_q2216 AND symb_decoder(16#13#)) OR
 					(reg_q2216 AND symb_decoder(16#7b#)) OR
 					(reg_q2216 AND symb_decoder(16#60#)) OR
 					(reg_q2216 AND symb_decoder(16#dd#)) OR
 					(reg_q2216 AND symb_decoder(16#ba#)) OR
 					(reg_q2216 AND symb_decoder(16#47#)) OR
 					(reg_q2216 AND symb_decoder(16#d4#)) OR
 					(reg_q2216 AND symb_decoder(16#23#)) OR
 					(reg_q2216 AND symb_decoder(16#4c#)) OR
 					(reg_q2216 AND symb_decoder(16#f9#)) OR
 					(reg_q2216 AND symb_decoder(16#a6#)) OR
 					(reg_q2216 AND symb_decoder(16#26#)) OR
 					(reg_q2216 AND symb_decoder(16#e8#)) OR
 					(reg_q2216 AND symb_decoder(16#7e#)) OR
 					(reg_q2216 AND symb_decoder(16#89#)) OR
 					(reg_q2216 AND symb_decoder(16#34#)) OR
 					(reg_q2216 AND symb_decoder(16#c3#)) OR
 					(reg_q2216 AND symb_decoder(16#c8#)) OR
 					(reg_q2216 AND symb_decoder(16#01#)) OR
 					(reg_q2216 AND symb_decoder(16#43#)) OR
 					(reg_q2216 AND symb_decoder(16#e4#)) OR
 					(reg_q2216 AND symb_decoder(16#9c#)) OR
 					(reg_q2216 AND symb_decoder(16#71#)) OR
 					(reg_q2216 AND symb_decoder(16#19#)) OR
 					(reg_q2216 AND symb_decoder(16#97#)) OR
 					(reg_q2216 AND symb_decoder(16#95#)) OR
 					(reg_q2216 AND symb_decoder(16#8b#)) OR
 					(reg_q2216 AND symb_decoder(16#d3#)) OR
 					(reg_q2216 AND symb_decoder(16#e2#)) OR
 					(reg_q2216 AND symb_decoder(16#9f#)) OR
 					(reg_q2216 AND symb_decoder(16#0b#)) OR
 					(reg_q2216 AND symb_decoder(16#80#)) OR
 					(reg_q2216 AND symb_decoder(16#3d#)) OR
 					(reg_q2216 AND symb_decoder(16#d9#)) OR
 					(reg_q2216 AND symb_decoder(16#c1#)) OR
 					(reg_q2216 AND symb_decoder(16#a4#)) OR
 					(reg_q2216 AND symb_decoder(16#84#)) OR
 					(reg_q2216 AND symb_decoder(16#0f#)) OR
 					(reg_q2216 AND symb_decoder(16#35#)) OR
 					(reg_q2216 AND symb_decoder(16#c2#)) OR
 					(reg_q2216 AND symb_decoder(16#e6#)) OR
 					(reg_q2216 AND symb_decoder(16#02#)) OR
 					(reg_q2216 AND symb_decoder(16#61#)) OR
 					(reg_q2216 AND symb_decoder(16#e3#)) OR
 					(reg_q2216 AND symb_decoder(16#ec#)) OR
 					(reg_q2216 AND symb_decoder(16#a5#)) OR
 					(reg_q2216 AND symb_decoder(16#10#)) OR
 					(reg_q2216 AND symb_decoder(16#eb#)) OR
 					(reg_q2216 AND symb_decoder(16#a2#)) OR
 					(reg_q2216 AND symb_decoder(16#f5#)) OR
 					(reg_q2216 AND symb_decoder(16#5e#)) OR
 					(reg_q2216 AND symb_decoder(16#c5#)) OR
 					(reg_q2216 AND symb_decoder(16#e9#)) OR
 					(reg_q2216 AND symb_decoder(16#67#)) OR
 					(reg_q2216 AND symb_decoder(16#4d#)) OR
 					(reg_q2216 AND symb_decoder(16#f2#)) OR
 					(reg_q2216 AND symb_decoder(16#2e#)) OR
 					(reg_q2216 AND symb_decoder(16#86#)) OR
 					(reg_q2216 AND symb_decoder(16#d6#)) OR
 					(reg_q2216 AND symb_decoder(16#44#)) OR
 					(reg_q2216 AND symb_decoder(16#d5#)) OR
 					(reg_q2216 AND symb_decoder(16#03#)) OR
 					(reg_q2216 AND symb_decoder(16#22#)) OR
 					(reg_q2216 AND symb_decoder(16#f7#)) OR
 					(reg_q2216 AND symb_decoder(16#59#)) OR
 					(reg_q2216 AND symb_decoder(16#f1#)) OR
 					(reg_q2216 AND symb_decoder(16#09#)) OR
 					(reg_q2216 AND symb_decoder(16#bc#)) OR
 					(reg_q2216 AND symb_decoder(16#52#)) OR
 					(reg_q2216 AND symb_decoder(16#0c#)) OR
 					(reg_q2216 AND symb_decoder(16#f0#)) OR
 					(reg_q2216 AND symb_decoder(16#d2#)) OR
 					(reg_q2216 AND symb_decoder(16#fd#)) OR
 					(reg_q2216 AND symb_decoder(16#8a#)) OR
 					(reg_q2216 AND symb_decoder(16#aa#)) OR
 					(reg_q2216 AND symb_decoder(16#df#)) OR
 					(reg_q2216 AND symb_decoder(16#06#)) OR
 					(reg_q2216 AND symb_decoder(16#0e#)) OR
 					(reg_q2216 AND symb_decoder(16#11#)) OR
 					(reg_q2216 AND symb_decoder(16#50#)) OR
 					(reg_q2216 AND symb_decoder(16#dc#)) OR
 					(reg_q2216 AND symb_decoder(16#99#)) OR
 					(reg_q2216 AND symb_decoder(16#f6#)) OR
 					(reg_q2216 AND symb_decoder(16#bb#)) OR
 					(reg_q2216 AND symb_decoder(16#a9#)) OR
 					(reg_q2216 AND symb_decoder(16#85#)) OR
 					(reg_q2216 AND symb_decoder(16#f8#)) OR
 					(reg_q2216 AND symb_decoder(16#98#)) OR
 					(reg_q2216 AND symb_decoder(16#af#)) OR
 					(reg_q2216 AND symb_decoder(16#ed#)) OR
 					(reg_q2216 AND symb_decoder(16#64#)) OR
 					(reg_q2216 AND symb_decoder(16#e1#)) OR
 					(reg_q2216 AND symb_decoder(16#ad#)) OR
 					(reg_q2216 AND symb_decoder(16#6e#)) OR
 					(reg_q2216 AND symb_decoder(16#46#)) OR
 					(reg_q2216 AND symb_decoder(16#7f#)) OR
 					(reg_q2216 AND symb_decoder(16#ce#)) OR
 					(reg_q2216 AND symb_decoder(16#12#)) OR
 					(reg_q2216 AND symb_decoder(16#b0#)) OR
 					(reg_q2216 AND symb_decoder(16#b5#)) OR
 					(reg_q2216 AND symb_decoder(16#fc#)) OR
 					(reg_q2216 AND symb_decoder(16#9d#)) OR
 					(reg_q2216 AND symb_decoder(16#25#)) OR
 					(reg_q2216 AND symb_decoder(16#d8#)) OR
 					(reg_q2216 AND symb_decoder(16#27#)) OR
 					(reg_q2216 AND symb_decoder(16#b4#)) OR
 					(reg_q2216 AND symb_decoder(16#b9#)) OR
 					(reg_q2216 AND symb_decoder(16#30#)) OR
 					(reg_q2216 AND symb_decoder(16#5d#)) OR
 					(reg_q2216 AND symb_decoder(16#55#)) OR
 					(reg_q2216 AND symb_decoder(16#e7#)) OR
 					(reg_q2216 AND symb_decoder(16#9a#)) OR
 					(reg_q2216 AND symb_decoder(16#a0#)) OR
 					(reg_q2216 AND symb_decoder(16#b8#)) OR
 					(reg_q2216 AND symb_decoder(16#cc#)) OR
 					(reg_q2216 AND symb_decoder(16#6f#)) OR
 					(reg_q2216 AND symb_decoder(16#66#)) OR
 					(reg_q2216 AND symb_decoder(16#3f#)) OR
 					(reg_q2216 AND symb_decoder(16#2b#)) OR
 					(reg_q2216 AND symb_decoder(16#51#)) OR
 					(reg_q2216 AND symb_decoder(16#49#)) OR
 					(reg_q2216 AND symb_decoder(16#6d#)) OR
 					(reg_q2216 AND symb_decoder(16#e5#)) OR
 					(reg_q2216 AND symb_decoder(16#fe#)) OR
 					(reg_q2216 AND symb_decoder(16#5b#)) OR
 					(reg_q2216 AND symb_decoder(16#c9#)) OR
 					(reg_q2216 AND symb_decoder(16#70#)) OR
 					(reg_q2216 AND symb_decoder(16#5c#)) OR
 					(reg_q2216 AND symb_decoder(16#08#)) OR
 					(reg_q2216 AND symb_decoder(16#7c#)) OR
 					(reg_q2216 AND symb_decoder(16#92#)) OR
 					(reg_q2216 AND symb_decoder(16#53#)) OR
 					(reg_q2216 AND symb_decoder(16#20#)) OR
 					(reg_q2216 AND symb_decoder(16#21#)) OR
 					(reg_q2216 AND symb_decoder(16#88#)) OR
 					(reg_q2216 AND symb_decoder(16#28#)) OR
 					(reg_q2216 AND symb_decoder(16#b6#)) OR
 					(reg_q2216 AND symb_decoder(16#ab#)) OR
 					(reg_q2216 AND symb_decoder(16#2d#)) OR
 					(reg_q2216 AND symb_decoder(16#4b#)) OR
 					(reg_q2216 AND symb_decoder(16#5f#)) OR
 					(reg_q2216 AND symb_decoder(16#1f#)) OR
 					(reg_q2216 AND symb_decoder(16#8d#)) OR
 					(reg_q2216 AND symb_decoder(16#b7#)) OR
 					(reg_q2216 AND symb_decoder(16#81#)) OR
 					(reg_q2216 AND symb_decoder(16#45#)) OR
 					(reg_q2216 AND symb_decoder(16#73#)) OR
 					(reg_q2216 AND symb_decoder(16#68#)) OR
 					(reg_q2216 AND symb_decoder(16#d1#)) OR
 					(reg_q2216 AND symb_decoder(16#96#)) OR
 					(reg_q2216 AND symb_decoder(16#6a#)) OR
 					(reg_q2216 AND symb_decoder(16#1c#)) OR
 					(reg_q2216 AND symb_decoder(16#ac#)) OR
 					(reg_q2216 AND symb_decoder(16#05#)) OR
 					(reg_q2216 AND symb_decoder(16#3a#)) OR
 					(reg_q2216 AND symb_decoder(16#7d#)) OR
 					(reg_q2216 AND symb_decoder(16#ea#)) OR
 					(reg_q2216 AND symb_decoder(16#c7#)) OR
 					(reg_q2216 AND symb_decoder(16#2c#)) OR
 					(reg_q2216 AND symb_decoder(16#8e#)) OR
 					(reg_q2216 AND symb_decoder(16#2a#)) OR
 					(reg_q2216 AND symb_decoder(16#e0#)) OR
 					(reg_q2216 AND symb_decoder(16#1e#)) OR
 					(reg_q2216 AND symb_decoder(16#fa#)) OR
 					(reg_q2216 AND symb_decoder(16#62#)) OR
 					(reg_q2216 AND symb_decoder(16#cf#)) OR
 					(reg_q2216 AND symb_decoder(16#33#)) OR
 					(reg_q2216 AND symb_decoder(16#3e#)) OR
 					(reg_q2216 AND symb_decoder(16#d0#)) OR
 					(reg_q2216 AND symb_decoder(16#17#)) OR
 					(reg_q2216 AND symb_decoder(16#c4#)) OR
 					(reg_q2216 AND symb_decoder(16#6b#)) OR
 					(reg_q2216 AND symb_decoder(16#a1#)) OR
 					(reg_q2216 AND symb_decoder(16#24#)) OR
 					(reg_q2216 AND symb_decoder(16#42#)) OR
 					(reg_q2216 AND symb_decoder(16#db#)) OR
 					(reg_q2216 AND symb_decoder(16#72#)) OR
 					(reg_q2216 AND symb_decoder(16#91#)) OR
 					(reg_q2216 AND symb_decoder(16#79#)) OR
 					(reg_q2216 AND symb_decoder(16#78#)) OR
 					(reg_q2216 AND symb_decoder(16#bd#)) OR
 					(reg_q2216 AND symb_decoder(16#1a#)) OR
 					(reg_q2216 AND symb_decoder(16#94#)) OR
 					(reg_q2216 AND symb_decoder(16#8f#)) OR
 					(reg_q2216 AND symb_decoder(16#48#)) OR
 					(reg_q2216 AND symb_decoder(16#57#)) OR
 					(reg_q2216 AND symb_decoder(16#16#)) OR
 					(reg_q2216 AND symb_decoder(16#40#)) OR
 					(reg_q2216 AND symb_decoder(16#1b#)) OR
 					(reg_q2216 AND symb_decoder(16#74#)) OR
 					(reg_q2216 AND symb_decoder(16#32#)) OR
 					(reg_q2216 AND symb_decoder(16#c6#)) OR
 					(reg_q2216 AND symb_decoder(16#b2#)) OR
 					(reg_q2216 AND symb_decoder(16#39#)) OR
 					(reg_q2216 AND symb_decoder(16#a8#)) OR
 					(reg_q2216 AND symb_decoder(16#15#)) OR
 					(reg_q2150 AND symb_decoder(16#13#)) OR
 					(reg_q2150 AND symb_decoder(16#6c#)) OR
 					(reg_q2150 AND symb_decoder(16#6e#)) OR
 					(reg_q2150 AND symb_decoder(16#f6#)) OR
 					(reg_q2150 AND symb_decoder(16#ad#)) OR
 					(reg_q2150 AND symb_decoder(16#5c#)) OR
 					(reg_q2150 AND symb_decoder(16#39#)) OR
 					(reg_q2150 AND symb_decoder(16#be#)) OR
 					(reg_q2150 AND symb_decoder(16#c3#)) OR
 					(reg_q2150 AND symb_decoder(16#27#)) OR
 					(reg_q2150 AND symb_decoder(16#3a#)) OR
 					(reg_q2150 AND symb_decoder(16#a7#)) OR
 					(reg_q2150 AND symb_decoder(16#b4#)) OR
 					(reg_q2150 AND symb_decoder(16#3f#)) OR
 					(reg_q2150 AND symb_decoder(16#f5#)) OR
 					(reg_q2150 AND symb_decoder(16#47#)) OR
 					(reg_q2150 AND symb_decoder(16#ab#)) OR
 					(reg_q2150 AND symb_decoder(16#a2#)) OR
 					(reg_q2150 AND symb_decoder(16#96#)) OR
 					(reg_q2150 AND symb_decoder(16#4f#)) OR
 					(reg_q2150 AND symb_decoder(16#1e#)) OR
 					(reg_q2150 AND symb_decoder(16#63#)) OR
 					(reg_q2150 AND symb_decoder(16#0b#)) OR
 					(reg_q2150 AND symb_decoder(16#60#)) OR
 					(reg_q2150 AND symb_decoder(16#fd#)) OR
 					(reg_q2150 AND symb_decoder(16#21#)) OR
 					(reg_q2150 AND symb_decoder(16#44#)) OR
 					(reg_q2150 AND symb_decoder(16#8a#)) OR
 					(reg_q2150 AND symb_decoder(16#ed#)) OR
 					(reg_q2150 AND symb_decoder(16#6f#)) OR
 					(reg_q2150 AND symb_decoder(16#4d#)) OR
 					(reg_q2150 AND symb_decoder(16#00#)) OR
 					(reg_q2150 AND symb_decoder(16#23#)) OR
 					(reg_q2150 AND symb_decoder(16#b3#)) OR
 					(reg_q2150 AND symb_decoder(16#7e#)) OR
 					(reg_q2150 AND symb_decoder(16#d8#)) OR
 					(reg_q2150 AND symb_decoder(16#48#)) OR
 					(reg_q2150 AND symb_decoder(16#7c#)) OR
 					(reg_q2150 AND symb_decoder(16#10#)) OR
 					(reg_q2150 AND symb_decoder(16#8d#)) OR
 					(reg_q2150 AND symb_decoder(16#d9#)) OR
 					(reg_q2150 AND symb_decoder(16#0e#)) OR
 					(reg_q2150 AND symb_decoder(16#49#)) OR
 					(reg_q2150 AND symb_decoder(16#a6#)) OR
 					(reg_q2150 AND symb_decoder(16#e6#)) OR
 					(reg_q2150 AND symb_decoder(16#bd#)) OR
 					(reg_q2150 AND symb_decoder(16#bb#)) OR
 					(reg_q2150 AND symb_decoder(16#62#)) OR
 					(reg_q2150 AND symb_decoder(16#c0#)) OR
 					(reg_q2150 AND symb_decoder(16#99#)) OR
 					(reg_q2150 AND symb_decoder(16#83#)) OR
 					(reg_q2150 AND symb_decoder(16#19#)) OR
 					(reg_q2150 AND symb_decoder(16#cf#)) OR
 					(reg_q2150 AND symb_decoder(16#85#)) OR
 					(reg_q2150 AND symb_decoder(16#75#)) OR
 					(reg_q2150 AND symb_decoder(16#fc#)) OR
 					(reg_q2150 AND symb_decoder(16#16#)) OR
 					(reg_q2150 AND symb_decoder(16#32#)) OR
 					(reg_q2150 AND symb_decoder(16#30#)) OR
 					(reg_q2150 AND symb_decoder(16#6a#)) OR
 					(reg_q2150 AND symb_decoder(16#34#)) OR
 					(reg_q2150 AND symb_decoder(16#66#)) OR
 					(reg_q2150 AND symb_decoder(16#f4#)) OR
 					(reg_q2150 AND symb_decoder(16#2a#)) OR
 					(reg_q2150 AND symb_decoder(16#20#)) OR
 					(reg_q2150 AND symb_decoder(16#e0#)) OR
 					(reg_q2150 AND symb_decoder(16#02#)) OR
 					(reg_q2150 AND symb_decoder(16#05#)) OR
 					(reg_q2150 AND symb_decoder(16#eb#)) OR
 					(reg_q2150 AND symb_decoder(16#e3#)) OR
 					(reg_q2150 AND symb_decoder(16#93#)) OR
 					(reg_q2150 AND symb_decoder(16#92#)) OR
 					(reg_q2150 AND symb_decoder(16#3c#)) OR
 					(reg_q2150 AND symb_decoder(16#73#)) OR
 					(reg_q2150 AND symb_decoder(16#bc#)) OR
 					(reg_q2150 AND symb_decoder(16#1a#)) OR
 					(reg_q2150 AND symb_decoder(16#d4#)) OR
 					(reg_q2150 AND symb_decoder(16#e2#)) OR
 					(reg_q2150 AND symb_decoder(16#c8#)) OR
 					(reg_q2150 AND symb_decoder(16#57#)) OR
 					(reg_q2150 AND symb_decoder(16#42#)) OR
 					(reg_q2150 AND symb_decoder(16#db#)) OR
 					(reg_q2150 AND symb_decoder(16#71#)) OR
 					(reg_q2150 AND symb_decoder(16#9e#)) OR
 					(reg_q2150 AND symb_decoder(16#f3#)) OR
 					(reg_q2150 AND symb_decoder(16#ee#)) OR
 					(reg_q2150 AND symb_decoder(16#3d#)) OR
 					(reg_q2150 AND symb_decoder(16#88#)) OR
 					(reg_q2150 AND symb_decoder(16#2d#)) OR
 					(reg_q2150 AND symb_decoder(16#76#)) OR
 					(reg_q2150 AND symb_decoder(16#b0#)) OR
 					(reg_q2150 AND symb_decoder(16#4b#)) OR
 					(reg_q2150 AND symb_decoder(16#d2#)) OR
 					(reg_q2150 AND symb_decoder(16#b5#)) OR
 					(reg_q2150 AND symb_decoder(16#98#)) OR
 					(reg_q2150 AND symb_decoder(16#9d#)) OR
 					(reg_q2150 AND symb_decoder(16#08#)) OR
 					(reg_q2150 AND symb_decoder(16#86#)) OR
 					(reg_q2150 AND symb_decoder(16#65#)) OR
 					(reg_q2150 AND symb_decoder(16#b9#)) OR
 					(reg_q2150 AND symb_decoder(16#68#)) OR
 					(reg_q2150 AND symb_decoder(16#7b#)) OR
 					(reg_q2150 AND symb_decoder(16#56#)) OR
 					(reg_q2150 AND symb_decoder(16#da#)) OR
 					(reg_q2150 AND symb_decoder(16#b2#)) OR
 					(reg_q2150 AND symb_decoder(16#0f#)) OR
 					(reg_q2150 AND symb_decoder(16#4c#)) OR
 					(reg_q2150 AND symb_decoder(16#1d#)) OR
 					(reg_q2150 AND symb_decoder(16#72#)) OR
 					(reg_q2150 AND symb_decoder(16#31#)) OR
 					(reg_q2150 AND symb_decoder(16#b7#)) OR
 					(reg_q2150 AND symb_decoder(16#af#)) OR
 					(reg_q2150 AND symb_decoder(16#04#)) OR
 					(reg_q2150 AND symb_decoder(16#4e#)) OR
 					(reg_q2150 AND symb_decoder(16#37#)) OR
 					(reg_q2150 AND symb_decoder(16#25#)) OR
 					(reg_q2150 AND symb_decoder(16#1b#)) OR
 					(reg_q2150 AND symb_decoder(16#7d#)) OR
 					(reg_q2150 AND symb_decoder(16#9b#)) OR
 					(reg_q2150 AND symb_decoder(16#7a#)) OR
 					(reg_q2150 AND symb_decoder(16#52#)) OR
 					(reg_q2150 AND symb_decoder(16#5f#)) OR
 					(reg_q2150 AND symb_decoder(16#3b#)) OR
 					(reg_q2150 AND symb_decoder(16#d7#)) OR
 					(reg_q2150 AND symb_decoder(16#d5#)) OR
 					(reg_q2150 AND symb_decoder(16#e7#)) OR
 					(reg_q2150 AND symb_decoder(16#ce#)) OR
 					(reg_q2150 AND symb_decoder(16#91#)) OR
 					(reg_q2150 AND symb_decoder(16#3e#)) OR
 					(reg_q2150 AND symb_decoder(16#b8#)) OR
 					(reg_q2150 AND symb_decoder(16#c1#)) OR
 					(reg_q2150 AND symb_decoder(16#c6#)) OR
 					(reg_q2150 AND symb_decoder(16#f9#)) OR
 					(reg_q2150 AND symb_decoder(16#64#)) OR
 					(reg_q2150 AND symb_decoder(16#a1#)) OR
 					(reg_q2150 AND symb_decoder(16#d1#)) OR
 					(reg_q2150 AND symb_decoder(16#f8#)) OR
 					(reg_q2150 AND symb_decoder(16#1f#)) OR
 					(reg_q2150 AND symb_decoder(16#e5#)) OR
 					(reg_q2150 AND symb_decoder(16#c9#)) OR
 					(reg_q2150 AND symb_decoder(16#cc#)) OR
 					(reg_q2150 AND symb_decoder(16#61#)) OR
 					(reg_q2150 AND symb_decoder(16#c5#)) OR
 					(reg_q2150 AND symb_decoder(16#51#)) OR
 					(reg_q2150 AND symb_decoder(16#17#)) OR
 					(reg_q2150 AND symb_decoder(16#69#)) OR
 					(reg_q2150 AND symb_decoder(16#f7#)) OR
 					(reg_q2150 AND symb_decoder(16#35#)) OR
 					(reg_q2150 AND symb_decoder(16#e9#)) OR
 					(reg_q2150 AND symb_decoder(16#87#)) OR
 					(reg_q2150 AND symb_decoder(16#b6#)) OR
 					(reg_q2150 AND symb_decoder(16#e4#)) OR
 					(reg_q2150 AND symb_decoder(16#d3#)) OR
 					(reg_q2150 AND symb_decoder(16#18#)) OR
 					(reg_q2150 AND symb_decoder(16#03#)) OR
 					(reg_q2150 AND symb_decoder(16#0c#)) OR
 					(reg_q2150 AND symb_decoder(16#6b#)) OR
 					(reg_q2150 AND symb_decoder(16#b1#)) OR
 					(reg_q2150 AND symb_decoder(16#80#)) OR
 					(reg_q2150 AND symb_decoder(16#14#)) OR
 					(reg_q2150 AND symb_decoder(16#9f#)) OR
 					(reg_q2150 AND symb_decoder(16#11#)) OR
 					(reg_q2150 AND symb_decoder(16#fa#)) OR
 					(reg_q2150 AND symb_decoder(16#c7#)) OR
 					(reg_q2150 AND symb_decoder(16#06#)) OR
 					(reg_q2150 AND symb_decoder(16#de#)) OR
 					(reg_q2150 AND symb_decoder(16#e8#)) OR
 					(reg_q2150 AND symb_decoder(16#a3#)) OR
 					(reg_q2150 AND symb_decoder(16#41#)) OR
 					(reg_q2150 AND symb_decoder(16#fe#)) OR
 					(reg_q2150 AND symb_decoder(16#28#)) OR
 					(reg_q2150 AND symb_decoder(16#82#)) OR
 					(reg_q2150 AND symb_decoder(16#c4#)) OR
 					(reg_q2150 AND symb_decoder(16#81#)) OR
 					(reg_q2150 AND symb_decoder(16#dc#)) OR
 					(reg_q2150 AND symb_decoder(16#ea#)) OR
 					(reg_q2150 AND symb_decoder(16#53#)) OR
 					(reg_q2150 AND symb_decoder(16#fb#)) OR
 					(reg_q2150 AND symb_decoder(16#97#)) OR
 					(reg_q2150 AND symb_decoder(16#77#)) OR
 					(reg_q2150 AND symb_decoder(16#29#)) OR
 					(reg_q2150 AND symb_decoder(16#c2#)) OR
 					(reg_q2150 AND symb_decoder(16#54#)) OR
 					(reg_q2150 AND symb_decoder(16#46#)) OR
 					(reg_q2150 AND symb_decoder(16#6d#)) OR
 					(reg_q2150 AND symb_decoder(16#70#)) OR
 					(reg_q2150 AND symb_decoder(16#74#)) OR
 					(reg_q2150 AND symb_decoder(16#36#)) OR
 					(reg_q2150 AND symb_decoder(16#4a#)) OR
 					(reg_q2150 AND symb_decoder(16#01#)) OR
 					(reg_q2150 AND symb_decoder(16#f0#)) OR
 					(reg_q2150 AND symb_decoder(16#58#)) OR
 					(reg_q2150 AND symb_decoder(16#12#)) OR
 					(reg_q2150 AND symb_decoder(16#55#)) OR
 					(reg_q2150 AND symb_decoder(16#45#)) OR
 					(reg_q2150 AND symb_decoder(16#15#)) OR
 					(reg_q2150 AND symb_decoder(16#f1#)) OR
 					(reg_q2150 AND symb_decoder(16#ae#)) OR
 					(reg_q2150 AND symb_decoder(16#ca#)) OR
 					(reg_q2150 AND symb_decoder(16#8b#)) OR
 					(reg_q2150 AND symb_decoder(16#8c#)) OR
 					(reg_q2150 AND symb_decoder(16#9c#)) OR
 					(reg_q2150 AND symb_decoder(16#dd#)) OR
 					(reg_q2150 AND symb_decoder(16#aa#)) OR
 					(reg_q2150 AND symb_decoder(16#78#)) OR
 					(reg_q2150 AND symb_decoder(16#2c#)) OR
 					(reg_q2150 AND symb_decoder(16#84#)) OR
 					(reg_q2150 AND symb_decoder(16#43#)) OR
 					(reg_q2150 AND symb_decoder(16#ef#)) OR
 					(reg_q2150 AND symb_decoder(16#a8#)) OR
 					(reg_q2150 AND symb_decoder(16#a4#)) OR
 					(reg_q2150 AND symb_decoder(16#5d#)) OR
 					(reg_q2150 AND symb_decoder(16#ba#)) OR
 					(reg_q2150 AND symb_decoder(16#79#)) OR
 					(reg_q2150 AND symb_decoder(16#33#)) OR
 					(reg_q2150 AND symb_decoder(16#8f#)) OR
 					(reg_q2150 AND symb_decoder(16#d0#)) OR
 					(reg_q2150 AND symb_decoder(16#ac#)) OR
 					(reg_q2150 AND symb_decoder(16#95#)) OR
 					(reg_q2150 AND symb_decoder(16#e1#)) OR
 					(reg_q2150 AND symb_decoder(16#ff#)) OR
 					(reg_q2150 AND symb_decoder(16#90#)) OR
 					(reg_q2150 AND symb_decoder(16#26#)) OR
 					(reg_q2150 AND symb_decoder(16#cd#)) OR
 					(reg_q2150 AND symb_decoder(16#5e#)) OR
 					(reg_q2150 AND symb_decoder(16#ec#)) OR
 					(reg_q2150 AND symb_decoder(16#8e#)) OR
 					(reg_q2150 AND symb_decoder(16#24#)) OR
 					(reg_q2150 AND symb_decoder(16#89#)) OR
 					(reg_q2150 AND symb_decoder(16#2e#)) OR
 					(reg_q2150 AND symb_decoder(16#a9#)) OR
 					(reg_q2150 AND symb_decoder(16#df#)) OR
 					(reg_q2150 AND symb_decoder(16#50#)) OR
 					(reg_q2150 AND symb_decoder(16#59#)) OR
 					(reg_q2150 AND symb_decoder(16#a0#)) OR
 					(reg_q2150 AND symb_decoder(16#2f#)) OR
 					(reg_q2150 AND symb_decoder(16#09#)) OR
 					(reg_q2150 AND symb_decoder(16#bf#)) OR
 					(reg_q2150 AND symb_decoder(16#07#)) OR
 					(reg_q2150 AND symb_decoder(16#7f#)) OR
 					(reg_q2150 AND symb_decoder(16#cb#)) OR
 					(reg_q2150 AND symb_decoder(16#94#)) OR
 					(reg_q2150 AND symb_decoder(16#9a#)) OR
 					(reg_q2150 AND symb_decoder(16#d6#)) OR
 					(reg_q2150 AND symb_decoder(16#40#)) OR
 					(reg_q2150 AND symb_decoder(16#38#)) OR
 					(reg_q2150 AND symb_decoder(16#a5#)) OR
 					(reg_q2150 AND symb_decoder(16#5b#)) OR
 					(reg_q2150 AND symb_decoder(16#f2#)) OR
 					(reg_q2150 AND symb_decoder(16#5a#)) OR
 					(reg_q2150 AND symb_decoder(16#2b#)) OR
 					(reg_q2150 AND symb_decoder(16#67#)) OR
 					(reg_q2150 AND symb_decoder(16#1c#)) OR
 					(reg_q2150 AND symb_decoder(16#22#));
reg_q117_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q116 AND symb_decoder(16#0a#)) OR
 					(reg_q116 AND symb_decoder(16#0d#));
reg_q805_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q804 AND symb_decoder(16#53#)) OR
 					(reg_q804 AND symb_decoder(16#73#));
reg_fullgraph38_init <= "00";

reg_fullgraph38_sel <= "0" & reg_q805_in & reg_q117_in & reg_q2216_in;

	--coder fullgraph38
with reg_fullgraph38_sel select
reg_fullgraph38_in <=
	"01" when "0001",
	"10" when "0010",
	"11" when "0100",
	"00" when others;
 --end coder

	p_reg_fullgraph38: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph38 <= reg_fullgraph38_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph38 <= reg_fullgraph38_init;
        else
          reg_fullgraph38 <= reg_fullgraph38_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph38

		reg_q2216 <= '1' when reg_fullgraph38 = "01" else '0'; 
		reg_q117 <= '1' when reg_fullgraph38 = "10" else '0'; 
		reg_q805 <= '1' when reg_fullgraph38 = "11" else '0'; 
--end decoder 
--######################################################
--fullgraph39

reg_q397_in <= (reg_q359 AND symb_decoder(16#c3#)) OR
 					(reg_q359 AND symb_decoder(16#15#)) OR
 					(reg_q359 AND symb_decoder(16#fb#)) OR
 					(reg_q359 AND symb_decoder(16#fd#)) OR
 					(reg_q359 AND symb_decoder(16#8d#)) OR
 					(reg_q359 AND symb_decoder(16#b5#)) OR
 					(reg_q359 AND symb_decoder(16#07#)) OR
 					(reg_q359 AND symb_decoder(16#9a#)) OR
 					(reg_q359 AND symb_decoder(16#b8#)) OR
 					(reg_q359 AND symb_decoder(16#2c#)) OR
 					(reg_q359 AND symb_decoder(16#e6#)) OR
 					(reg_q359 AND symb_decoder(16#94#)) OR
 					(reg_q359 AND symb_decoder(16#37#)) OR
 					(reg_q359 AND symb_decoder(16#36#)) OR
 					(reg_q359 AND symb_decoder(16#74#)) OR
 					(reg_q359 AND symb_decoder(16#1d#)) OR
 					(reg_q359 AND symb_decoder(16#6c#)) OR
 					(reg_q359 AND symb_decoder(16#b4#)) OR
 					(reg_q359 AND symb_decoder(16#0e#)) OR
 					(reg_q359 AND symb_decoder(16#97#)) OR
 					(reg_q359 AND symb_decoder(16#c2#)) OR
 					(reg_q359 AND symb_decoder(16#4c#)) OR
 					(reg_q359 AND symb_decoder(16#f4#)) OR
 					(reg_q359 AND symb_decoder(16#e1#)) OR
 					(reg_q359 AND symb_decoder(16#f5#)) OR
 					(reg_q359 AND symb_decoder(16#6d#)) OR
 					(reg_q359 AND symb_decoder(16#a8#)) OR
 					(reg_q359 AND symb_decoder(16#26#)) OR
 					(reg_q359 AND symb_decoder(16#ed#)) OR
 					(reg_q359 AND symb_decoder(16#b3#)) OR
 					(reg_q359 AND symb_decoder(16#f9#)) OR
 					(reg_q359 AND symb_decoder(16#f1#)) OR
 					(reg_q359 AND symb_decoder(16#a2#)) OR
 					(reg_q359 AND symb_decoder(16#c4#)) OR
 					(reg_q359 AND symb_decoder(16#a3#)) OR
 					(reg_q359 AND symb_decoder(16#80#)) OR
 					(reg_q359 AND symb_decoder(16#34#)) OR
 					(reg_q359 AND symb_decoder(16#14#)) OR
 					(reg_q359 AND symb_decoder(16#b7#)) OR
 					(reg_q359 AND symb_decoder(16#aa#)) OR
 					(reg_q359 AND symb_decoder(16#62#)) OR
 					(reg_q359 AND symb_decoder(16#08#)) OR
 					(reg_q359 AND symb_decoder(16#7f#)) OR
 					(reg_q359 AND symb_decoder(16#8a#)) OR
 					(reg_q359 AND symb_decoder(16#4d#)) OR
 					(reg_q359 AND symb_decoder(16#ab#)) OR
 					(reg_q359 AND symb_decoder(16#40#)) OR
 					(reg_q359 AND symb_decoder(16#ce#)) OR
 					(reg_q359 AND symb_decoder(16#7a#)) OR
 					(reg_q359 AND symb_decoder(16#ff#)) OR
 					(reg_q359 AND symb_decoder(16#c6#)) OR
 					(reg_q359 AND symb_decoder(16#95#)) OR
 					(reg_q359 AND symb_decoder(16#c1#)) OR
 					(reg_q359 AND symb_decoder(16#5f#)) OR
 					(reg_q359 AND symb_decoder(16#a0#)) OR
 					(reg_q359 AND symb_decoder(16#20#)) OR
 					(reg_q359 AND symb_decoder(16#a7#)) OR
 					(reg_q359 AND symb_decoder(16#99#)) OR
 					(reg_q359 AND symb_decoder(16#e2#)) OR
 					(reg_q359 AND symb_decoder(16#f0#)) OR
 					(reg_q359 AND symb_decoder(16#3f#)) OR
 					(reg_q359 AND symb_decoder(16#c8#)) OR
 					(reg_q359 AND symb_decoder(16#e0#)) OR
 					(reg_q359 AND symb_decoder(16#6f#)) OR
 					(reg_q359 AND symb_decoder(16#d5#)) OR
 					(reg_q359 AND symb_decoder(16#8b#)) OR
 					(reg_q359 AND symb_decoder(16#1c#)) OR
 					(reg_q359 AND symb_decoder(16#32#)) OR
 					(reg_q359 AND symb_decoder(16#30#)) OR
 					(reg_q359 AND symb_decoder(16#f6#)) OR
 					(reg_q359 AND symb_decoder(16#db#)) OR
 					(reg_q359 AND symb_decoder(16#cb#)) OR
 					(reg_q359 AND symb_decoder(16#f7#)) OR
 					(reg_q359 AND symb_decoder(16#48#)) OR
 					(reg_q359 AND symb_decoder(16#52#)) OR
 					(reg_q359 AND symb_decoder(16#d0#)) OR
 					(reg_q359 AND symb_decoder(16#38#)) OR
 					(reg_q359 AND symb_decoder(16#4e#)) OR
 					(reg_q359 AND symb_decoder(16#2b#)) OR
 					(reg_q359 AND symb_decoder(16#bb#)) OR
 					(reg_q359 AND symb_decoder(16#c7#)) OR
 					(reg_q359 AND symb_decoder(16#67#)) OR
 					(reg_q359 AND symb_decoder(16#e7#)) OR
 					(reg_q359 AND symb_decoder(16#68#)) OR
 					(reg_q359 AND symb_decoder(16#5b#)) OR
 					(reg_q359 AND symb_decoder(16#d2#)) OR
 					(reg_q359 AND symb_decoder(16#33#)) OR
 					(reg_q359 AND symb_decoder(16#89#)) OR
 					(reg_q359 AND symb_decoder(16#8c#)) OR
 					(reg_q359 AND symb_decoder(16#a9#)) OR
 					(reg_q359 AND symb_decoder(16#0c#)) OR
 					(reg_q359 AND symb_decoder(16#46#)) OR
 					(reg_q359 AND symb_decoder(16#e5#)) OR
 					(reg_q359 AND symb_decoder(16#42#)) OR
 					(reg_q359 AND symb_decoder(16#ca#)) OR
 					(reg_q359 AND symb_decoder(16#24#)) OR
 					(reg_q359 AND symb_decoder(16#4a#)) OR
 					(reg_q359 AND symb_decoder(16#11#)) OR
 					(reg_q359 AND symb_decoder(16#b1#)) OR
 					(reg_q359 AND symb_decoder(16#4f#)) OR
 					(reg_q359 AND symb_decoder(16#53#)) OR
 					(reg_q359 AND symb_decoder(16#81#)) OR
 					(reg_q359 AND symb_decoder(16#59#)) OR
 					(reg_q359 AND symb_decoder(16#55#)) OR
 					(reg_q359 AND symb_decoder(16#df#)) OR
 					(reg_q359 AND symb_decoder(16#2f#)) OR
 					(reg_q359 AND symb_decoder(16#96#)) OR
 					(reg_q359 AND symb_decoder(16#01#)) OR
 					(reg_q359 AND symb_decoder(16#45#)) OR
 					(reg_q359 AND symb_decoder(16#02#)) OR
 					(reg_q359 AND symb_decoder(16#9d#)) OR
 					(reg_q359 AND symb_decoder(16#0f#)) OR
 					(reg_q359 AND symb_decoder(16#7c#)) OR
 					(reg_q359 AND symb_decoder(16#3b#)) OR
 					(reg_q359 AND symb_decoder(16#09#)) OR
 					(reg_q359 AND symb_decoder(16#18#)) OR
 					(reg_q359 AND symb_decoder(16#de#)) OR
 					(reg_q359 AND symb_decoder(16#1e#)) OR
 					(reg_q359 AND symb_decoder(16#9f#)) OR
 					(reg_q359 AND symb_decoder(16#12#)) OR
 					(reg_q359 AND symb_decoder(16#04#)) OR
 					(reg_q359 AND symb_decoder(16#1a#)) OR
 					(reg_q359 AND symb_decoder(16#6b#)) OR
 					(reg_q359 AND symb_decoder(16#f8#)) OR
 					(reg_q359 AND symb_decoder(16#71#)) OR
 					(reg_q359 AND symb_decoder(16#91#)) OR
 					(reg_q359 AND symb_decoder(16#65#)) OR
 					(reg_q359 AND symb_decoder(16#4b#)) OR
 					(reg_q359 AND symb_decoder(16#49#)) OR
 					(reg_q359 AND symb_decoder(16#8f#)) OR
 					(reg_q359 AND symb_decoder(16#e3#)) OR
 					(reg_q359 AND symb_decoder(16#6a#)) OR
 					(reg_q359 AND symb_decoder(16#2e#)) OR
 					(reg_q359 AND symb_decoder(16#78#)) OR
 					(reg_q359 AND symb_decoder(16#d9#)) OR
 					(reg_q359 AND symb_decoder(16#84#)) OR
 					(reg_q359 AND symb_decoder(16#93#)) OR
 					(reg_q359 AND symb_decoder(16#d3#)) OR
 					(reg_q359 AND symb_decoder(16#a4#)) OR
 					(reg_q359 AND symb_decoder(16#88#)) OR
 					(reg_q359 AND symb_decoder(16#27#)) OR
 					(reg_q359 AND symb_decoder(16#cc#)) OR
 					(reg_q359 AND symb_decoder(16#ad#)) OR
 					(reg_q359 AND symb_decoder(16#b6#)) OR
 					(reg_q359 AND symb_decoder(16#a1#)) OR
 					(reg_q359 AND symb_decoder(16#05#)) OR
 					(reg_q359 AND symb_decoder(16#ba#)) OR
 					(reg_q359 AND symb_decoder(16#66#)) OR
 					(reg_q359 AND symb_decoder(16#d6#)) OR
 					(reg_q359 AND symb_decoder(16#9e#)) OR
 					(reg_q359 AND symb_decoder(16#35#)) OR
 					(reg_q359 AND symb_decoder(16#50#)) OR
 					(reg_q359 AND symb_decoder(16#3c#)) OR
 					(reg_q359 AND symb_decoder(16#85#)) OR
 					(reg_q359 AND symb_decoder(16#60#)) OR
 					(reg_q359 AND symb_decoder(16#72#)) OR
 					(reg_q359 AND symb_decoder(16#eb#)) OR
 					(reg_q359 AND symb_decoder(16#83#)) OR
 					(reg_q359 AND symb_decoder(16#17#)) OR
 					(reg_q359 AND symb_decoder(16#bc#)) OR
 					(reg_q359 AND symb_decoder(16#61#)) OR
 					(reg_q359 AND symb_decoder(16#bf#)) OR
 					(reg_q359 AND symb_decoder(16#c0#)) OR
 					(reg_q359 AND symb_decoder(16#25#)) OR
 					(reg_q359 AND symb_decoder(16#e8#)) OR
 					(reg_q359 AND symb_decoder(16#16#)) OR
 					(reg_q359 AND symb_decoder(16#79#)) OR
 					(reg_q359 AND symb_decoder(16#d1#)) OR
 					(reg_q359 AND symb_decoder(16#3e#)) OR
 					(reg_q359 AND symb_decoder(16#54#)) OR
 					(reg_q359 AND symb_decoder(16#d8#)) OR
 					(reg_q359 AND symb_decoder(16#64#)) OR
 					(reg_q359 AND symb_decoder(16#d4#)) OR
 					(reg_q359 AND symb_decoder(16#87#)) OR
 					(reg_q359 AND symb_decoder(16#f3#)) OR
 					(reg_q359 AND symb_decoder(16#c9#)) OR
 					(reg_q359 AND symb_decoder(16#fe#)) OR
 					(reg_q359 AND symb_decoder(16#b2#)) OR
 					(reg_q359 AND symb_decoder(16#13#)) OR
 					(reg_q359 AND symb_decoder(16#f2#)) OR
 					(reg_q359 AND symb_decoder(16#92#)) OR
 					(reg_q359 AND symb_decoder(16#03#)) OR
 					(reg_q359 AND symb_decoder(16#21#)) OR
 					(reg_q359 AND symb_decoder(16#51#)) OR
 					(reg_q359 AND symb_decoder(16#8e#)) OR
 					(reg_q359 AND symb_decoder(16#31#)) OR
 					(reg_q359 AND symb_decoder(16#77#)) OR
 					(reg_q359 AND symb_decoder(16#be#)) OR
 					(reg_q359 AND symb_decoder(16#86#)) OR
 					(reg_q359 AND symb_decoder(16#fa#)) OR
 					(reg_q359 AND symb_decoder(16#57#)) OR
 					(reg_q359 AND symb_decoder(16#56#)) OR
 					(reg_q359 AND symb_decoder(16#5c#)) OR
 					(reg_q359 AND symb_decoder(16#9c#)) OR
 					(reg_q359 AND symb_decoder(16#a6#)) OR
 					(reg_q359 AND symb_decoder(16#22#)) OR
 					(reg_q359 AND symb_decoder(16#5a#)) OR
 					(reg_q359 AND symb_decoder(16#90#)) OR
 					(reg_q359 AND symb_decoder(16#76#)) OR
 					(reg_q359 AND symb_decoder(16#00#)) OR
 					(reg_q359 AND symb_decoder(16#a5#)) OR
 					(reg_q359 AND symb_decoder(16#b0#)) OR
 					(reg_q359 AND symb_decoder(16#19#)) OR
 					(reg_q359 AND symb_decoder(16#c5#)) OR
 					(reg_q359 AND symb_decoder(16#d7#)) OR
 					(reg_q359 AND symb_decoder(16#7b#)) OR
 					(reg_q359 AND symb_decoder(16#0b#)) OR
 					(reg_q359 AND symb_decoder(16#73#)) OR
 					(reg_q359 AND symb_decoder(16#7d#)) OR
 					(reg_q359 AND symb_decoder(16#69#)) OR
 					(reg_q359 AND symb_decoder(16#da#)) OR
 					(reg_q359 AND symb_decoder(16#39#)) OR
 					(reg_q359 AND symb_decoder(16#47#)) OR
 					(reg_q359 AND symb_decoder(16#e4#)) OR
 					(reg_q359 AND symb_decoder(16#28#)) OR
 					(reg_q359 AND symb_decoder(16#9b#)) OR
 					(reg_q359 AND symb_decoder(16#82#)) OR
 					(reg_q359 AND symb_decoder(16#29#)) OR
 					(reg_q359 AND symb_decoder(16#cd#)) OR
 					(reg_q359 AND symb_decoder(16#cf#)) OR
 					(reg_q359 AND symb_decoder(16#23#)) OR
 					(reg_q359 AND symb_decoder(16#ec#)) OR
 					(reg_q359 AND symb_decoder(16#43#)) OR
 					(reg_q359 AND symb_decoder(16#6e#)) OR
 					(reg_q359 AND symb_decoder(16#ac#)) OR
 					(reg_q359 AND symb_decoder(16#ee#)) OR
 					(reg_q359 AND symb_decoder(16#bd#)) OR
 					(reg_q359 AND symb_decoder(16#3a#)) OR
 					(reg_q359 AND symb_decoder(16#1f#)) OR
 					(reg_q359 AND symb_decoder(16#2a#)) OR
 					(reg_q359 AND symb_decoder(16#06#)) OR
 					(reg_q359 AND symb_decoder(16#63#)) OR
 					(reg_q359 AND symb_decoder(16#3d#)) OR
 					(reg_q359 AND symb_decoder(16#5d#)) OR
 					(reg_q359 AND symb_decoder(16#ae#)) OR
 					(reg_q359 AND symb_decoder(16#58#)) OR
 					(reg_q359 AND symb_decoder(16#44#)) OR
 					(reg_q359 AND symb_decoder(16#ea#)) OR
 					(reg_q359 AND symb_decoder(16#98#)) OR
 					(reg_q359 AND symb_decoder(16#af#)) OR
 					(reg_q359 AND symb_decoder(16#2d#)) OR
 					(reg_q359 AND symb_decoder(16#70#)) OR
 					(reg_q359 AND symb_decoder(16#7e#)) OR
 					(reg_q359 AND symb_decoder(16#5e#)) OR
 					(reg_q359 AND symb_decoder(16#ef#)) OR
 					(reg_q359 AND symb_decoder(16#10#)) OR
 					(reg_q359 AND symb_decoder(16#b9#)) OR
 					(reg_q359 AND symb_decoder(16#fc#)) OR
 					(reg_q359 AND symb_decoder(16#e9#)) OR
 					(reg_q359 AND symb_decoder(16#75#)) OR
 					(reg_q359 AND symb_decoder(16#dd#)) OR
 					(reg_q359 AND symb_decoder(16#dc#)) OR
 					(reg_q359 AND symb_decoder(16#1b#)) OR
 					(reg_q359 AND symb_decoder(16#41#)) OR
 					(reg_q397 AND symb_decoder(16#24#)) OR
 					(reg_q397 AND symb_decoder(16#34#)) OR
 					(reg_q397 AND symb_decoder(16#51#)) OR
 					(reg_q397 AND symb_decoder(16#2e#)) OR
 					(reg_q397 AND symb_decoder(16#59#)) OR
 					(reg_q397 AND symb_decoder(16#f1#)) OR
 					(reg_q397 AND symb_decoder(16#ea#)) OR
 					(reg_q397 AND symb_decoder(16#20#)) OR
 					(reg_q397 AND symb_decoder(16#e0#)) OR
 					(reg_q397 AND symb_decoder(16#ca#)) OR
 					(reg_q397 AND symb_decoder(16#5c#)) OR
 					(reg_q397 AND symb_decoder(16#9b#)) OR
 					(reg_q397 AND symb_decoder(16#14#)) OR
 					(reg_q397 AND symb_decoder(16#c2#)) OR
 					(reg_q397 AND symb_decoder(16#d6#)) OR
 					(reg_q397 AND symb_decoder(16#e1#)) OR
 					(reg_q397 AND symb_decoder(16#df#)) OR
 					(reg_q397 AND symb_decoder(16#75#)) OR
 					(reg_q397 AND symb_decoder(16#ff#)) OR
 					(reg_q397 AND symb_decoder(16#61#)) OR
 					(reg_q397 AND symb_decoder(16#00#)) OR
 					(reg_q397 AND symb_decoder(16#b2#)) OR
 					(reg_q397 AND symb_decoder(16#6a#)) OR
 					(reg_q397 AND symb_decoder(16#1a#)) OR
 					(reg_q397 AND symb_decoder(16#1c#)) OR
 					(reg_q397 AND symb_decoder(16#f9#)) OR
 					(reg_q397 AND symb_decoder(16#77#)) OR
 					(reg_q397 AND symb_decoder(16#07#)) OR
 					(reg_q397 AND symb_decoder(16#65#)) OR
 					(reg_q397 AND symb_decoder(16#ac#)) OR
 					(reg_q397 AND symb_decoder(16#e4#)) OR
 					(reg_q397 AND symb_decoder(16#ce#)) OR
 					(reg_q397 AND symb_decoder(16#d7#)) OR
 					(reg_q397 AND symb_decoder(16#af#)) OR
 					(reg_q397 AND symb_decoder(16#cc#)) OR
 					(reg_q397 AND symb_decoder(16#3c#)) OR
 					(reg_q397 AND symb_decoder(16#3f#)) OR
 					(reg_q397 AND symb_decoder(16#9c#)) OR
 					(reg_q397 AND symb_decoder(16#02#)) OR
 					(reg_q397 AND symb_decoder(16#ad#)) OR
 					(reg_q397 AND symb_decoder(16#18#)) OR
 					(reg_q397 AND symb_decoder(16#7a#)) OR
 					(reg_q397 AND symb_decoder(16#79#)) OR
 					(reg_q397 AND symb_decoder(16#c0#)) OR
 					(reg_q397 AND symb_decoder(16#0c#)) OR
 					(reg_q397 AND symb_decoder(16#85#)) OR
 					(reg_q397 AND symb_decoder(16#87#)) OR
 					(reg_q397 AND symb_decoder(16#7d#)) OR
 					(reg_q397 AND symb_decoder(16#3e#)) OR
 					(reg_q397 AND symb_decoder(16#aa#)) OR
 					(reg_q397 AND symb_decoder(16#ec#)) OR
 					(reg_q397 AND symb_decoder(16#31#)) OR
 					(reg_q397 AND symb_decoder(16#4f#)) OR
 					(reg_q397 AND symb_decoder(16#21#)) OR
 					(reg_q397 AND symb_decoder(16#5b#)) OR
 					(reg_q397 AND symb_decoder(16#fe#)) OR
 					(reg_q397 AND symb_decoder(16#d4#)) OR
 					(reg_q397 AND symb_decoder(16#ab#)) OR
 					(reg_q397 AND symb_decoder(16#99#)) OR
 					(reg_q397 AND symb_decoder(16#6d#)) OR
 					(reg_q397 AND symb_decoder(16#04#)) OR
 					(reg_q397 AND symb_decoder(16#80#)) OR
 					(reg_q397 AND symb_decoder(16#5d#)) OR
 					(reg_q397 AND symb_decoder(16#3d#)) OR
 					(reg_q397 AND symb_decoder(16#68#)) OR
 					(reg_q397 AND symb_decoder(16#63#)) OR
 					(reg_q397 AND symb_decoder(16#6c#)) OR
 					(reg_q397 AND symb_decoder(16#bd#)) OR
 					(reg_q397 AND symb_decoder(16#e3#)) OR
 					(reg_q397 AND symb_decoder(16#d5#)) OR
 					(reg_q397 AND symb_decoder(16#54#)) OR
 					(reg_q397 AND symb_decoder(16#94#)) OR
 					(reg_q397 AND symb_decoder(16#90#)) OR
 					(reg_q397 AND symb_decoder(16#0e#)) OR
 					(reg_q397 AND symb_decoder(16#d9#)) OR
 					(reg_q397 AND symb_decoder(16#de#)) OR
 					(reg_q397 AND symb_decoder(16#40#)) OR
 					(reg_q397 AND symb_decoder(16#06#)) OR
 					(reg_q397 AND symb_decoder(16#47#)) OR
 					(reg_q397 AND symb_decoder(16#82#)) OR
 					(reg_q397 AND symb_decoder(16#23#)) OR
 					(reg_q397 AND symb_decoder(16#8a#)) OR
 					(reg_q397 AND symb_decoder(16#45#)) OR
 					(reg_q397 AND symb_decoder(16#74#)) OR
 					(reg_q397 AND symb_decoder(16#bc#)) OR
 					(reg_q397 AND symb_decoder(16#60#)) OR
 					(reg_q397 AND symb_decoder(16#72#)) OR
 					(reg_q397 AND symb_decoder(16#d8#)) OR
 					(reg_q397 AND symb_decoder(16#fd#)) OR
 					(reg_q397 AND symb_decoder(16#52#)) OR
 					(reg_q397 AND symb_decoder(16#2f#)) OR
 					(reg_q397 AND symb_decoder(16#73#)) OR
 					(reg_q397 AND symb_decoder(16#c4#)) OR
 					(reg_q397 AND symb_decoder(16#6b#)) OR
 					(reg_q397 AND symb_decoder(16#ba#)) OR
 					(reg_q397 AND symb_decoder(16#a0#)) OR
 					(reg_q397 AND symb_decoder(16#9f#)) OR
 					(reg_q397 AND symb_decoder(16#81#)) OR
 					(reg_q397 AND symb_decoder(16#13#)) OR
 					(reg_q397 AND symb_decoder(16#4c#)) OR
 					(reg_q397 AND symb_decoder(16#b6#)) OR
 					(reg_q397 AND symb_decoder(16#30#)) OR
 					(reg_q397 AND symb_decoder(16#e9#)) OR
 					(reg_q397 AND symb_decoder(16#fc#)) OR
 					(reg_q397 AND symb_decoder(16#95#)) OR
 					(reg_q397 AND symb_decoder(16#41#)) OR
 					(reg_q397 AND symb_decoder(16#10#)) OR
 					(reg_q397 AND symb_decoder(16#e6#)) OR
 					(reg_q397 AND symb_decoder(16#cd#)) OR
 					(reg_q397 AND symb_decoder(16#8c#)) OR
 					(reg_q397 AND symb_decoder(16#4e#)) OR
 					(reg_q397 AND symb_decoder(16#b1#)) OR
 					(reg_q397 AND symb_decoder(16#6e#)) OR
 					(reg_q397 AND symb_decoder(16#03#)) OR
 					(reg_q397 AND symb_decoder(16#be#)) OR
 					(reg_q397 AND symb_decoder(16#c5#)) OR
 					(reg_q397 AND symb_decoder(16#83#)) OR
 					(reg_q397 AND symb_decoder(16#a7#)) OR
 					(reg_q397 AND symb_decoder(16#ed#)) OR
 					(reg_q397 AND symb_decoder(16#a3#)) OR
 					(reg_q397 AND symb_decoder(16#78#)) OR
 					(reg_q397 AND symb_decoder(16#69#)) OR
 					(reg_q397 AND symb_decoder(16#1e#)) OR
 					(reg_q397 AND symb_decoder(16#d1#)) OR
 					(reg_q397 AND symb_decoder(16#33#)) OR
 					(reg_q397 AND symb_decoder(16#86#)) OR
 					(reg_q397 AND symb_decoder(16#5a#)) OR
 					(reg_q397 AND symb_decoder(16#c7#)) OR
 					(reg_q397 AND symb_decoder(16#89#)) OR
 					(reg_q397 AND symb_decoder(16#7f#)) OR
 					(reg_q397 AND symb_decoder(16#0f#)) OR
 					(reg_q397 AND symb_decoder(16#44#)) OR
 					(reg_q397 AND symb_decoder(16#8e#)) OR
 					(reg_q397 AND symb_decoder(16#bf#)) OR
 					(reg_q397 AND symb_decoder(16#12#)) OR
 					(reg_q397 AND symb_decoder(16#28#)) OR
 					(reg_q397 AND symb_decoder(16#97#)) OR
 					(reg_q397 AND symb_decoder(16#b0#)) OR
 					(reg_q397 AND symb_decoder(16#42#)) OR
 					(reg_q397 AND symb_decoder(16#8d#)) OR
 					(reg_q397 AND symb_decoder(16#50#)) OR
 					(reg_q397 AND symb_decoder(16#c3#)) OR
 					(reg_q397 AND symb_decoder(16#0b#)) OR
 					(reg_q397 AND symb_decoder(16#15#)) OR
 					(reg_q397 AND symb_decoder(16#4b#)) OR
 					(reg_q397 AND symb_decoder(16#8b#)) OR
 					(reg_q397 AND symb_decoder(16#92#)) OR
 					(reg_q397 AND symb_decoder(16#b3#)) OR
 					(reg_q397 AND symb_decoder(16#1f#)) OR
 					(reg_q397 AND symb_decoder(16#56#)) OR
 					(reg_q397 AND symb_decoder(16#9e#)) OR
 					(reg_q397 AND symb_decoder(16#da#)) OR
 					(reg_q397 AND symb_decoder(16#e5#)) OR
 					(reg_q397 AND symb_decoder(16#9a#)) OR
 					(reg_q397 AND symb_decoder(16#cb#)) OR
 					(reg_q397 AND symb_decoder(16#09#)) OR
 					(reg_q397 AND symb_decoder(16#b4#)) OR
 					(reg_q397 AND symb_decoder(16#dd#)) OR
 					(reg_q397 AND symb_decoder(16#96#)) OR
 					(reg_q397 AND symb_decoder(16#db#)) OR
 					(reg_q397 AND symb_decoder(16#b9#)) OR
 					(reg_q397 AND symb_decoder(16#c1#)) OR
 					(reg_q397 AND symb_decoder(16#17#)) OR
 					(reg_q397 AND symb_decoder(16#f7#)) OR
 					(reg_q397 AND symb_decoder(16#3a#)) OR
 					(reg_q397 AND symb_decoder(16#c6#)) OR
 					(reg_q397 AND symb_decoder(16#35#)) OR
 					(reg_q397 AND symb_decoder(16#2d#)) OR
 					(reg_q397 AND symb_decoder(16#d3#)) OR
 					(reg_q397 AND symb_decoder(16#ef#)) OR
 					(reg_q397 AND symb_decoder(16#a6#)) OR
 					(reg_q397 AND symb_decoder(16#eb#)) OR
 					(reg_q397 AND symb_decoder(16#27#)) OR
 					(reg_q397 AND symb_decoder(16#39#)) OR
 					(reg_q397 AND symb_decoder(16#66#)) OR
 					(reg_q397 AND symb_decoder(16#e7#)) OR
 					(reg_q397 AND symb_decoder(16#a9#)) OR
 					(reg_q397 AND symb_decoder(16#1b#)) OR
 					(reg_q397 AND symb_decoder(16#64#)) OR
 					(reg_q397 AND symb_decoder(16#5e#)) OR
 					(reg_q397 AND symb_decoder(16#f0#)) OR
 					(reg_q397 AND symb_decoder(16#2a#)) OR
 					(reg_q397 AND symb_decoder(16#29#)) OR
 					(reg_q397 AND symb_decoder(16#84#)) OR
 					(reg_q397 AND symb_decoder(16#25#)) OR
 					(reg_q397 AND symb_decoder(16#2b#)) OR
 					(reg_q397 AND symb_decoder(16#11#)) OR
 					(reg_q397 AND symb_decoder(16#cf#)) OR
 					(reg_q397 AND symb_decoder(16#01#)) OR
 					(reg_q397 AND symb_decoder(16#62#)) OR
 					(reg_q397 AND symb_decoder(16#36#)) OR
 					(reg_q397 AND symb_decoder(16#b7#)) OR
 					(reg_q397 AND symb_decoder(16#8f#)) OR
 					(reg_q397 AND symb_decoder(16#08#)) OR
 					(reg_q397 AND symb_decoder(16#7e#)) OR
 					(reg_q397 AND symb_decoder(16#55#)) OR
 					(reg_q397 AND symb_decoder(16#c8#)) OR
 					(reg_q397 AND symb_decoder(16#f2#)) OR
 					(reg_q397 AND symb_decoder(16#f3#)) OR
 					(reg_q397 AND symb_decoder(16#7c#)) OR
 					(reg_q397 AND symb_decoder(16#98#)) OR
 					(reg_q397 AND symb_decoder(16#c9#)) OR
 					(reg_q397 AND symb_decoder(16#a1#)) OR
 					(reg_q397 AND symb_decoder(16#b5#)) OR
 					(reg_q397 AND symb_decoder(16#e2#)) OR
 					(reg_q397 AND symb_decoder(16#d0#)) OR
 					(reg_q397 AND symb_decoder(16#05#)) OR
 					(reg_q397 AND symb_decoder(16#76#)) OR
 					(reg_q397 AND symb_decoder(16#f5#)) OR
 					(reg_q397 AND symb_decoder(16#4d#)) OR
 					(reg_q397 AND symb_decoder(16#9d#)) OR
 					(reg_q397 AND symb_decoder(16#19#)) OR
 					(reg_q397 AND symb_decoder(16#38#)) OR
 					(reg_q397 AND symb_decoder(16#f4#)) OR
 					(reg_q397 AND symb_decoder(16#48#)) OR
 					(reg_q397 AND symb_decoder(16#26#)) OR
 					(reg_q397 AND symb_decoder(16#fb#)) OR
 					(reg_q397 AND symb_decoder(16#1d#)) OR
 					(reg_q397 AND symb_decoder(16#a4#)) OR
 					(reg_q397 AND symb_decoder(16#3b#)) OR
 					(reg_q397 AND symb_decoder(16#5f#)) OR
 					(reg_q397 AND symb_decoder(16#57#)) OR
 					(reg_q397 AND symb_decoder(16#dc#)) OR
 					(reg_q397 AND symb_decoder(16#46#)) OR
 					(reg_q397 AND symb_decoder(16#4a#)) OR
 					(reg_q397 AND symb_decoder(16#bb#)) OR
 					(reg_q397 AND symb_decoder(16#f6#)) OR
 					(reg_q397 AND symb_decoder(16#a8#)) OR
 					(reg_q397 AND symb_decoder(16#b8#)) OR
 					(reg_q397 AND symb_decoder(16#a2#)) OR
 					(reg_q397 AND symb_decoder(16#49#)) OR
 					(reg_q397 AND symb_decoder(16#f8#)) OR
 					(reg_q397 AND symb_decoder(16#22#)) OR
 					(reg_q397 AND symb_decoder(16#91#)) OR
 					(reg_q397 AND symb_decoder(16#2c#)) OR
 					(reg_q397 AND symb_decoder(16#67#)) OR
 					(reg_q397 AND symb_decoder(16#a5#)) OR
 					(reg_q397 AND symb_decoder(16#58#)) OR
 					(reg_q397 AND symb_decoder(16#6f#)) OR
 					(reg_q397 AND symb_decoder(16#70#)) OR
 					(reg_q397 AND symb_decoder(16#71#)) OR
 					(reg_q397 AND symb_decoder(16#93#)) OR
 					(reg_q397 AND symb_decoder(16#ae#)) OR
 					(reg_q397 AND symb_decoder(16#d2#)) OR
 					(reg_q397 AND symb_decoder(16#7b#)) OR
 					(reg_q397 AND symb_decoder(16#ee#)) OR
 					(reg_q397 AND symb_decoder(16#fa#)) OR
 					(reg_q397 AND symb_decoder(16#16#)) OR
 					(reg_q397 AND symb_decoder(16#43#)) OR
 					(reg_q397 AND symb_decoder(16#e8#)) OR
 					(reg_q397 AND symb_decoder(16#37#)) OR
 					(reg_q397 AND symb_decoder(16#32#)) OR
 					(reg_q397 AND symb_decoder(16#53#)) OR
 					(reg_q397 AND symb_decoder(16#88#));
reg_q540_in <= (reg_q526 AND symb_decoder(16#69#)) OR
 					(reg_q526 AND symb_decoder(16#04#)) OR
 					(reg_q526 AND symb_decoder(16#b3#)) OR
 					(reg_q526 AND symb_decoder(16#60#)) OR
 					(reg_q526 AND symb_decoder(16#a2#)) OR
 					(reg_q526 AND symb_decoder(16#d3#)) OR
 					(reg_q526 AND symb_decoder(16#21#)) OR
 					(reg_q526 AND symb_decoder(16#d0#)) OR
 					(reg_q526 AND symb_decoder(16#7e#)) OR
 					(reg_q526 AND symb_decoder(16#0b#)) OR
 					(reg_q526 AND symb_decoder(16#b0#)) OR
 					(reg_q526 AND symb_decoder(16#31#)) OR
 					(reg_q526 AND symb_decoder(16#b4#)) OR
 					(reg_q526 AND symb_decoder(16#9a#)) OR
 					(reg_q526 AND symb_decoder(16#09#)) OR
 					(reg_q526 AND symb_decoder(16#64#)) OR
 					(reg_q526 AND symb_decoder(16#db#)) OR
 					(reg_q526 AND symb_decoder(16#f8#)) OR
 					(reg_q526 AND symb_decoder(16#f4#)) OR
 					(reg_q526 AND symb_decoder(16#89#)) OR
 					(reg_q526 AND symb_decoder(16#6b#)) OR
 					(reg_q526 AND symb_decoder(16#ad#)) OR
 					(reg_q526 AND symb_decoder(16#9c#)) OR
 					(reg_q526 AND symb_decoder(16#a4#)) OR
 					(reg_q526 AND symb_decoder(16#aa#)) OR
 					(reg_q526 AND symb_decoder(16#61#)) OR
 					(reg_q526 AND symb_decoder(16#7d#)) OR
 					(reg_q526 AND symb_decoder(16#47#)) OR
 					(reg_q526 AND symb_decoder(16#4a#)) OR
 					(reg_q526 AND symb_decoder(16#3b#)) OR
 					(reg_q526 AND symb_decoder(16#ec#)) OR
 					(reg_q526 AND symb_decoder(16#19#)) OR
 					(reg_q526 AND symb_decoder(16#ed#)) OR
 					(reg_q526 AND symb_decoder(16#f7#)) OR
 					(reg_q526 AND symb_decoder(16#eb#)) OR
 					(reg_q526 AND symb_decoder(16#e8#)) OR
 					(reg_q526 AND symb_decoder(16#fd#)) OR
 					(reg_q526 AND symb_decoder(16#9b#)) OR
 					(reg_q526 AND symb_decoder(16#29#)) OR
 					(reg_q526 AND symb_decoder(16#39#)) OR
 					(reg_q526 AND symb_decoder(16#a6#)) OR
 					(reg_q526 AND symb_decoder(16#18#)) OR
 					(reg_q526 AND symb_decoder(16#25#)) OR
 					(reg_q526 AND symb_decoder(16#5c#)) OR
 					(reg_q526 AND symb_decoder(16#d9#)) OR
 					(reg_q526 AND symb_decoder(16#bd#)) OR
 					(reg_q526 AND symb_decoder(16#02#)) OR
 					(reg_q526 AND symb_decoder(16#f2#)) OR
 					(reg_q526 AND symb_decoder(16#e6#)) OR
 					(reg_q526 AND symb_decoder(16#44#)) OR
 					(reg_q526 AND symb_decoder(16#da#)) OR
 					(reg_q526 AND symb_decoder(16#3d#)) OR
 					(reg_q526 AND symb_decoder(16#07#)) OR
 					(reg_q526 AND symb_decoder(16#d1#)) OR
 					(reg_q526 AND symb_decoder(16#16#)) OR
 					(reg_q526 AND symb_decoder(16#77#)) OR
 					(reg_q526 AND symb_decoder(16#2c#)) OR
 					(reg_q526 AND symb_decoder(16#c6#)) OR
 					(reg_q526 AND symb_decoder(16#f6#)) OR
 					(reg_q526 AND symb_decoder(16#56#)) OR
 					(reg_q526 AND symb_decoder(16#0c#)) OR
 					(reg_q526 AND symb_decoder(16#5f#)) OR
 					(reg_q526 AND symb_decoder(16#ff#)) OR
 					(reg_q526 AND symb_decoder(16#e0#)) OR
 					(reg_q526 AND symb_decoder(16#4f#)) OR
 					(reg_q526 AND symb_decoder(16#10#)) OR
 					(reg_q526 AND symb_decoder(16#58#)) OR
 					(reg_q526 AND symb_decoder(16#f9#)) OR
 					(reg_q526 AND symb_decoder(16#75#)) OR
 					(reg_q526 AND symb_decoder(16#11#)) OR
 					(reg_q526 AND symb_decoder(16#fa#)) OR
 					(reg_q526 AND symb_decoder(16#98#)) OR
 					(reg_q526 AND symb_decoder(16#af#)) OR
 					(reg_q526 AND symb_decoder(16#2f#)) OR
 					(reg_q526 AND symb_decoder(16#a1#)) OR
 					(reg_q526 AND symb_decoder(16#12#)) OR
 					(reg_q526 AND symb_decoder(16#4e#)) OR
 					(reg_q526 AND symb_decoder(16#7f#)) OR
 					(reg_q526 AND symb_decoder(16#6a#)) OR
 					(reg_q526 AND symb_decoder(16#8e#)) OR
 					(reg_q526 AND symb_decoder(16#13#)) OR
 					(reg_q526 AND symb_decoder(16#95#)) OR
 					(reg_q526 AND symb_decoder(16#e2#)) OR
 					(reg_q526 AND symb_decoder(16#f1#)) OR
 					(reg_q526 AND symb_decoder(16#32#)) OR
 					(reg_q526 AND symb_decoder(16#a0#)) OR
 					(reg_q526 AND symb_decoder(16#6c#)) OR
 					(reg_q526 AND symb_decoder(16#22#)) OR
 					(reg_q526 AND symb_decoder(16#08#)) OR
 					(reg_q526 AND symb_decoder(16#0e#)) OR
 					(reg_q526 AND symb_decoder(16#70#)) OR
 					(reg_q526 AND symb_decoder(16#1d#)) OR
 					(reg_q526 AND symb_decoder(16#91#)) OR
 					(reg_q526 AND symb_decoder(16#1b#)) OR
 					(reg_q526 AND symb_decoder(16#59#)) OR
 					(reg_q526 AND symb_decoder(16#63#)) OR
 					(reg_q526 AND symb_decoder(16#ca#)) OR
 					(reg_q526 AND symb_decoder(16#7c#)) OR
 					(reg_q526 AND symb_decoder(16#38#)) OR
 					(reg_q526 AND symb_decoder(16#66#)) OR
 					(reg_q526 AND symb_decoder(16#93#)) OR
 					(reg_q526 AND symb_decoder(16#54#)) OR
 					(reg_q526 AND symb_decoder(16#b9#)) OR
 					(reg_q526 AND symb_decoder(16#73#)) OR
 					(reg_q526 AND symb_decoder(16#00#)) OR
 					(reg_q526 AND symb_decoder(16#f0#)) OR
 					(reg_q526 AND symb_decoder(16#ba#)) OR
 					(reg_q526 AND symb_decoder(16#8d#)) OR
 					(reg_q526 AND symb_decoder(16#c0#)) OR
 					(reg_q526 AND symb_decoder(16#2b#)) OR
 					(reg_q526 AND symb_decoder(16#e5#)) OR
 					(reg_q526 AND symb_decoder(16#bc#)) OR
 					(reg_q526 AND symb_decoder(16#0f#)) OR
 					(reg_q526 AND symb_decoder(16#c5#)) OR
 					(reg_q526 AND symb_decoder(16#d2#)) OR
 					(reg_q526 AND symb_decoder(16#43#)) OR
 					(reg_q526 AND symb_decoder(16#2d#)) OR
 					(reg_q526 AND symb_decoder(16#ea#)) OR
 					(reg_q526 AND symb_decoder(16#28#)) OR
 					(reg_q526 AND symb_decoder(16#99#)) OR
 					(reg_q526 AND symb_decoder(16#20#)) OR
 					(reg_q526 AND symb_decoder(16#7a#)) OR
 					(reg_q526 AND symb_decoder(16#1a#)) OR
 					(reg_q526 AND symb_decoder(16#2a#)) OR
 					(reg_q526 AND symb_decoder(16#45#)) OR
 					(reg_q526 AND symb_decoder(16#fc#)) OR
 					(reg_q526 AND symb_decoder(16#79#)) OR
 					(reg_q526 AND symb_decoder(16#4d#)) OR
 					(reg_q526 AND symb_decoder(16#9e#)) OR
 					(reg_q526 AND symb_decoder(16#46#)) OR
 					(reg_q526 AND symb_decoder(16#cd#)) OR
 					(reg_q526 AND symb_decoder(16#cf#)) OR
 					(reg_q526 AND symb_decoder(16#97#)) OR
 					(reg_q526 AND symb_decoder(16#9f#)) OR
 					(reg_q526 AND symb_decoder(16#42#)) OR
 					(reg_q526 AND symb_decoder(16#be#)) OR
 					(reg_q526 AND symb_decoder(16#84#)) OR
 					(reg_q526 AND symb_decoder(16#b2#)) OR
 					(reg_q526 AND symb_decoder(16#83#)) OR
 					(reg_q526 AND symb_decoder(16#37#)) OR
 					(reg_q526 AND symb_decoder(16#94#)) OR
 					(reg_q526 AND symb_decoder(16#d5#)) OR
 					(reg_q526 AND symb_decoder(16#03#)) OR
 					(reg_q526 AND symb_decoder(16#87#)) OR
 					(reg_q526 AND symb_decoder(16#27#)) OR
 					(reg_q526 AND symb_decoder(16#8c#)) OR
 					(reg_q526 AND symb_decoder(16#41#)) OR
 					(reg_q526 AND symb_decoder(16#48#)) OR
 					(reg_q526 AND symb_decoder(16#bf#)) OR
 					(reg_q526 AND symb_decoder(16#78#)) OR
 					(reg_q526 AND symb_decoder(16#8f#)) OR
 					(reg_q526 AND symb_decoder(16#35#)) OR
 					(reg_q526 AND symb_decoder(16#74#)) OR
 					(reg_q526 AND symb_decoder(16#34#)) OR
 					(reg_q526 AND symb_decoder(16#49#)) OR
 					(reg_q526 AND symb_decoder(16#01#)) OR
 					(reg_q526 AND symb_decoder(16#15#)) OR
 					(reg_q526 AND symb_decoder(16#d6#)) OR
 					(reg_q526 AND symb_decoder(16#81#)) OR
 					(reg_q526 AND symb_decoder(16#92#)) OR
 					(reg_q526 AND symb_decoder(16#72#)) OR
 					(reg_q526 AND symb_decoder(16#1c#)) OR
 					(reg_q526 AND symb_decoder(16#a9#)) OR
 					(reg_q526 AND symb_decoder(16#67#)) OR
 					(reg_q526 AND symb_decoder(16#3f#)) OR
 					(reg_q526 AND symb_decoder(16#b6#)) OR
 					(reg_q526 AND symb_decoder(16#c4#)) OR
 					(reg_q526 AND symb_decoder(16#b7#)) OR
 					(reg_q526 AND symb_decoder(16#8a#)) OR
 					(reg_q526 AND symb_decoder(16#e1#)) OR
 					(reg_q526 AND symb_decoder(16#ce#)) OR
 					(reg_q526 AND symb_decoder(16#c8#)) OR
 					(reg_q526 AND symb_decoder(16#24#)) OR
 					(reg_q526 AND symb_decoder(16#ae#)) OR
 					(reg_q526 AND symb_decoder(16#8b#)) OR
 					(reg_q526 AND symb_decoder(16#5e#)) OR
 					(reg_q526 AND symb_decoder(16#f3#)) OR
 					(reg_q526 AND symb_decoder(16#14#)) OR
 					(reg_q526 AND symb_decoder(16#dc#)) OR
 					(reg_q526 AND symb_decoder(16#fe#)) OR
 					(reg_q526 AND symb_decoder(16#1e#)) OR
 					(reg_q526 AND symb_decoder(16#a3#)) OR
 					(reg_q526 AND symb_decoder(16#ac#)) OR
 					(reg_q526 AND symb_decoder(16#6e#)) OR
 					(reg_q526 AND symb_decoder(16#ab#)) OR
 					(reg_q526 AND symb_decoder(16#c2#)) OR
 					(reg_q526 AND symb_decoder(16#96#)) OR
 					(reg_q526 AND symb_decoder(16#4b#)) OR
 					(reg_q526 AND symb_decoder(16#2e#)) OR
 					(reg_q526 AND symb_decoder(16#26#)) OR
 					(reg_q526 AND symb_decoder(16#d4#)) OR
 					(reg_q526 AND symb_decoder(16#a7#)) OR
 					(reg_q526 AND symb_decoder(16#05#)) OR
 					(reg_q526 AND symb_decoder(16#dd#)) OR
 					(reg_q526 AND symb_decoder(16#e4#)) OR
 					(reg_q526 AND symb_decoder(16#ee#)) OR
 					(reg_q526 AND symb_decoder(16#b8#)) OR
 					(reg_q526 AND symb_decoder(16#88#)) OR
 					(reg_q526 AND symb_decoder(16#cc#)) OR
 					(reg_q526 AND symb_decoder(16#4c#)) OR
 					(reg_q526 AND symb_decoder(16#d8#)) OR
 					(reg_q526 AND symb_decoder(16#cb#)) OR
 					(reg_q526 AND symb_decoder(16#e9#)) OR
 					(reg_q526 AND symb_decoder(16#52#)) OR
 					(reg_q526 AND symb_decoder(16#ef#)) OR
 					(reg_q526 AND symb_decoder(16#17#)) OR
 					(reg_q526 AND symb_decoder(16#85#)) OR
 					(reg_q526 AND symb_decoder(16#df#)) OR
 					(reg_q526 AND symb_decoder(16#de#)) OR
 					(reg_q526 AND symb_decoder(16#33#)) OR
 					(reg_q526 AND symb_decoder(16#b5#)) OR
 					(reg_q526 AND symb_decoder(16#c9#)) OR
 					(reg_q526 AND symb_decoder(16#1f#)) OR
 					(reg_q526 AND symb_decoder(16#e7#)) OR
 					(reg_q526 AND symb_decoder(16#50#)) OR
 					(reg_q526 AND symb_decoder(16#b1#)) OR
 					(reg_q526 AND symb_decoder(16#c3#)) OR
 					(reg_q526 AND symb_decoder(16#5d#)) OR
 					(reg_q526 AND symb_decoder(16#3c#)) OR
 					(reg_q526 AND symb_decoder(16#51#)) OR
 					(reg_q526 AND symb_decoder(16#f5#)) OR
 					(reg_q526 AND symb_decoder(16#82#)) OR
 					(reg_q526 AND symb_decoder(16#80#)) OR
 					(reg_q526 AND symb_decoder(16#36#)) OR
 					(reg_q526 AND symb_decoder(16#86#)) OR
 					(reg_q526 AND symb_decoder(16#6d#)) OR
 					(reg_q526 AND symb_decoder(16#76#)) OR
 					(reg_q526 AND symb_decoder(16#90#)) OR
 					(reg_q526 AND symb_decoder(16#6f#)) OR
 					(reg_q526 AND symb_decoder(16#fb#)) OR
 					(reg_q526 AND symb_decoder(16#65#)) OR
 					(reg_q526 AND symb_decoder(16#62#)) OR
 					(reg_q526 AND symb_decoder(16#23#)) OR
 					(reg_q526 AND symb_decoder(16#68#)) OR
 					(reg_q526 AND symb_decoder(16#55#)) OR
 					(reg_q526 AND symb_decoder(16#c1#)) OR
 					(reg_q526 AND symb_decoder(16#53#)) OR
 					(reg_q526 AND symb_decoder(16#71#)) OR
 					(reg_q526 AND symb_decoder(16#06#)) OR
 					(reg_q526 AND symb_decoder(16#40#)) OR
 					(reg_q526 AND symb_decoder(16#3a#)) OR
 					(reg_q526 AND symb_decoder(16#9d#)) OR
 					(reg_q526 AND symb_decoder(16#5a#)) OR
 					(reg_q526 AND symb_decoder(16#a5#)) OR
 					(reg_q526 AND symb_decoder(16#c7#)) OR
 					(reg_q526 AND symb_decoder(16#d7#)) OR
 					(reg_q526 AND symb_decoder(16#30#)) OR
 					(reg_q526 AND symb_decoder(16#7b#)) OR
 					(reg_q526 AND symb_decoder(16#5b#)) OR
 					(reg_q526 AND symb_decoder(16#e3#)) OR
 					(reg_q526 AND symb_decoder(16#57#)) OR
 					(reg_q526 AND symb_decoder(16#3e#)) OR
 					(reg_q526 AND symb_decoder(16#a8#)) OR
 					(reg_q526 AND symb_decoder(16#bb#)) OR
 					(reg_q540 AND symb_decoder(16#d6#)) OR
 					(reg_q540 AND symb_decoder(16#1b#)) OR
 					(reg_q540 AND symb_decoder(16#c5#)) OR
 					(reg_q540 AND symb_decoder(16#5a#)) OR
 					(reg_q540 AND symb_decoder(16#0b#)) OR
 					(reg_q540 AND symb_decoder(16#56#)) OR
 					(reg_q540 AND symb_decoder(16#a6#)) OR
 					(reg_q540 AND symb_decoder(16#99#)) OR
 					(reg_q540 AND symb_decoder(16#d3#)) OR
 					(reg_q540 AND symb_decoder(16#6b#)) OR
 					(reg_q540 AND symb_decoder(16#ed#)) OR
 					(reg_q540 AND symb_decoder(16#8d#)) OR
 					(reg_q540 AND symb_decoder(16#e2#)) OR
 					(reg_q540 AND symb_decoder(16#55#)) OR
 					(reg_q540 AND symb_decoder(16#78#)) OR
 					(reg_q540 AND symb_decoder(16#6e#)) OR
 					(reg_q540 AND symb_decoder(16#90#)) OR
 					(reg_q540 AND symb_decoder(16#b2#)) OR
 					(reg_q540 AND symb_decoder(16#21#)) OR
 					(reg_q540 AND symb_decoder(16#19#)) OR
 					(reg_q540 AND symb_decoder(16#d9#)) OR
 					(reg_q540 AND symb_decoder(16#61#)) OR
 					(reg_q540 AND symb_decoder(16#0e#)) OR
 					(reg_q540 AND symb_decoder(16#b5#)) OR
 					(reg_q540 AND symb_decoder(16#12#)) OR
 					(reg_q540 AND symb_decoder(16#a9#)) OR
 					(reg_q540 AND symb_decoder(16#25#)) OR
 					(reg_q540 AND symb_decoder(16#e1#)) OR
 					(reg_q540 AND symb_decoder(16#52#)) OR
 					(reg_q540 AND symb_decoder(16#ac#)) OR
 					(reg_q540 AND symb_decoder(16#f7#)) OR
 					(reg_q540 AND symb_decoder(16#35#)) OR
 					(reg_q540 AND symb_decoder(16#0f#)) OR
 					(reg_q540 AND symb_decoder(16#26#)) OR
 					(reg_q540 AND symb_decoder(16#29#)) OR
 					(reg_q540 AND symb_decoder(16#5f#)) OR
 					(reg_q540 AND symb_decoder(16#5d#)) OR
 					(reg_q540 AND symb_decoder(16#ea#)) OR
 					(reg_q540 AND symb_decoder(16#41#)) OR
 					(reg_q540 AND symb_decoder(16#a2#)) OR
 					(reg_q540 AND symb_decoder(16#97#)) OR
 					(reg_q540 AND symb_decoder(16#bf#)) OR
 					(reg_q540 AND symb_decoder(16#f2#)) OR
 					(reg_q540 AND symb_decoder(16#8f#)) OR
 					(reg_q540 AND symb_decoder(16#49#)) OR
 					(reg_q540 AND symb_decoder(16#f5#)) OR
 					(reg_q540 AND symb_decoder(16#e8#)) OR
 					(reg_q540 AND symb_decoder(16#37#)) OR
 					(reg_q540 AND symb_decoder(16#c0#)) OR
 					(reg_q540 AND symb_decoder(16#bb#)) OR
 					(reg_q540 AND symb_decoder(16#18#)) OR
 					(reg_q540 AND symb_decoder(16#5c#)) OR
 					(reg_q540 AND symb_decoder(16#d5#)) OR
 					(reg_q540 AND symb_decoder(16#9e#)) OR
 					(reg_q540 AND symb_decoder(16#66#)) OR
 					(reg_q540 AND symb_decoder(16#87#)) OR
 					(reg_q540 AND symb_decoder(16#1e#)) OR
 					(reg_q540 AND symb_decoder(16#28#)) OR
 					(reg_q540 AND symb_decoder(16#1c#)) OR
 					(reg_q540 AND symb_decoder(16#93#)) OR
 					(reg_q540 AND symb_decoder(16#77#)) OR
 					(reg_q540 AND symb_decoder(16#05#)) OR
 					(reg_q540 AND symb_decoder(16#ca#)) OR
 					(reg_q540 AND symb_decoder(16#53#)) OR
 					(reg_q540 AND symb_decoder(16#64#)) OR
 					(reg_q540 AND symb_decoder(16#16#)) OR
 					(reg_q540 AND symb_decoder(16#96#)) OR
 					(reg_q540 AND symb_decoder(16#13#)) OR
 					(reg_q540 AND symb_decoder(16#24#)) OR
 					(reg_q540 AND symb_decoder(16#15#)) OR
 					(reg_q540 AND symb_decoder(16#ff#)) OR
 					(reg_q540 AND symb_decoder(16#cf#)) OR
 					(reg_q540 AND symb_decoder(16#c6#)) OR
 					(reg_q540 AND symb_decoder(16#68#)) OR
 					(reg_q540 AND symb_decoder(16#b8#)) OR
 					(reg_q540 AND symb_decoder(16#9b#)) OR
 					(reg_q540 AND symb_decoder(16#e0#)) OR
 					(reg_q540 AND symb_decoder(16#7a#)) OR
 					(reg_q540 AND symb_decoder(16#f9#)) OR
 					(reg_q540 AND symb_decoder(16#07#)) OR
 					(reg_q540 AND symb_decoder(16#6d#)) OR
 					(reg_q540 AND symb_decoder(16#50#)) OR
 					(reg_q540 AND symb_decoder(16#69#)) OR
 					(reg_q540 AND symb_decoder(16#9c#)) OR
 					(reg_q540 AND symb_decoder(16#74#)) OR
 					(reg_q540 AND symb_decoder(16#02#)) OR
 					(reg_q540 AND symb_decoder(16#b3#)) OR
 					(reg_q540 AND symb_decoder(16#14#)) OR
 					(reg_q540 AND symb_decoder(16#57#)) OR
 					(reg_q540 AND symb_decoder(16#a5#)) OR
 					(reg_q540 AND symb_decoder(16#e7#)) OR
 					(reg_q540 AND symb_decoder(16#d8#)) OR
 					(reg_q540 AND symb_decoder(16#ab#)) OR
 					(reg_q540 AND symb_decoder(16#09#)) OR
 					(reg_q540 AND symb_decoder(16#fd#)) OR
 					(reg_q540 AND symb_decoder(16#3a#)) OR
 					(reg_q540 AND symb_decoder(16#08#)) OR
 					(reg_q540 AND symb_decoder(16#e3#)) OR
 					(reg_q540 AND symb_decoder(16#76#)) OR
 					(reg_q540 AND symb_decoder(16#e6#)) OR
 					(reg_q540 AND symb_decoder(16#23#)) OR
 					(reg_q540 AND symb_decoder(16#63#)) OR
 					(reg_q540 AND symb_decoder(16#f1#)) OR
 					(reg_q540 AND symb_decoder(16#59#)) OR
 					(reg_q540 AND symb_decoder(16#de#)) OR
 					(reg_q540 AND symb_decoder(16#3b#)) OR
 					(reg_q540 AND symb_decoder(16#5e#)) OR
 					(reg_q540 AND symb_decoder(16#22#)) OR
 					(reg_q540 AND symb_decoder(16#30#)) OR
 					(reg_q540 AND symb_decoder(16#bc#)) OR
 					(reg_q540 AND symb_decoder(16#8e#)) OR
 					(reg_q540 AND symb_decoder(16#94#)) OR
 					(reg_q540 AND symb_decoder(16#60#)) OR
 					(reg_q540 AND symb_decoder(16#2e#)) OR
 					(reg_q540 AND symb_decoder(16#a7#)) OR
 					(reg_q540 AND symb_decoder(16#42#)) OR
 					(reg_q540 AND symb_decoder(16#b6#)) OR
 					(reg_q540 AND symb_decoder(16#95#)) OR
 					(reg_q540 AND symb_decoder(16#ec#)) OR
 					(reg_q540 AND symb_decoder(16#1f#)) OR
 					(reg_q540 AND symb_decoder(16#d1#)) OR
 					(reg_q540 AND symb_decoder(16#39#)) OR
 					(reg_q540 AND symb_decoder(16#33#)) OR
 					(reg_q540 AND symb_decoder(16#3d#)) OR
 					(reg_q540 AND symb_decoder(16#04#)) OR
 					(reg_q540 AND symb_decoder(16#40#)) OR
 					(reg_q540 AND symb_decoder(16#f4#)) OR
 					(reg_q540 AND symb_decoder(16#e5#)) OR
 					(reg_q540 AND symb_decoder(16#5b#)) OR
 					(reg_q540 AND symb_decoder(16#8c#)) OR
 					(reg_q540 AND symb_decoder(16#54#)) OR
 					(reg_q540 AND symb_decoder(16#17#)) OR
 					(reg_q540 AND symb_decoder(16#be#)) OR
 					(reg_q540 AND symb_decoder(16#65#)) OR
 					(reg_q540 AND symb_decoder(16#d4#)) OR
 					(reg_q540 AND symb_decoder(16#cd#)) OR
 					(reg_q540 AND symb_decoder(16#4d#)) OR
 					(reg_q540 AND symb_decoder(16#f0#)) OR
 					(reg_q540 AND symb_decoder(16#aa#)) OR
 					(reg_q540 AND symb_decoder(16#0c#)) OR
 					(reg_q540 AND symb_decoder(16#06#)) OR
 					(reg_q540 AND symb_decoder(16#c1#)) OR
 					(reg_q540 AND symb_decoder(16#cb#)) OR
 					(reg_q540 AND symb_decoder(16#1d#)) OR
 					(reg_q540 AND symb_decoder(16#eb#)) OR
 					(reg_q540 AND symb_decoder(16#4e#)) OR
 					(reg_q540 AND symb_decoder(16#9f#)) OR
 					(reg_q540 AND symb_decoder(16#d0#)) OR
 					(reg_q540 AND symb_decoder(16#1a#)) OR
 					(reg_q540 AND symb_decoder(16#4a#)) OR
 					(reg_q540 AND symb_decoder(16#7c#)) OR
 					(reg_q540 AND symb_decoder(16#a4#)) OR
 					(reg_q540 AND symb_decoder(16#48#)) OR
 					(reg_q540 AND symb_decoder(16#af#)) OR
 					(reg_q540 AND symb_decoder(16#fc#)) OR
 					(reg_q540 AND symb_decoder(16#a8#)) OR
 					(reg_q540 AND symb_decoder(16#9d#)) OR
 					(reg_q540 AND symb_decoder(16#d2#)) OR
 					(reg_q540 AND symb_decoder(16#2b#)) OR
 					(reg_q540 AND symb_decoder(16#d7#)) OR
 					(reg_q540 AND symb_decoder(16#34#)) OR
 					(reg_q540 AND symb_decoder(16#85#)) OR
 					(reg_q540 AND symb_decoder(16#70#)) OR
 					(reg_q540 AND symb_decoder(16#62#)) OR
 					(reg_q540 AND symb_decoder(16#b7#)) OR
 					(reg_q540 AND symb_decoder(16#f8#)) OR
 					(reg_q540 AND symb_decoder(16#8a#)) OR
 					(reg_q540 AND symb_decoder(16#27#)) OR
 					(reg_q540 AND symb_decoder(16#58#)) OR
 					(reg_q540 AND symb_decoder(16#bd#)) OR
 					(reg_q540 AND symb_decoder(16#ad#)) OR
 					(reg_q540 AND symb_decoder(16#7d#)) OR
 					(reg_q540 AND symb_decoder(16#31#)) OR
 					(reg_q540 AND symb_decoder(16#8b#)) OR
 					(reg_q540 AND symb_decoder(16#c3#)) OR
 					(reg_q540 AND symb_decoder(16#c4#)) OR
 					(reg_q540 AND symb_decoder(16#6a#)) OR
 					(reg_q540 AND symb_decoder(16#92#)) OR
 					(reg_q540 AND symb_decoder(16#67#)) OR
 					(reg_q540 AND symb_decoder(16#88#)) OR
 					(reg_q540 AND symb_decoder(16#43#)) OR
 					(reg_q540 AND symb_decoder(16#b0#)) OR
 					(reg_q540 AND symb_decoder(16#11#)) OR
 					(reg_q540 AND symb_decoder(16#b4#)) OR
 					(reg_q540 AND symb_decoder(16#e4#)) OR
 					(reg_q540 AND symb_decoder(16#32#)) OR
 					(reg_q540 AND symb_decoder(16#ee#)) OR
 					(reg_q540 AND symb_decoder(16#86#)) OR
 					(reg_q540 AND symb_decoder(16#ef#)) OR
 					(reg_q540 AND symb_decoder(16#44#)) OR
 					(reg_q540 AND symb_decoder(16#79#)) OR
 					(reg_q540 AND symb_decoder(16#4b#)) OR
 					(reg_q540 AND symb_decoder(16#ae#)) OR
 					(reg_q540 AND symb_decoder(16#2c#)) OR
 					(reg_q540 AND symb_decoder(16#01#)) OR
 					(reg_q540 AND symb_decoder(16#da#)) OR
 					(reg_q540 AND symb_decoder(16#3f#)) OR
 					(reg_q540 AND symb_decoder(16#4f#)) OR
 					(reg_q540 AND symb_decoder(16#6c#)) OR
 					(reg_q540 AND symb_decoder(16#2f#)) OR
 					(reg_q540 AND symb_decoder(16#db#)) OR
 					(reg_q540 AND symb_decoder(16#b1#)) OR
 					(reg_q540 AND symb_decoder(16#ce#)) OR
 					(reg_q540 AND symb_decoder(16#b9#)) OR
 					(reg_q540 AND symb_decoder(16#f3#)) OR
 					(reg_q540 AND symb_decoder(16#4c#)) OR
 					(reg_q540 AND symb_decoder(16#dd#)) OR
 					(reg_q540 AND symb_decoder(16#7f#)) OR
 					(reg_q540 AND symb_decoder(16#df#)) OR
 					(reg_q540 AND symb_decoder(16#36#)) OR
 					(reg_q540 AND symb_decoder(16#c9#)) OR
 					(reg_q540 AND symb_decoder(16#82#)) OR
 					(reg_q540 AND symb_decoder(16#83#)) OR
 					(reg_q540 AND symb_decoder(16#dc#)) OR
 					(reg_q540 AND symb_decoder(16#c7#)) OR
 					(reg_q540 AND symb_decoder(16#fe#)) OR
 					(reg_q540 AND symb_decoder(16#fa#)) OR
 					(reg_q540 AND symb_decoder(16#e9#)) OR
 					(reg_q540 AND symb_decoder(16#c2#)) OR
 					(reg_q540 AND symb_decoder(16#72#)) OR
 					(reg_q540 AND symb_decoder(16#f6#)) OR
 					(reg_q540 AND symb_decoder(16#75#)) OR
 					(reg_q540 AND symb_decoder(16#80#)) OR
 					(reg_q540 AND symb_decoder(16#45#)) OR
 					(reg_q540 AND symb_decoder(16#a1#)) OR
 					(reg_q540 AND symb_decoder(16#6f#)) OR
 					(reg_q540 AND symb_decoder(16#3e#)) OR
 					(reg_q540 AND symb_decoder(16#71#)) OR
 					(reg_q540 AND symb_decoder(16#89#)) OR
 					(reg_q540 AND symb_decoder(16#81#)) OR
 					(reg_q540 AND symb_decoder(16#c8#)) OR
 					(reg_q540 AND symb_decoder(16#3c#)) OR
 					(reg_q540 AND symb_decoder(16#20#)) OR
 					(reg_q540 AND symb_decoder(16#47#)) OR
 					(reg_q540 AND symb_decoder(16#73#)) OR
 					(reg_q540 AND symb_decoder(16#7e#)) OR
 					(reg_q540 AND symb_decoder(16#84#)) OR
 					(reg_q540 AND symb_decoder(16#7b#)) OR
 					(reg_q540 AND symb_decoder(16#a3#)) OR
 					(reg_q540 AND symb_decoder(16#a0#)) OR
 					(reg_q540 AND symb_decoder(16#46#)) OR
 					(reg_q540 AND symb_decoder(16#10#)) OR
 					(reg_q540 AND symb_decoder(16#51#)) OR
 					(reg_q540 AND symb_decoder(16#03#)) OR
 					(reg_q540 AND symb_decoder(16#fb#)) OR
 					(reg_q540 AND symb_decoder(16#98#)) OR
 					(reg_q540 AND symb_decoder(16#00#)) OR
 					(reg_q540 AND symb_decoder(16#9a#)) OR
 					(reg_q540 AND symb_decoder(16#ba#)) OR
 					(reg_q540 AND symb_decoder(16#91#)) OR
 					(reg_q540 AND symb_decoder(16#cc#)) OR
 					(reg_q540 AND symb_decoder(16#2a#)) OR
 					(reg_q540 AND symb_decoder(16#2d#)) OR
 					(reg_q540 AND symb_decoder(16#38#));
reg_q847_in <= (reg_q847 AND symb_decoder(16#35#)) OR
 					(reg_q847 AND symb_decoder(16#32#)) OR
 					(reg_q847 AND symb_decoder(16#31#)) OR
 					(reg_q847 AND symb_decoder(16#38#)) OR
 					(reg_q847 AND symb_decoder(16#33#)) OR
 					(reg_q847 AND symb_decoder(16#30#)) OR
 					(reg_q847 AND symb_decoder(16#37#)) OR
 					(reg_q847 AND symb_decoder(16#36#)) OR
 					(reg_q847 AND symb_decoder(16#34#)) OR
 					(reg_q847 AND symb_decoder(16#39#)) OR
 					(reg_q845 AND symb_decoder(16#33#)) OR
 					(reg_q845 AND symb_decoder(16#30#)) OR
 					(reg_q845 AND symb_decoder(16#37#)) OR
 					(reg_q845 AND symb_decoder(16#31#)) OR
 					(reg_q845 AND symb_decoder(16#36#)) OR
 					(reg_q845 AND symb_decoder(16#39#)) OR
 					(reg_q845 AND symb_decoder(16#34#)) OR
 					(reg_q845 AND symb_decoder(16#35#)) OR
 					(reg_q845 AND symb_decoder(16#32#)) OR
 					(reg_q845 AND symb_decoder(16#38#));
reg_q855_in <= (reg_q855 AND symb_decoder(16#39#)) OR
 					(reg_q855 AND symb_decoder(16#33#)) OR
 					(reg_q855 AND symb_decoder(16#31#)) OR
 					(reg_q855 AND symb_decoder(16#37#)) OR
 					(reg_q855 AND symb_decoder(16#38#)) OR
 					(reg_q855 AND symb_decoder(16#34#)) OR
 					(reg_q855 AND symb_decoder(16#30#)) OR
 					(reg_q855 AND symb_decoder(16#35#)) OR
 					(reg_q855 AND symb_decoder(16#36#)) OR
 					(reg_q855 AND symb_decoder(16#32#)) OR
 					(reg_q853 AND symb_decoder(16#39#)) OR
 					(reg_q853 AND symb_decoder(16#38#)) OR
 					(reg_q853 AND symb_decoder(16#35#)) OR
 					(reg_q853 AND symb_decoder(16#37#)) OR
 					(reg_q853 AND symb_decoder(16#32#)) OR
 					(reg_q853 AND symb_decoder(16#33#)) OR
 					(reg_q853 AND symb_decoder(16#36#)) OR
 					(reg_q853 AND symb_decoder(16#31#)) OR
 					(reg_q853 AND symb_decoder(16#30#)) OR
 					(reg_q853 AND symb_decoder(16#34#));
reg_q823_in <= (reg_q819 AND symb_decoder(16#69#)) OR
 					(reg_q819 AND symb_decoder(16#49#)) OR
 					(reg_q857 AND symb_decoder(16#69#)) OR
 					(reg_q857 AND symb_decoder(16#49#));
reg_q853_in <= (reg_q851 AND symb_decoder(16#2e#));
reg_q845_in <= (reg_q843 AND symb_decoder(16#2e#));
reg_q843_in <= (reg_q841 AND symb_decoder(16#30#)) OR
 					(reg_q841 AND symb_decoder(16#31#)) OR
 					(reg_q841 AND symb_decoder(16#38#)) OR
 					(reg_q841 AND symb_decoder(16#34#)) OR
 					(reg_q841 AND symb_decoder(16#33#)) OR
 					(reg_q841 AND symb_decoder(16#39#)) OR
 					(reg_q841 AND symb_decoder(16#37#)) OR
 					(reg_q841 AND symb_decoder(16#32#)) OR
 					(reg_q841 AND symb_decoder(16#35#)) OR
 					(reg_q841 AND symb_decoder(16#36#)) OR
 					(reg_q843 AND symb_decoder(16#34#)) OR
 					(reg_q843 AND symb_decoder(16#31#)) OR
 					(reg_q843 AND symb_decoder(16#37#)) OR
 					(reg_q843 AND symb_decoder(16#38#)) OR
 					(reg_q843 AND symb_decoder(16#30#)) OR
 					(reg_q843 AND symb_decoder(16#36#)) OR
 					(reg_q843 AND symb_decoder(16#32#)) OR
 					(reg_q843 AND symb_decoder(16#39#)) OR
 					(reg_q843 AND symb_decoder(16#35#)) OR
 					(reg_q843 AND symb_decoder(16#33#));
reg_q1146_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q1145 AND symb_decoder(16#0a#)) OR
 					(reg_q1145 AND symb_decoder(16#0d#));
reg_q849_in <= (reg_q847 AND symb_decoder(16#2e#));
reg_q851_in <= (reg_q849 AND symb_decoder(16#35#)) OR
 					(reg_q849 AND symb_decoder(16#37#)) OR
 					(reg_q849 AND symb_decoder(16#39#)) OR
 					(reg_q849 AND symb_decoder(16#38#)) OR
 					(reg_q849 AND symb_decoder(16#34#)) OR
 					(reg_q849 AND symb_decoder(16#30#)) OR
 					(reg_q849 AND symb_decoder(16#31#)) OR
 					(reg_q849 AND symb_decoder(16#33#)) OR
 					(reg_q849 AND symb_decoder(16#36#)) OR
 					(reg_q849 AND symb_decoder(16#32#)) OR
 					(reg_q851 AND symb_decoder(16#30#)) OR
 					(reg_q851 AND symb_decoder(16#31#)) OR
 					(reg_q851 AND symb_decoder(16#34#)) OR
 					(reg_q851 AND symb_decoder(16#36#)) OR
 					(reg_q851 AND symb_decoder(16#32#)) OR
 					(reg_q851 AND symb_decoder(16#35#)) OR
 					(reg_q851 AND symb_decoder(16#37#)) OR
 					(reg_q851 AND symb_decoder(16#38#)) OR
 					(reg_q851 AND symb_decoder(16#39#)) OR
 					(reg_q851 AND symb_decoder(16#33#));
reg_q347_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q346 AND symb_decoder(16#53#)) OR
 					(reg_q346 AND symb_decoder(16#73#));
reg_q880_in <= (reg_q876 AND symb_decoder(16#6e#)) OR
 					(reg_q876 AND symb_decoder(16#4e#)) OR
 					(reg_q942 AND symb_decoder(16#6e#)) OR
 					(reg_q942 AND symb_decoder(16#4e#));
reg_q884_in <= (reg_q882 AND symb_decoder(16#74#)) OR
 					(reg_q882 AND symb_decoder(16#54#));
reg_q882_in <= (reg_q880 AND symb_decoder(16#65#)) OR
 					(reg_q880 AND symb_decoder(16#45#));
reg_fullgraph39_init <= "0000";

reg_fullgraph39_sel <= "0" & reg_q882_in & reg_q884_in & reg_q880_in & reg_q347_in & reg_q851_in & reg_q849_in & reg_q1146_in & reg_q843_in & reg_q845_in & reg_q853_in & reg_q823_in & reg_q855_in & reg_q847_in & reg_q540_in & reg_q397_in;

	--coder fullgraph39
with reg_fullgraph39_sel select
reg_fullgraph39_in <=
	"0001" when "0000000000000001",
	"0010" when "0000000000000010",
	"0011" when "0000000000000100",
	"0100" when "0000000000001000",
	"0101" when "0000000000010000",
	"0110" when "0000000000100000",
	"0111" when "0000000001000000",
	"1000" when "0000000010000000",
	"1001" when "0000000100000000",
	"1010" when "0000001000000000",
	"1011" when "0000010000000000",
	"1100" when "0000100000000000",
	"1101" when "0001000000000000",
	"1110" when "0010000000000000",
	"1111" when "0100000000000000",
	"0000" when others;
 --end coder

	p_reg_fullgraph39: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph39 <= reg_fullgraph39_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph39 <= reg_fullgraph39_init;
        else
          reg_fullgraph39 <= reg_fullgraph39_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph39

		reg_q397 <= '1' when reg_fullgraph39 = "0001" else '0'; 
		reg_q540 <= '1' when reg_fullgraph39 = "0010" else '0'; 
		reg_q847 <= '1' when reg_fullgraph39 = "0011" else '0'; 
		reg_q855 <= '1' when reg_fullgraph39 = "0100" else '0'; 
		reg_q823 <= '1' when reg_fullgraph39 = "0101" else '0'; 
		reg_q853 <= '1' when reg_fullgraph39 = "0110" else '0'; 
		reg_q845 <= '1' when reg_fullgraph39 = "0111" else '0'; 
		reg_q843 <= '1' when reg_fullgraph39 = "1000" else '0'; 
		reg_q1146 <= '1' when reg_fullgraph39 = "1001" else '0'; 
		reg_q849 <= '1' when reg_fullgraph39 = "1010" else '0'; 
		reg_q851 <= '1' when reg_fullgraph39 = "1011" else '0'; 
		reg_q347 <= '1' when reg_fullgraph39 = "1100" else '0'; 
		reg_q880 <= '1' when reg_fullgraph39 = "1101" else '0'; 
		reg_q884 <= '1' when reg_fullgraph39 = "1110" else '0'; 
		reg_q882 <= '1' when reg_fullgraph39 = "1111" else '0'; 
--end decoder 

reg_q970_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q970 AND symb_decoder(16#9a#)) OR
 					(reg_q970 AND symb_decoder(16#ab#)) OR
 					(reg_q970 AND symb_decoder(16#c3#)) OR
 					(reg_q970 AND symb_decoder(16#20#)) OR
 					(reg_q970 AND symb_decoder(16#c6#)) OR
 					(reg_q970 AND symb_decoder(16#1a#)) OR
 					(reg_q970 AND symb_decoder(16#fe#)) OR
 					(reg_q970 AND symb_decoder(16#b5#)) OR
 					(reg_q970 AND symb_decoder(16#31#)) OR
 					(reg_q970 AND symb_decoder(16#12#)) OR
 					(reg_q970 AND symb_decoder(16#ae#)) OR
 					(reg_q970 AND symb_decoder(16#b9#)) OR
 					(reg_q970 AND symb_decoder(16#2b#)) OR
 					(reg_q970 AND symb_decoder(16#fa#)) OR
 					(reg_q970 AND symb_decoder(16#19#)) OR
 					(reg_q970 AND symb_decoder(16#27#)) OR
 					(reg_q970 AND symb_decoder(16#5f#)) OR
 					(reg_q970 AND symb_decoder(16#8a#)) OR
 					(reg_q970 AND symb_decoder(16#5b#)) OR
 					(reg_q970 AND symb_decoder(16#18#)) OR
 					(reg_q970 AND symb_decoder(16#4b#)) OR
 					(reg_q970 AND symb_decoder(16#25#)) OR
 					(reg_q970 AND symb_decoder(16#9c#)) OR
 					(reg_q970 AND symb_decoder(16#82#)) OR
 					(reg_q970 AND symb_decoder(16#2c#)) OR
 					(reg_q970 AND symb_decoder(16#be#)) OR
 					(reg_q970 AND symb_decoder(16#21#)) OR
 					(reg_q970 AND symb_decoder(16#08#)) OR
 					(reg_q970 AND symb_decoder(16#09#)) OR
 					(reg_q970 AND symb_decoder(16#64#)) OR
 					(reg_q970 AND symb_decoder(16#d7#)) OR
 					(reg_q970 AND symb_decoder(16#80#)) OR
 					(reg_q970 AND symb_decoder(16#f4#)) OR
 					(reg_q970 AND symb_decoder(16#fc#)) OR
 					(reg_q970 AND symb_decoder(16#59#)) OR
 					(reg_q970 AND symb_decoder(16#9f#)) OR
 					(reg_q970 AND symb_decoder(16#77#)) OR
 					(reg_q970 AND symb_decoder(16#22#)) OR
 					(reg_q970 AND symb_decoder(16#c5#)) OR
 					(reg_q970 AND symb_decoder(16#0d#)) OR
 					(reg_q970 AND symb_decoder(16#b1#)) OR
 					(reg_q970 AND symb_decoder(16#16#)) OR
 					(reg_q970 AND symb_decoder(16#13#)) OR
 					(reg_q970 AND symb_decoder(16#bc#)) OR
 					(reg_q970 AND symb_decoder(16#a6#)) OR
 					(reg_q970 AND symb_decoder(16#9d#)) OR
 					(reg_q970 AND symb_decoder(16#69#)) OR
 					(reg_q970 AND symb_decoder(16#94#)) OR
 					(reg_q970 AND symb_decoder(16#7e#)) OR
 					(reg_q970 AND symb_decoder(16#5c#)) OR
 					(reg_q970 AND symb_decoder(16#9e#)) OR
 					(reg_q970 AND symb_decoder(16#b3#)) OR
 					(reg_q970 AND symb_decoder(16#6e#)) OR
 					(reg_q970 AND symb_decoder(16#7c#)) OR
 					(reg_q970 AND symb_decoder(16#43#)) OR
 					(reg_q970 AND symb_decoder(16#35#)) OR
 					(reg_q970 AND symb_decoder(16#54#)) OR
 					(reg_q970 AND symb_decoder(16#56#)) OR
 					(reg_q970 AND symb_decoder(16#58#)) OR
 					(reg_q970 AND symb_decoder(16#63#)) OR
 					(reg_q970 AND symb_decoder(16#0b#)) OR
 					(reg_q970 AND symb_decoder(16#c0#)) OR
 					(reg_q970 AND symb_decoder(16#72#)) OR
 					(reg_q970 AND symb_decoder(16#2f#)) OR
 					(reg_q970 AND symb_decoder(16#36#)) OR
 					(reg_q970 AND symb_decoder(16#ff#)) OR
 					(reg_q970 AND symb_decoder(16#04#)) OR
 					(reg_q970 AND symb_decoder(16#47#)) OR
 					(reg_q970 AND symb_decoder(16#e5#)) OR
 					(reg_q970 AND symb_decoder(16#ef#)) OR
 					(reg_q970 AND symb_decoder(16#0a#)) OR
 					(reg_q970 AND symb_decoder(16#99#)) OR
 					(reg_q970 AND symb_decoder(16#7a#)) OR
 					(reg_q970 AND symb_decoder(16#e4#)) OR
 					(reg_q970 AND symb_decoder(16#c7#)) OR
 					(reg_q970 AND symb_decoder(16#f8#)) OR
 					(reg_q970 AND symb_decoder(16#84#)) OR
 					(reg_q970 AND symb_decoder(16#b7#)) OR
 					(reg_q970 AND symb_decoder(16#67#)) OR
 					(reg_q970 AND symb_decoder(16#a8#)) OR
 					(reg_q970 AND symb_decoder(16#00#)) OR
 					(reg_q970 AND symb_decoder(16#0f#)) OR
 					(reg_q970 AND symb_decoder(16#ba#)) OR
 					(reg_q970 AND symb_decoder(16#48#)) OR
 					(reg_q970 AND symb_decoder(16#d1#)) OR
 					(reg_q970 AND symb_decoder(16#b6#)) OR
 					(reg_q970 AND symb_decoder(16#d5#)) OR
 					(reg_q970 AND symb_decoder(16#4a#)) OR
 					(reg_q970 AND symb_decoder(16#87#)) OR
 					(reg_q970 AND symb_decoder(16#e7#)) OR
 					(reg_q970 AND symb_decoder(16#24#)) OR
 					(reg_q970 AND symb_decoder(16#3e#)) OR
 					(reg_q970 AND symb_decoder(16#a1#)) OR
 					(reg_q970 AND symb_decoder(16#6d#)) OR
 					(reg_q970 AND symb_decoder(16#e3#)) OR
 					(reg_q970 AND symb_decoder(16#ce#)) OR
 					(reg_q970 AND symb_decoder(16#b4#)) OR
 					(reg_q970 AND symb_decoder(16#d3#)) OR
 					(reg_q970 AND symb_decoder(16#37#)) OR
 					(reg_q970 AND symb_decoder(16#df#)) OR
 					(reg_q970 AND symb_decoder(16#86#)) OR
 					(reg_q970 AND symb_decoder(16#38#)) OR
 					(reg_q970 AND symb_decoder(16#8e#)) OR
 					(reg_q970 AND symb_decoder(16#66#)) OR
 					(reg_q970 AND symb_decoder(16#1d#)) OR
 					(reg_q970 AND symb_decoder(16#f5#)) OR
 					(reg_q970 AND symb_decoder(16#a9#)) OR
 					(reg_q970 AND symb_decoder(16#97#)) OR
 					(reg_q970 AND symb_decoder(16#db#)) OR
 					(reg_q970 AND symb_decoder(16#dc#)) OR
 					(reg_q970 AND symb_decoder(16#fb#)) OR
 					(reg_q970 AND symb_decoder(16#ec#)) OR
 					(reg_q970 AND symb_decoder(16#11#)) OR
 					(reg_q970 AND symb_decoder(16#a5#)) OR
 					(reg_q970 AND symb_decoder(16#42#)) OR
 					(reg_q970 AND symb_decoder(16#70#)) OR
 					(reg_q970 AND symb_decoder(16#e0#)) OR
 					(reg_q970 AND symb_decoder(16#d9#)) OR
 					(reg_q970 AND symb_decoder(16#40#)) OR
 					(reg_q970 AND symb_decoder(16#d2#)) OR
 					(reg_q970 AND symb_decoder(16#f0#)) OR
 					(reg_q970 AND symb_decoder(16#f2#)) OR
 					(reg_q970 AND symb_decoder(16#da#)) OR
 					(reg_q970 AND symb_decoder(16#62#)) OR
 					(reg_q970 AND symb_decoder(16#30#)) OR
 					(reg_q970 AND symb_decoder(16#c9#)) OR
 					(reg_q970 AND symb_decoder(16#af#)) OR
 					(reg_q970 AND symb_decoder(16#75#)) OR
 					(reg_q970 AND symb_decoder(16#5e#)) OR
 					(reg_q970 AND symb_decoder(16#46#)) OR
 					(reg_q970 AND symb_decoder(16#dd#)) OR
 					(reg_q970 AND symb_decoder(16#73#)) OR
 					(reg_q970 AND symb_decoder(16#14#)) OR
 					(reg_q970 AND symb_decoder(16#51#)) OR
 					(reg_q970 AND symb_decoder(16#8b#)) OR
 					(reg_q970 AND symb_decoder(16#26#)) OR
 					(reg_q970 AND symb_decoder(16#f1#)) OR
 					(reg_q970 AND symb_decoder(16#f6#)) OR
 					(reg_q970 AND symb_decoder(16#bb#)) OR
 					(reg_q970 AND symb_decoder(16#1e#)) OR
 					(reg_q970 AND symb_decoder(16#ed#)) OR
 					(reg_q970 AND symb_decoder(16#c1#)) OR
 					(reg_q970 AND symb_decoder(16#2d#)) OR
 					(reg_q970 AND symb_decoder(16#45#)) OR
 					(reg_q970 AND symb_decoder(16#1b#)) OR
 					(reg_q970 AND symb_decoder(16#a0#)) OR
 					(reg_q970 AND symb_decoder(16#ca#)) OR
 					(reg_q970 AND symb_decoder(16#10#)) OR
 					(reg_q970 AND symb_decoder(16#91#)) OR
 					(reg_q970 AND symb_decoder(16#5d#)) OR
 					(reg_q970 AND symb_decoder(16#d4#)) OR
 					(reg_q970 AND symb_decoder(16#28#)) OR
 					(reg_q970 AND symb_decoder(16#34#)) OR
 					(reg_q970 AND symb_decoder(16#ea#)) OR
 					(reg_q970 AND symb_decoder(16#d6#)) OR
 					(reg_q970 AND symb_decoder(16#e2#)) OR
 					(reg_q970 AND symb_decoder(16#1f#)) OR
 					(reg_q970 AND symb_decoder(16#01#)) OR
 					(reg_q970 AND symb_decoder(16#98#)) OR
 					(reg_q970 AND symb_decoder(16#8f#)) OR
 					(reg_q970 AND symb_decoder(16#96#)) OR
 					(reg_q970 AND symb_decoder(16#78#)) OR
 					(reg_q970 AND symb_decoder(16#fd#)) OR
 					(reg_q970 AND symb_decoder(16#2e#)) OR
 					(reg_q970 AND symb_decoder(16#4f#)) OR
 					(reg_q970 AND symb_decoder(16#d8#)) OR
 					(reg_q970 AND symb_decoder(16#cc#)) OR
 					(reg_q970 AND symb_decoder(16#7f#)) OR
 					(reg_q970 AND symb_decoder(16#55#)) OR
 					(reg_q970 AND symb_decoder(16#6f#)) OR
 					(reg_q970 AND symb_decoder(16#e9#)) OR
 					(reg_q970 AND symb_decoder(16#76#)) OR
 					(reg_q970 AND symb_decoder(16#17#)) OR
 					(reg_q970 AND symb_decoder(16#e1#)) OR
 					(reg_q970 AND symb_decoder(16#c2#)) OR
 					(reg_q970 AND symb_decoder(16#53#)) OR
 					(reg_q970 AND symb_decoder(16#f3#)) OR
 					(reg_q970 AND symb_decoder(16#5a#)) OR
 					(reg_q970 AND symb_decoder(16#60#)) OR
 					(reg_q970 AND symb_decoder(16#6c#)) OR
 					(reg_q970 AND symb_decoder(16#c4#)) OR
 					(reg_q970 AND symb_decoder(16#05#)) OR
 					(reg_q970 AND symb_decoder(16#44#)) OR
 					(reg_q970 AND symb_decoder(16#2a#)) OR
 					(reg_q970 AND symb_decoder(16#92#)) OR
 					(reg_q970 AND symb_decoder(16#ee#)) OR
 					(reg_q970 AND symb_decoder(16#39#)) OR
 					(reg_q970 AND symb_decoder(16#aa#)) OR
 					(reg_q970 AND symb_decoder(16#03#)) OR
 					(reg_q970 AND symb_decoder(16#3d#)) OR
 					(reg_q970 AND symb_decoder(16#1c#)) OR
 					(reg_q970 AND symb_decoder(16#74#)) OR
 					(reg_q970 AND symb_decoder(16#89#)) OR
 					(reg_q970 AND symb_decoder(16#79#)) OR
 					(reg_q970 AND symb_decoder(16#ac#)) OR
 					(reg_q970 AND symb_decoder(16#bf#)) OR
 					(reg_q970 AND symb_decoder(16#8d#)) OR
 					(reg_q970 AND symb_decoder(16#b0#)) OR
 					(reg_q970 AND symb_decoder(16#cd#)) OR
 					(reg_q970 AND symb_decoder(16#0c#)) OR
 					(reg_q970 AND symb_decoder(16#07#)) OR
 					(reg_q970 AND symb_decoder(16#61#)) OR
 					(reg_q970 AND symb_decoder(16#88#)) OR
 					(reg_q970 AND symb_decoder(16#de#)) OR
 					(reg_q970 AND symb_decoder(16#a7#)) OR
 					(reg_q970 AND symb_decoder(16#d0#)) OR
 					(reg_q970 AND symb_decoder(16#90#)) OR
 					(reg_q970 AND symb_decoder(16#f9#)) OR
 					(reg_q970 AND symb_decoder(16#eb#)) OR
 					(reg_q970 AND symb_decoder(16#41#)) OR
 					(reg_q970 AND symb_decoder(16#bd#)) OR
 					(reg_q970 AND symb_decoder(16#06#)) OR
 					(reg_q970 AND symb_decoder(16#4d#)) OR
 					(reg_q970 AND symb_decoder(16#50#)) OR
 					(reg_q970 AND symb_decoder(16#0e#)) OR
 					(reg_q970 AND symb_decoder(16#a3#)) OR
 					(reg_q970 AND symb_decoder(16#a4#)) OR
 					(reg_q970 AND symb_decoder(16#7d#)) OR
 					(reg_q970 AND symb_decoder(16#7b#)) OR
 					(reg_q970 AND symb_decoder(16#33#)) OR
 					(reg_q970 AND symb_decoder(16#83#)) OR
 					(reg_q970 AND symb_decoder(16#52#)) OR
 					(reg_q970 AND symb_decoder(16#68#)) OR
 					(reg_q970 AND symb_decoder(16#3b#)) OR
 					(reg_q970 AND symb_decoder(16#3c#)) OR
 					(reg_q970 AND symb_decoder(16#c8#)) OR
 					(reg_q970 AND symb_decoder(16#b8#)) OR
 					(reg_q970 AND symb_decoder(16#85#)) OR
 					(reg_q970 AND symb_decoder(16#81#)) OR
 					(reg_q970 AND symb_decoder(16#9b#)) OR
 					(reg_q970 AND symb_decoder(16#cf#)) OR
 					(reg_q970 AND symb_decoder(16#29#)) OR
 					(reg_q970 AND symb_decoder(16#6b#)) OR
 					(reg_q970 AND symb_decoder(16#3f#)) OR
 					(reg_q970 AND symb_decoder(16#93#)) OR
 					(reg_q970 AND symb_decoder(16#95#)) OR
 					(reg_q970 AND symb_decoder(16#49#)) OR
 					(reg_q970 AND symb_decoder(16#ad#)) OR
 					(reg_q970 AND symb_decoder(16#02#)) OR
 					(reg_q970 AND symb_decoder(16#e8#)) OR
 					(reg_q970 AND symb_decoder(16#32#)) OR
 					(reg_q970 AND symb_decoder(16#8c#)) OR
 					(reg_q970 AND symb_decoder(16#6a#)) OR
 					(reg_q970 AND symb_decoder(16#4e#)) OR
 					(reg_q970 AND symb_decoder(16#71#)) OR
 					(reg_q970 AND symb_decoder(16#57#)) OR
 					(reg_q970 AND symb_decoder(16#f7#)) OR
 					(reg_q970 AND symb_decoder(16#4c#)) OR
 					(reg_q970 AND symb_decoder(16#b2#)) OR
 					(reg_q970 AND symb_decoder(16#e6#)) OR
 					(reg_q970 AND symb_decoder(16#23#)) OR
 					(reg_q970 AND symb_decoder(16#a2#)) OR
 					(reg_q970 AND symb_decoder(16#15#)) OR
 					(reg_q970 AND symb_decoder(16#cb#)) OR
 					(reg_q970 AND symb_decoder(16#65#)) OR
 					(reg_q970 AND symb_decoder(16#3a#));
reg_q970_init <= '0' ;
	p_reg_q970: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q970 <= reg_q970_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q970 <= reg_q970_init;
        else
          reg_q970 <= reg_q970_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1096_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1096 AND symb_decoder(16#6a#)) OR
 					(reg_q1096 AND symb_decoder(16#c9#)) OR
 					(reg_q1096 AND symb_decoder(16#8c#)) OR
 					(reg_q1096 AND symb_decoder(16#1b#)) OR
 					(reg_q1096 AND symb_decoder(16#c8#)) OR
 					(reg_q1096 AND symb_decoder(16#f5#)) OR
 					(reg_q1096 AND symb_decoder(16#58#)) OR
 					(reg_q1096 AND symb_decoder(16#a2#)) OR
 					(reg_q1096 AND symb_decoder(16#b8#)) OR
 					(reg_q1096 AND symb_decoder(16#06#)) OR
 					(reg_q1096 AND symb_decoder(16#80#)) OR
 					(reg_q1096 AND symb_decoder(16#5d#)) OR
 					(reg_q1096 AND symb_decoder(16#f1#)) OR
 					(reg_q1096 AND symb_decoder(16#b3#)) OR
 					(reg_q1096 AND symb_decoder(16#69#)) OR
 					(reg_q1096 AND symb_decoder(16#cc#)) OR
 					(reg_q1096 AND symb_decoder(16#ea#)) OR
 					(reg_q1096 AND symb_decoder(16#13#)) OR
 					(reg_q1096 AND symb_decoder(16#2b#)) OR
 					(reg_q1096 AND symb_decoder(16#e7#)) OR
 					(reg_q1096 AND symb_decoder(16#ed#)) OR
 					(reg_q1096 AND symb_decoder(16#7c#)) OR
 					(reg_q1096 AND symb_decoder(16#b2#)) OR
 					(reg_q1096 AND symb_decoder(16#d3#)) OR
 					(reg_q1096 AND symb_decoder(16#bd#)) OR
 					(reg_q1096 AND symb_decoder(16#78#)) OR
 					(reg_q1096 AND symb_decoder(16#59#)) OR
 					(reg_q1096 AND symb_decoder(16#3f#)) OR
 					(reg_q1096 AND symb_decoder(16#17#)) OR
 					(reg_q1096 AND symb_decoder(16#ac#)) OR
 					(reg_q1096 AND symb_decoder(16#53#)) OR
 					(reg_q1096 AND symb_decoder(16#f9#)) OR
 					(reg_q1096 AND symb_decoder(16#a0#)) OR
 					(reg_q1096 AND symb_decoder(16#e5#)) OR
 					(reg_q1096 AND symb_decoder(16#34#)) OR
 					(reg_q1096 AND symb_decoder(16#4f#)) OR
 					(reg_q1096 AND symb_decoder(16#10#)) OR
 					(reg_q1096 AND symb_decoder(16#56#)) OR
 					(reg_q1096 AND symb_decoder(16#b7#)) OR
 					(reg_q1096 AND symb_decoder(16#cf#)) OR
 					(reg_q1096 AND symb_decoder(16#d1#)) OR
 					(reg_q1096 AND symb_decoder(16#50#)) OR
 					(reg_q1096 AND symb_decoder(16#01#)) OR
 					(reg_q1096 AND symb_decoder(16#0b#)) OR
 					(reg_q1096 AND symb_decoder(16#c7#)) OR
 					(reg_q1096 AND symb_decoder(16#f4#)) OR
 					(reg_q1096 AND symb_decoder(16#87#)) OR
 					(reg_q1096 AND symb_decoder(16#fa#)) OR
 					(reg_q1096 AND symb_decoder(16#9c#)) OR
 					(reg_q1096 AND symb_decoder(16#e6#)) OR
 					(reg_q1096 AND symb_decoder(16#48#)) OR
 					(reg_q1096 AND symb_decoder(16#15#)) OR
 					(reg_q1096 AND symb_decoder(16#f3#)) OR
 					(reg_q1096 AND symb_decoder(16#36#)) OR
 					(reg_q1096 AND symb_decoder(16#1d#)) OR
 					(reg_q1096 AND symb_decoder(16#e3#)) OR
 					(reg_q1096 AND symb_decoder(16#38#)) OR
 					(reg_q1096 AND symb_decoder(16#ce#)) OR
 					(reg_q1096 AND symb_decoder(16#2a#)) OR
 					(reg_q1096 AND symb_decoder(16#fc#)) OR
 					(reg_q1096 AND symb_decoder(16#d0#)) OR
 					(reg_q1096 AND symb_decoder(16#55#)) OR
 					(reg_q1096 AND symb_decoder(16#33#)) OR
 					(reg_q1096 AND symb_decoder(16#ec#)) OR
 					(reg_q1096 AND symb_decoder(16#5a#)) OR
 					(reg_q1096 AND symb_decoder(16#c3#)) OR
 					(reg_q1096 AND symb_decoder(16#81#)) OR
 					(reg_q1096 AND symb_decoder(16#a1#)) OR
 					(reg_q1096 AND symb_decoder(16#96#)) OR
 					(reg_q1096 AND symb_decoder(16#22#)) OR
 					(reg_q1096 AND symb_decoder(16#75#)) OR
 					(reg_q1096 AND symb_decoder(16#be#)) OR
 					(reg_q1096 AND symb_decoder(16#9b#)) OR
 					(reg_q1096 AND symb_decoder(16#7d#)) OR
 					(reg_q1096 AND symb_decoder(16#27#)) OR
 					(reg_q1096 AND symb_decoder(16#0e#)) OR
 					(reg_q1096 AND symb_decoder(16#e2#)) OR
 					(reg_q1096 AND symb_decoder(16#0a#)) OR
 					(reg_q1096 AND symb_decoder(16#7a#)) OR
 					(reg_q1096 AND symb_decoder(16#de#)) OR
 					(reg_q1096 AND symb_decoder(16#2f#)) OR
 					(reg_q1096 AND symb_decoder(16#41#)) OR
 					(reg_q1096 AND symb_decoder(16#29#)) OR
 					(reg_q1096 AND symb_decoder(16#88#)) OR
 					(reg_q1096 AND symb_decoder(16#0c#)) OR
 					(reg_q1096 AND symb_decoder(16#12#)) OR
 					(reg_q1096 AND symb_decoder(16#d5#)) OR
 					(reg_q1096 AND symb_decoder(16#ef#)) OR
 					(reg_q1096 AND symb_decoder(16#43#)) OR
 					(reg_q1096 AND symb_decoder(16#b4#)) OR
 					(reg_q1096 AND symb_decoder(16#25#)) OR
 					(reg_q1096 AND symb_decoder(16#ff#)) OR
 					(reg_q1096 AND symb_decoder(16#54#)) OR
 					(reg_q1096 AND symb_decoder(16#4c#)) OR
 					(reg_q1096 AND symb_decoder(16#6b#)) OR
 					(reg_q1096 AND symb_decoder(16#0d#)) OR
 					(reg_q1096 AND symb_decoder(16#a8#)) OR
 					(reg_q1096 AND symb_decoder(16#c0#)) OR
 					(reg_q1096 AND symb_decoder(16#11#)) OR
 					(reg_q1096 AND symb_decoder(16#19#)) OR
 					(reg_q1096 AND symb_decoder(16#b9#)) OR
 					(reg_q1096 AND symb_decoder(16#bc#)) OR
 					(reg_q1096 AND symb_decoder(16#83#)) OR
 					(reg_q1096 AND symb_decoder(16#ae#)) OR
 					(reg_q1096 AND symb_decoder(16#dd#)) OR
 					(reg_q1096 AND symb_decoder(16#14#)) OR
 					(reg_q1096 AND symb_decoder(16#d2#)) OR
 					(reg_q1096 AND symb_decoder(16#61#)) OR
 					(reg_q1096 AND symb_decoder(16#89#)) OR
 					(reg_q1096 AND symb_decoder(16#5b#)) OR
 					(reg_q1096 AND symb_decoder(16#bf#)) OR
 					(reg_q1096 AND symb_decoder(16#4a#)) OR
 					(reg_q1096 AND symb_decoder(16#71#)) OR
 					(reg_q1096 AND symb_decoder(16#ee#)) OR
 					(reg_q1096 AND symb_decoder(16#66#)) OR
 					(reg_q1096 AND symb_decoder(16#af#)) OR
 					(reg_q1096 AND symb_decoder(16#95#)) OR
 					(reg_q1096 AND symb_decoder(16#23#)) OR
 					(reg_q1096 AND symb_decoder(16#63#)) OR
 					(reg_q1096 AND symb_decoder(16#9e#)) OR
 					(reg_q1096 AND symb_decoder(16#e0#)) OR
 					(reg_q1096 AND symb_decoder(16#8a#)) OR
 					(reg_q1096 AND symb_decoder(16#07#)) OR
 					(reg_q1096 AND symb_decoder(16#8f#)) OR
 					(reg_q1096 AND symb_decoder(16#a6#)) OR
 					(reg_q1096 AND symb_decoder(16#ca#)) OR
 					(reg_q1096 AND symb_decoder(16#cd#)) OR
 					(reg_q1096 AND symb_decoder(16#df#)) OR
 					(reg_q1096 AND symb_decoder(16#45#)) OR
 					(reg_q1096 AND symb_decoder(16#b6#)) OR
 					(reg_q1096 AND symb_decoder(16#e9#)) OR
 					(reg_q1096 AND symb_decoder(16#00#)) OR
 					(reg_q1096 AND symb_decoder(16#2d#)) OR
 					(reg_q1096 AND symb_decoder(16#f8#)) OR
 					(reg_q1096 AND symb_decoder(16#72#)) OR
 					(reg_q1096 AND symb_decoder(16#f6#)) OR
 					(reg_q1096 AND symb_decoder(16#9d#)) OR
 					(reg_q1096 AND symb_decoder(16#dc#)) OR
 					(reg_q1096 AND symb_decoder(16#0f#)) OR
 					(reg_q1096 AND symb_decoder(16#28#)) OR
 					(reg_q1096 AND symb_decoder(16#8d#)) OR
 					(reg_q1096 AND symb_decoder(16#a7#)) OR
 					(reg_q1096 AND symb_decoder(16#62#)) OR
 					(reg_q1096 AND symb_decoder(16#52#)) OR
 					(reg_q1096 AND symb_decoder(16#3b#)) OR
 					(reg_q1096 AND symb_decoder(16#d6#)) OR
 					(reg_q1096 AND symb_decoder(16#44#)) OR
 					(reg_q1096 AND symb_decoder(16#85#)) OR
 					(reg_q1096 AND symb_decoder(16#7b#)) OR
 					(reg_q1096 AND symb_decoder(16#5f#)) OR
 					(reg_q1096 AND symb_decoder(16#37#)) OR
 					(reg_q1096 AND symb_decoder(16#1c#)) OR
 					(reg_q1096 AND symb_decoder(16#e8#)) OR
 					(reg_q1096 AND symb_decoder(16#c2#)) OR
 					(reg_q1096 AND symb_decoder(16#90#)) OR
 					(reg_q1096 AND symb_decoder(16#68#)) OR
 					(reg_q1096 AND symb_decoder(16#76#)) OR
 					(reg_q1096 AND symb_decoder(16#09#)) OR
 					(reg_q1096 AND symb_decoder(16#a9#)) OR
 					(reg_q1096 AND symb_decoder(16#73#)) OR
 					(reg_q1096 AND symb_decoder(16#3a#)) OR
 					(reg_q1096 AND symb_decoder(16#8e#)) OR
 					(reg_q1096 AND symb_decoder(16#84#)) OR
 					(reg_q1096 AND symb_decoder(16#05#)) OR
 					(reg_q1096 AND symb_decoder(16#aa#)) OR
 					(reg_q1096 AND symb_decoder(16#a3#)) OR
 					(reg_q1096 AND symb_decoder(16#a5#)) OR
 					(reg_q1096 AND symb_decoder(16#c5#)) OR
 					(reg_q1096 AND symb_decoder(16#f0#)) OR
 					(reg_q1096 AND symb_decoder(16#93#)) OR
 					(reg_q1096 AND symb_decoder(16#ba#)) OR
 					(reg_q1096 AND symb_decoder(16#b0#)) OR
 					(reg_q1096 AND symb_decoder(16#9a#)) OR
 					(reg_q1096 AND symb_decoder(16#47#)) OR
 					(reg_q1096 AND symb_decoder(16#74#)) OR
 					(reg_q1096 AND symb_decoder(16#1f#)) OR
 					(reg_q1096 AND symb_decoder(16#51#)) OR
 					(reg_q1096 AND symb_decoder(16#03#)) OR
 					(reg_q1096 AND symb_decoder(16#64#)) OR
 					(reg_q1096 AND symb_decoder(16#e1#)) OR
 					(reg_q1096 AND symb_decoder(16#5e#)) OR
 					(reg_q1096 AND symb_decoder(16#31#)) OR
 					(reg_q1096 AND symb_decoder(16#3d#)) OR
 					(reg_q1096 AND symb_decoder(16#26#)) OR
 					(reg_q1096 AND symb_decoder(16#30#)) OR
 					(reg_q1096 AND symb_decoder(16#fb#)) OR
 					(reg_q1096 AND symb_decoder(16#6c#)) OR
 					(reg_q1096 AND symb_decoder(16#49#)) OR
 					(reg_q1096 AND symb_decoder(16#ab#)) OR
 					(reg_q1096 AND symb_decoder(16#94#)) OR
 					(reg_q1096 AND symb_decoder(16#cb#)) OR
 					(reg_q1096 AND symb_decoder(16#d8#)) OR
 					(reg_q1096 AND symb_decoder(16#99#)) OR
 					(reg_q1096 AND symb_decoder(16#7e#)) OR
 					(reg_q1096 AND symb_decoder(16#1a#)) OR
 					(reg_q1096 AND symb_decoder(16#d9#)) OR
 					(reg_q1096 AND symb_decoder(16#92#)) OR
 					(reg_q1096 AND symb_decoder(16#f7#)) OR
 					(reg_q1096 AND symb_decoder(16#79#)) OR
 					(reg_q1096 AND symb_decoder(16#c6#)) OR
 					(reg_q1096 AND symb_decoder(16#fe#)) OR
 					(reg_q1096 AND symb_decoder(16#97#)) OR
 					(reg_q1096 AND symb_decoder(16#3e#)) OR
 					(reg_q1096 AND symb_decoder(16#d7#)) OR
 					(reg_q1096 AND symb_decoder(16#65#)) OR
 					(reg_q1096 AND symb_decoder(16#9f#)) OR
 					(reg_q1096 AND symb_decoder(16#a4#)) OR
 					(reg_q1096 AND symb_decoder(16#6f#)) OR
 					(reg_q1096 AND symb_decoder(16#42#)) OR
 					(reg_q1096 AND symb_decoder(16#67#)) OR
 					(reg_q1096 AND symb_decoder(16#04#)) OR
 					(reg_q1096 AND symb_decoder(16#91#)) OR
 					(reg_q1096 AND symb_decoder(16#98#)) OR
 					(reg_q1096 AND symb_decoder(16#c1#)) OR
 					(reg_q1096 AND symb_decoder(16#bb#)) OR
 					(reg_q1096 AND symb_decoder(16#2c#)) OR
 					(reg_q1096 AND symb_decoder(16#16#)) OR
 					(reg_q1096 AND symb_decoder(16#57#)) OR
 					(reg_q1096 AND symb_decoder(16#4e#)) OR
 					(reg_q1096 AND symb_decoder(16#35#)) OR
 					(reg_q1096 AND symb_decoder(16#8b#)) OR
 					(reg_q1096 AND symb_decoder(16#46#)) OR
 					(reg_q1096 AND symb_decoder(16#08#)) OR
 					(reg_q1096 AND symb_decoder(16#eb#)) OR
 					(reg_q1096 AND symb_decoder(16#fd#)) OR
 					(reg_q1096 AND symb_decoder(16#2e#)) OR
 					(reg_q1096 AND symb_decoder(16#f2#)) OR
 					(reg_q1096 AND symb_decoder(16#4b#)) OR
 					(reg_q1096 AND symb_decoder(16#b1#)) OR
 					(reg_q1096 AND symb_decoder(16#c4#)) OR
 					(reg_q1096 AND symb_decoder(16#21#)) OR
 					(reg_q1096 AND symb_decoder(16#86#)) OR
 					(reg_q1096 AND symb_decoder(16#24#)) OR
 					(reg_q1096 AND symb_decoder(16#1e#)) OR
 					(reg_q1096 AND symb_decoder(16#60#)) OR
 					(reg_q1096 AND symb_decoder(16#77#)) OR
 					(reg_q1096 AND symb_decoder(16#18#)) OR
 					(reg_q1096 AND symb_decoder(16#7f#)) OR
 					(reg_q1096 AND symb_decoder(16#b5#)) OR
 					(reg_q1096 AND symb_decoder(16#32#)) OR
 					(reg_q1096 AND symb_decoder(16#6d#)) OR
 					(reg_q1096 AND symb_decoder(16#20#)) OR
 					(reg_q1096 AND symb_decoder(16#e4#)) OR
 					(reg_q1096 AND symb_decoder(16#40#)) OR
 					(reg_q1096 AND symb_decoder(16#02#)) OR
 					(reg_q1096 AND symb_decoder(16#5c#)) OR
 					(reg_q1096 AND symb_decoder(16#4d#)) OR
 					(reg_q1096 AND symb_decoder(16#ad#)) OR
 					(reg_q1096 AND symb_decoder(16#d4#)) OR
 					(reg_q1096 AND symb_decoder(16#6e#)) OR
 					(reg_q1096 AND symb_decoder(16#3c#)) OR
 					(reg_q1096 AND symb_decoder(16#70#)) OR
 					(reg_q1096 AND symb_decoder(16#82#)) OR
 					(reg_q1096 AND symb_decoder(16#db#)) OR
 					(reg_q1096 AND symb_decoder(16#da#)) OR
 					(reg_q1096 AND symb_decoder(16#39#));
reg_q1096_init <= '0' ;
	p_reg_q1096: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1096 <= reg_q1096_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1096 <= reg_q1096_init;
        else
          reg_q1096 <= reg_q1096_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph42

reg_q2218_in <= (reg_q2218 AND symb_decoder(16#55#)) OR
 					(reg_q2218 AND symb_decoder(16#83#)) OR
 					(reg_q2218 AND symb_decoder(16#9f#)) OR
 					(reg_q2218 AND symb_decoder(16#c1#)) OR
 					(reg_q2218 AND symb_decoder(16#4c#)) OR
 					(reg_q2218 AND symb_decoder(16#47#)) OR
 					(reg_q2218 AND symb_decoder(16#58#)) OR
 					(reg_q2218 AND symb_decoder(16#95#)) OR
 					(reg_q2218 AND symb_decoder(16#2f#)) OR
 					(reg_q2218 AND symb_decoder(16#da#)) OR
 					(reg_q2218 AND symb_decoder(16#f7#)) OR
 					(reg_q2218 AND symb_decoder(16#89#)) OR
 					(reg_q2218 AND symb_decoder(16#68#)) OR
 					(reg_q2218 AND symb_decoder(16#2d#)) OR
 					(reg_q2218 AND symb_decoder(16#17#)) OR
 					(reg_q2218 AND symb_decoder(16#e3#)) OR
 					(reg_q2218 AND symb_decoder(16#1a#)) OR
 					(reg_q2218 AND symb_decoder(16#6e#)) OR
 					(reg_q2218 AND symb_decoder(16#79#)) OR
 					(reg_q2218 AND symb_decoder(16#c9#)) OR
 					(reg_q2218 AND symb_decoder(16#6b#)) OR
 					(reg_q2218 AND symb_decoder(16#3e#)) OR
 					(reg_q2218 AND symb_decoder(16#c4#)) OR
 					(reg_q2218 AND symb_decoder(16#c0#)) OR
 					(reg_q2218 AND symb_decoder(16#8f#)) OR
 					(reg_q2218 AND symb_decoder(16#04#)) OR
 					(reg_q2218 AND symb_decoder(16#72#)) OR
 					(reg_q2218 AND symb_decoder(16#73#)) OR
 					(reg_q2218 AND symb_decoder(16#02#)) OR
 					(reg_q2218 AND symb_decoder(16#c6#)) OR
 					(reg_q2218 AND symb_decoder(16#b1#)) OR
 					(reg_q2218 AND symb_decoder(16#3c#)) OR
 					(reg_q2218 AND symb_decoder(16#59#)) OR
 					(reg_q2218 AND symb_decoder(16#df#)) OR
 					(reg_q2218 AND symb_decoder(16#01#)) OR
 					(reg_q2218 AND symb_decoder(16#d5#)) OR
 					(reg_q2218 AND symb_decoder(16#0f#)) OR
 					(reg_q2218 AND symb_decoder(16#d3#)) OR
 					(reg_q2218 AND symb_decoder(16#bb#)) OR
 					(reg_q2218 AND symb_decoder(16#ec#)) OR
 					(reg_q2218 AND symb_decoder(16#13#)) OR
 					(reg_q2218 AND symb_decoder(16#42#)) OR
 					(reg_q2218 AND symb_decoder(16#f2#)) OR
 					(reg_q2218 AND symb_decoder(16#e6#)) OR
 					(reg_q2218 AND symb_decoder(16#35#)) OR
 					(reg_q2218 AND symb_decoder(16#93#)) OR
 					(reg_q2218 AND symb_decoder(16#8e#)) OR
 					(reg_q2218 AND symb_decoder(16#41#)) OR
 					(reg_q2218 AND symb_decoder(16#06#)) OR
 					(reg_q2218 AND symb_decoder(16#30#)) OR
 					(reg_q2218 AND symb_decoder(16#b3#)) OR
 					(reg_q2218 AND symb_decoder(16#96#)) OR
 					(reg_q2218 AND symb_decoder(16#e9#)) OR
 					(reg_q2218 AND symb_decoder(16#4e#)) OR
 					(reg_q2218 AND symb_decoder(16#34#)) OR
 					(reg_q2218 AND symb_decoder(16#84#)) OR
 					(reg_q2218 AND symb_decoder(16#e1#)) OR
 					(reg_q2218 AND symb_decoder(16#57#)) OR
 					(reg_q2218 AND symb_decoder(16#bc#)) OR
 					(reg_q2218 AND symb_decoder(16#5a#)) OR
 					(reg_q2218 AND symb_decoder(16#18#)) OR
 					(reg_q2218 AND symb_decoder(16#2a#)) OR
 					(reg_q2218 AND symb_decoder(16#f0#)) OR
 					(reg_q2218 AND symb_decoder(16#b7#)) OR
 					(reg_q2218 AND symb_decoder(16#bf#)) OR
 					(reg_q2218 AND symb_decoder(16#48#)) OR
 					(reg_q2218 AND symb_decoder(16#32#)) OR
 					(reg_q2218 AND symb_decoder(16#b6#)) OR
 					(reg_q2218 AND symb_decoder(16#d2#)) OR
 					(reg_q2218 AND symb_decoder(16#e2#)) OR
 					(reg_q2218 AND symb_decoder(16#44#)) OR
 					(reg_q2218 AND symb_decoder(16#54#)) OR
 					(reg_q2218 AND symb_decoder(16#52#)) OR
 					(reg_q2218 AND symb_decoder(16#29#)) OR
 					(reg_q2218 AND symb_decoder(16#cd#)) OR
 					(reg_q2218 AND symb_decoder(16#5b#)) OR
 					(reg_q2218 AND symb_decoder(16#6a#)) OR
 					(reg_q2218 AND symb_decoder(16#63#)) OR
 					(reg_q2218 AND symb_decoder(16#74#)) OR
 					(reg_q2218 AND symb_decoder(16#ef#)) OR
 					(reg_q2218 AND symb_decoder(16#92#)) OR
 					(reg_q2218 AND symb_decoder(16#e5#)) OR
 					(reg_q2218 AND symb_decoder(16#26#)) OR
 					(reg_q2218 AND symb_decoder(16#91#)) OR
 					(reg_q2218 AND symb_decoder(16#88#)) OR
 					(reg_q2218 AND symb_decoder(16#64#)) OR
 					(reg_q2218 AND symb_decoder(16#1d#)) OR
 					(reg_q2218 AND symb_decoder(16#85#)) OR
 					(reg_q2218 AND symb_decoder(16#8d#)) OR
 					(reg_q2218 AND symb_decoder(16#1e#)) OR
 					(reg_q2218 AND symb_decoder(16#7d#)) OR
 					(reg_q2218 AND symb_decoder(16#dc#)) OR
 					(reg_q2218 AND symb_decoder(16#cb#)) OR
 					(reg_q2218 AND symb_decoder(16#43#)) OR
 					(reg_q2218 AND symb_decoder(16#21#)) OR
 					(reg_q2218 AND symb_decoder(16#fd#)) OR
 					(reg_q2218 AND symb_decoder(16#cf#)) OR
 					(reg_q2218 AND symb_decoder(16#d4#)) OR
 					(reg_q2218 AND symb_decoder(16#82#)) OR
 					(reg_q2218 AND symb_decoder(16#fb#)) OR
 					(reg_q2218 AND symb_decoder(16#9d#)) OR
 					(reg_q2218 AND symb_decoder(16#f3#)) OR
 					(reg_q2218 AND symb_decoder(16#b2#)) OR
 					(reg_q2218 AND symb_decoder(16#9e#)) OR
 					(reg_q2218 AND symb_decoder(16#77#)) OR
 					(reg_q2218 AND symb_decoder(16#a6#)) OR
 					(reg_q2218 AND symb_decoder(16#45#)) OR
 					(reg_q2218 AND symb_decoder(16#10#)) OR
 					(reg_q2218 AND symb_decoder(16#a4#)) OR
 					(reg_q2218 AND symb_decoder(16#51#)) OR
 					(reg_q2218 AND symb_decoder(16#61#)) OR
 					(reg_q2218 AND symb_decoder(16#25#)) OR
 					(reg_q2218 AND symb_decoder(16#27#)) OR
 					(reg_q2218 AND symb_decoder(16#28#)) OR
 					(reg_q2218 AND symb_decoder(16#ee#)) OR
 					(reg_q2218 AND symb_decoder(16#7c#)) OR
 					(reg_q2218 AND symb_decoder(16#ff#)) OR
 					(reg_q2218 AND symb_decoder(16#a2#)) OR
 					(reg_q2218 AND symb_decoder(16#f8#)) OR
 					(reg_q2218 AND symb_decoder(16#cc#)) OR
 					(reg_q2218 AND symb_decoder(16#4d#)) OR
 					(reg_q2218 AND symb_decoder(16#66#)) OR
 					(reg_q2218 AND symb_decoder(16#d9#)) OR
 					(reg_q2218 AND symb_decoder(16#24#)) OR
 					(reg_q2218 AND symb_decoder(16#ed#)) OR
 					(reg_q2218 AND symb_decoder(16#eb#)) OR
 					(reg_q2218 AND symb_decoder(16#ce#)) OR
 					(reg_q2218 AND symb_decoder(16#1c#)) OR
 					(reg_q2218 AND symb_decoder(16#a7#)) OR
 					(reg_q2218 AND symb_decoder(16#75#)) OR
 					(reg_q2218 AND symb_decoder(16#7e#)) OR
 					(reg_q2218 AND symb_decoder(16#80#)) OR
 					(reg_q2218 AND symb_decoder(16#40#)) OR
 					(reg_q2218 AND symb_decoder(16#5f#)) OR
 					(reg_q2218 AND symb_decoder(16#c2#)) OR
 					(reg_q2218 AND symb_decoder(16#be#)) OR
 					(reg_q2218 AND symb_decoder(16#c3#)) OR
 					(reg_q2218 AND symb_decoder(16#90#)) OR
 					(reg_q2218 AND symb_decoder(16#fc#)) OR
 					(reg_q2218 AND symb_decoder(16#71#)) OR
 					(reg_q2218 AND symb_decoder(16#fe#)) OR
 					(reg_q2218 AND symb_decoder(16#db#)) OR
 					(reg_q2218 AND symb_decoder(16#00#)) OR
 					(reg_q2218 AND symb_decoder(16#49#)) OR
 					(reg_q2218 AND symb_decoder(16#6c#)) OR
 					(reg_q2218 AND symb_decoder(16#d8#)) OR
 					(reg_q2218 AND symb_decoder(16#7a#)) OR
 					(reg_q2218 AND symb_decoder(16#22#)) OR
 					(reg_q2218 AND symb_decoder(16#3f#)) OR
 					(reg_q2218 AND symb_decoder(16#af#)) OR
 					(reg_q2218 AND symb_decoder(16#f6#)) OR
 					(reg_q2218 AND symb_decoder(16#3d#)) OR
 					(reg_q2218 AND symb_decoder(16#56#)) OR
 					(reg_q2218 AND symb_decoder(16#ad#)) OR
 					(reg_q2218 AND symb_decoder(16#4f#)) OR
 					(reg_q2218 AND symb_decoder(16#12#)) OR
 					(reg_q2218 AND symb_decoder(16#ba#)) OR
 					(reg_q2218 AND symb_decoder(16#1b#)) OR
 					(reg_q2218 AND symb_decoder(16#f1#)) OR
 					(reg_q2218 AND symb_decoder(16#9a#)) OR
 					(reg_q2218 AND symb_decoder(16#87#)) OR
 					(reg_q2218 AND symb_decoder(16#b0#)) OR
 					(reg_q2218 AND symb_decoder(16#bd#)) OR
 					(reg_q2218 AND symb_decoder(16#ab#)) OR
 					(reg_q2218 AND symb_decoder(16#b4#)) OR
 					(reg_q2218 AND symb_decoder(16#d1#)) OR
 					(reg_q2218 AND symb_decoder(16#9b#)) OR
 					(reg_q2218 AND symb_decoder(16#ea#)) OR
 					(reg_q2218 AND symb_decoder(16#4b#)) OR
 					(reg_q2218 AND symb_decoder(16#8b#)) OR
 					(reg_q2218 AND symb_decoder(16#37#)) OR
 					(reg_q2218 AND symb_decoder(16#15#)) OR
 					(reg_q2218 AND symb_decoder(16#03#)) OR
 					(reg_q2218 AND symb_decoder(16#a3#)) OR
 					(reg_q2218 AND symb_decoder(16#78#)) OR
 					(reg_q2218 AND symb_decoder(16#6d#)) OR
 					(reg_q2218 AND symb_decoder(16#fa#)) OR
 					(reg_q2218 AND symb_decoder(16#b9#)) OR
 					(reg_q2218 AND symb_decoder(16#33#)) OR
 					(reg_q2218 AND symb_decoder(16#b5#)) OR
 					(reg_q2218 AND symb_decoder(16#e4#)) OR
 					(reg_q2218 AND symb_decoder(16#c5#)) OR
 					(reg_q2218 AND symb_decoder(16#7b#)) OR
 					(reg_q2218 AND symb_decoder(16#86#)) OR
 					(reg_q2218 AND symb_decoder(16#23#)) OR
 					(reg_q2218 AND symb_decoder(16#0e#)) OR
 					(reg_q2218 AND symb_decoder(16#0c#)) OR
 					(reg_q2218 AND symb_decoder(16#e8#)) OR
 					(reg_q2218 AND symb_decoder(16#d0#)) OR
 					(reg_q2218 AND symb_decoder(16#e0#)) OR
 					(reg_q2218 AND symb_decoder(16#5d#)) OR
 					(reg_q2218 AND symb_decoder(16#62#)) OR
 					(reg_q2218 AND symb_decoder(16#b8#)) OR
 					(reg_q2218 AND symb_decoder(16#8a#)) OR
 					(reg_q2218 AND symb_decoder(16#a5#)) OR
 					(reg_q2218 AND symb_decoder(16#ac#)) OR
 					(reg_q2218 AND symb_decoder(16#ae#)) OR
 					(reg_q2218 AND symb_decoder(16#6f#)) OR
 					(reg_q2218 AND symb_decoder(16#1f#)) OR
 					(reg_q2218 AND symb_decoder(16#3a#)) OR
 					(reg_q2218 AND symb_decoder(16#94#)) OR
 					(reg_q2218 AND symb_decoder(16#99#)) OR
 					(reg_q2218 AND symb_decoder(16#0b#)) OR
 					(reg_q2218 AND symb_decoder(16#50#)) OR
 					(reg_q2218 AND symb_decoder(16#c7#)) OR
 					(reg_q2218 AND symb_decoder(16#3b#)) OR
 					(reg_q2218 AND symb_decoder(16#98#)) OR
 					(reg_q2218 AND symb_decoder(16#36#)) OR
 					(reg_q2218 AND symb_decoder(16#69#)) OR
 					(reg_q2218 AND symb_decoder(16#e7#)) OR
 					(reg_q2218 AND symb_decoder(16#ca#)) OR
 					(reg_q2218 AND symb_decoder(16#53#)) OR
 					(reg_q2218 AND symb_decoder(16#20#)) OR
 					(reg_q2218 AND symb_decoder(16#f9#)) OR
 					(reg_q2218 AND symb_decoder(16#f4#)) OR
 					(reg_q2218 AND symb_decoder(16#09#)) OR
 					(reg_q2218 AND symb_decoder(16#14#)) OR
 					(reg_q2218 AND symb_decoder(16#65#)) OR
 					(reg_q2218 AND symb_decoder(16#5c#)) OR
 					(reg_q2218 AND symb_decoder(16#39#)) OR
 					(reg_q2218 AND symb_decoder(16#2b#)) OR
 					(reg_q2218 AND symb_decoder(16#60#)) OR
 					(reg_q2218 AND symb_decoder(16#67#)) OR
 					(reg_q2218 AND symb_decoder(16#2c#)) OR
 					(reg_q2218 AND symb_decoder(16#70#)) OR
 					(reg_q2218 AND symb_decoder(16#aa#)) OR
 					(reg_q2218 AND symb_decoder(16#a0#)) OR
 					(reg_q2218 AND symb_decoder(16#8c#)) OR
 					(reg_q2218 AND symb_decoder(16#de#)) OR
 					(reg_q2218 AND symb_decoder(16#2e#)) OR
 					(reg_q2218 AND symb_decoder(16#9c#)) OR
 					(reg_q2218 AND symb_decoder(16#a9#)) OR
 					(reg_q2218 AND symb_decoder(16#19#)) OR
 					(reg_q2218 AND symb_decoder(16#46#)) OR
 					(reg_q2218 AND symb_decoder(16#07#)) OR
 					(reg_q2218 AND symb_decoder(16#a8#)) OR
 					(reg_q2218 AND symb_decoder(16#38#)) OR
 					(reg_q2218 AND symb_decoder(16#d7#)) OR
 					(reg_q2218 AND symb_decoder(16#4a#)) OR
 					(reg_q2218 AND symb_decoder(16#08#)) OR
 					(reg_q2218 AND symb_decoder(16#11#)) OR
 					(reg_q2218 AND symb_decoder(16#7f#)) OR
 					(reg_q2218 AND symb_decoder(16#05#)) OR
 					(reg_q2218 AND symb_decoder(16#dd#)) OR
 					(reg_q2218 AND symb_decoder(16#97#)) OR
 					(reg_q2218 AND symb_decoder(16#16#)) OR
 					(reg_q2218 AND symb_decoder(16#76#)) OR
 					(reg_q2218 AND symb_decoder(16#81#)) OR
 					(reg_q2218 AND symb_decoder(16#5e#)) OR
 					(reg_q2218 AND symb_decoder(16#a1#)) OR
 					(reg_q2218 AND symb_decoder(16#c8#)) OR
 					(reg_q2218 AND symb_decoder(16#31#)) OR
 					(reg_q2218 AND symb_decoder(16#d6#)) OR
 					(reg_q2218 AND symb_decoder(16#f5#)) OR
 					(reg_q2112 AND symb_decoder(16#c2#)) OR
 					(reg_q2112 AND symb_decoder(16#19#)) OR
 					(reg_q2112 AND symb_decoder(16#70#)) OR
 					(reg_q2112 AND symb_decoder(16#e5#)) OR
 					(reg_q2112 AND symb_decoder(16#6e#)) OR
 					(reg_q2112 AND symb_decoder(16#a9#)) OR
 					(reg_q2112 AND symb_decoder(16#80#)) OR
 					(reg_q2112 AND symb_decoder(16#22#)) OR
 					(reg_q2112 AND symb_decoder(16#4e#)) OR
 					(reg_q2112 AND symb_decoder(16#02#)) OR
 					(reg_q2112 AND symb_decoder(16#ae#)) OR
 					(reg_q2112 AND symb_decoder(16#23#)) OR
 					(reg_q2112 AND symb_decoder(16#b8#)) OR
 					(reg_q2112 AND symb_decoder(16#f2#)) OR
 					(reg_q2112 AND symb_decoder(16#64#)) OR
 					(reg_q2112 AND symb_decoder(16#b5#)) OR
 					(reg_q2112 AND symb_decoder(16#96#)) OR
 					(reg_q2112 AND symb_decoder(16#c6#)) OR
 					(reg_q2112 AND symb_decoder(16#15#)) OR
 					(reg_q2112 AND symb_decoder(16#ee#)) OR
 					(reg_q2112 AND symb_decoder(16#00#)) OR
 					(reg_q2112 AND symb_decoder(16#9f#)) OR
 					(reg_q2112 AND symb_decoder(16#5d#)) OR
 					(reg_q2112 AND symb_decoder(16#60#)) OR
 					(reg_q2112 AND symb_decoder(16#f6#)) OR
 					(reg_q2112 AND symb_decoder(16#a7#)) OR
 					(reg_q2112 AND symb_decoder(16#af#)) OR
 					(reg_q2112 AND symb_decoder(16#52#)) OR
 					(reg_q2112 AND symb_decoder(16#ff#)) OR
 					(reg_q2112 AND symb_decoder(16#71#)) OR
 					(reg_q2112 AND symb_decoder(16#41#)) OR
 					(reg_q2112 AND symb_decoder(16#75#)) OR
 					(reg_q2112 AND symb_decoder(16#27#)) OR
 					(reg_q2112 AND symb_decoder(16#eb#)) OR
 					(reg_q2112 AND symb_decoder(16#4a#)) OR
 					(reg_q2112 AND symb_decoder(16#5c#)) OR
 					(reg_q2112 AND symb_decoder(16#24#)) OR
 					(reg_q2112 AND symb_decoder(16#a6#)) OR
 					(reg_q2112 AND symb_decoder(16#50#)) OR
 					(reg_q2112 AND symb_decoder(16#e3#)) OR
 					(reg_q2112 AND symb_decoder(16#62#)) OR
 					(reg_q2112 AND symb_decoder(16#7f#)) OR
 					(reg_q2112 AND symb_decoder(16#a5#)) OR
 					(reg_q2112 AND symb_decoder(16#3c#)) OR
 					(reg_q2112 AND symb_decoder(16#ce#)) OR
 					(reg_q2112 AND symb_decoder(16#34#)) OR
 					(reg_q2112 AND symb_decoder(16#e1#)) OR
 					(reg_q2112 AND symb_decoder(16#c9#)) OR
 					(reg_q2112 AND symb_decoder(16#b1#)) OR
 					(reg_q2112 AND symb_decoder(16#08#)) OR
 					(reg_q2112 AND symb_decoder(16#65#)) OR
 					(reg_q2112 AND symb_decoder(16#a2#)) OR
 					(reg_q2112 AND symb_decoder(16#29#)) OR
 					(reg_q2112 AND symb_decoder(16#f0#)) OR
 					(reg_q2112 AND symb_decoder(16#2f#)) OR
 					(reg_q2112 AND symb_decoder(16#33#)) OR
 					(reg_q2112 AND symb_decoder(16#59#)) OR
 					(reg_q2112 AND symb_decoder(16#c4#)) OR
 					(reg_q2112 AND symb_decoder(16#e7#)) OR
 					(reg_q2112 AND symb_decoder(16#95#)) OR
 					(reg_q2112 AND symb_decoder(16#4f#)) OR
 					(reg_q2112 AND symb_decoder(16#2d#)) OR
 					(reg_q2112 AND symb_decoder(16#f5#)) OR
 					(reg_q2112 AND symb_decoder(16#37#)) OR
 					(reg_q2112 AND symb_decoder(16#b0#)) OR
 					(reg_q2112 AND symb_decoder(16#1e#)) OR
 					(reg_q2112 AND symb_decoder(16#48#)) OR
 					(reg_q2112 AND symb_decoder(16#ac#)) OR
 					(reg_q2112 AND symb_decoder(16#40#)) OR
 					(reg_q2112 AND symb_decoder(16#17#)) OR
 					(reg_q2112 AND symb_decoder(16#ba#)) OR
 					(reg_q2112 AND symb_decoder(16#ec#)) OR
 					(reg_q2112 AND symb_decoder(16#55#)) OR
 					(reg_q2112 AND symb_decoder(16#77#)) OR
 					(reg_q2112 AND symb_decoder(16#e4#)) OR
 					(reg_q2112 AND symb_decoder(16#94#)) OR
 					(reg_q2112 AND symb_decoder(16#78#)) OR
 					(reg_q2112 AND symb_decoder(16#f4#)) OR
 					(reg_q2112 AND symb_decoder(16#82#)) OR
 					(reg_q2112 AND symb_decoder(16#74#)) OR
 					(reg_q2112 AND symb_decoder(16#a0#)) OR
 					(reg_q2112 AND symb_decoder(16#ab#)) OR
 					(reg_q2112 AND symb_decoder(16#35#)) OR
 					(reg_q2112 AND symb_decoder(16#07#)) OR
 					(reg_q2112 AND symb_decoder(16#6f#)) OR
 					(reg_q2112 AND symb_decoder(16#1a#)) OR
 					(reg_q2112 AND symb_decoder(16#3f#)) OR
 					(reg_q2112 AND symb_decoder(16#4b#)) OR
 					(reg_q2112 AND symb_decoder(16#fa#)) OR
 					(reg_q2112 AND symb_decoder(16#47#)) OR
 					(reg_q2112 AND symb_decoder(16#21#)) OR
 					(reg_q2112 AND symb_decoder(16#de#)) OR
 					(reg_q2112 AND symb_decoder(16#d7#)) OR
 					(reg_q2112 AND symb_decoder(16#93#)) OR
 					(reg_q2112 AND symb_decoder(16#5a#)) OR
 					(reg_q2112 AND symb_decoder(16#d0#)) OR
 					(reg_q2112 AND symb_decoder(16#c1#)) OR
 					(reg_q2112 AND symb_decoder(16#90#)) OR
 					(reg_q2112 AND symb_decoder(16#46#)) OR
 					(reg_q2112 AND symb_decoder(16#f1#)) OR
 					(reg_q2112 AND symb_decoder(16#a1#)) OR
 					(reg_q2112 AND symb_decoder(16#f7#)) OR
 					(reg_q2112 AND symb_decoder(16#c3#)) OR
 					(reg_q2112 AND symb_decoder(16#31#)) OR
 					(reg_q2112 AND symb_decoder(16#68#)) OR
 					(reg_q2112 AND symb_decoder(16#28#)) OR
 					(reg_q2112 AND symb_decoder(16#92#)) OR
 					(reg_q2112 AND symb_decoder(16#87#)) OR
 					(reg_q2112 AND symb_decoder(16#8e#)) OR
 					(reg_q2112 AND symb_decoder(16#d2#)) OR
 					(reg_q2112 AND symb_decoder(16#be#)) OR
 					(reg_q2112 AND symb_decoder(16#cd#)) OR
 					(reg_q2112 AND symb_decoder(16#6d#)) OR
 					(reg_q2112 AND symb_decoder(16#fb#)) OR
 					(reg_q2112 AND symb_decoder(16#5f#)) OR
 					(reg_q2112 AND symb_decoder(16#1d#)) OR
 					(reg_q2112 AND symb_decoder(16#6c#)) OR
 					(reg_q2112 AND symb_decoder(16#e6#)) OR
 					(reg_q2112 AND symb_decoder(16#fe#)) OR
 					(reg_q2112 AND symb_decoder(16#99#)) OR
 					(reg_q2112 AND symb_decoder(16#a4#)) OR
 					(reg_q2112 AND symb_decoder(16#0b#)) OR
 					(reg_q2112 AND symb_decoder(16#b2#)) OR
 					(reg_q2112 AND symb_decoder(16#bd#)) OR
 					(reg_q2112 AND symb_decoder(16#b6#)) OR
 					(reg_q2112 AND symb_decoder(16#61#)) OR
 					(reg_q2112 AND symb_decoder(16#45#)) OR
 					(reg_q2112 AND symb_decoder(16#25#)) OR
 					(reg_q2112 AND symb_decoder(16#57#)) OR
 					(reg_q2112 AND symb_decoder(16#0e#)) OR
 					(reg_q2112 AND symb_decoder(16#8b#)) OR
 					(reg_q2112 AND symb_decoder(16#7b#)) OR
 					(reg_q2112 AND symb_decoder(16#e8#)) OR
 					(reg_q2112 AND symb_decoder(16#3a#)) OR
 					(reg_q2112 AND symb_decoder(16#d4#)) OR
 					(reg_q2112 AND symb_decoder(16#2a#)) OR
 					(reg_q2112 AND symb_decoder(16#f9#)) OR
 					(reg_q2112 AND symb_decoder(16#1f#)) OR
 					(reg_q2112 AND symb_decoder(16#8a#)) OR
 					(reg_q2112 AND symb_decoder(16#e9#)) OR
 					(reg_q2112 AND symb_decoder(16#44#)) OR
 					(reg_q2112 AND symb_decoder(16#d9#)) OR
 					(reg_q2112 AND symb_decoder(16#b7#)) OR
 					(reg_q2112 AND symb_decoder(16#2e#)) OR
 					(reg_q2112 AND symb_decoder(16#b4#)) OR
 					(reg_q2112 AND symb_decoder(16#85#)) OR
 					(reg_q2112 AND symb_decoder(16#d6#)) OR
 					(reg_q2112 AND symb_decoder(16#0f#)) OR
 					(reg_q2112 AND symb_decoder(16#c7#)) OR
 					(reg_q2112 AND symb_decoder(16#32#)) OR
 					(reg_q2112 AND symb_decoder(16#7a#)) OR
 					(reg_q2112 AND symb_decoder(16#8d#)) OR
 					(reg_q2112 AND symb_decoder(16#98#)) OR
 					(reg_q2112 AND symb_decoder(16#0c#)) OR
 					(reg_q2112 AND symb_decoder(16#3b#)) OR
 					(reg_q2112 AND symb_decoder(16#a3#)) OR
 					(reg_q2112 AND symb_decoder(16#c8#)) OR
 					(reg_q2112 AND symb_decoder(16#dd#)) OR
 					(reg_q2112 AND symb_decoder(16#09#)) OR
 					(reg_q2112 AND symb_decoder(16#16#)) OR
 					(reg_q2112 AND symb_decoder(16#df#)) OR
 					(reg_q2112 AND symb_decoder(16#11#)) OR
 					(reg_q2112 AND symb_decoder(16#ef#)) OR
 					(reg_q2112 AND symb_decoder(16#04#)) OR
 					(reg_q2112 AND symb_decoder(16#14#)) OR
 					(reg_q2112 AND symb_decoder(16#89#)) OR
 					(reg_q2112 AND symb_decoder(16#aa#)) OR
 					(reg_q2112 AND symb_decoder(16#03#)) OR
 					(reg_q2112 AND symb_decoder(16#ed#)) OR
 					(reg_q2112 AND symb_decoder(16#2c#)) OR
 					(reg_q2112 AND symb_decoder(16#39#)) OR
 					(reg_q2112 AND symb_decoder(16#4c#)) OR
 					(reg_q2112 AND symb_decoder(16#bf#)) OR
 					(reg_q2112 AND symb_decoder(16#86#)) OR
 					(reg_q2112 AND symb_decoder(16#42#)) OR
 					(reg_q2112 AND symb_decoder(16#8c#)) OR
 					(reg_q2112 AND symb_decoder(16#18#)) OR
 					(reg_q2112 AND symb_decoder(16#ad#)) OR
 					(reg_q2112 AND symb_decoder(16#91#)) OR
 					(reg_q2112 AND symb_decoder(16#7e#)) OR
 					(reg_q2112 AND symb_decoder(16#1b#)) OR
 					(reg_q2112 AND symb_decoder(16#54#)) OR
 					(reg_q2112 AND symb_decoder(16#58#)) OR
 					(reg_q2112 AND symb_decoder(16#5b#)) OR
 					(reg_q2112 AND symb_decoder(16#da#)) OR
 					(reg_q2112 AND symb_decoder(16#63#)) OR
 					(reg_q2112 AND symb_decoder(16#9a#)) OR
 					(reg_q2112 AND symb_decoder(16#53#)) OR
 					(reg_q2112 AND symb_decoder(16#cb#)) OR
 					(reg_q2112 AND symb_decoder(16#e0#)) OR
 					(reg_q2112 AND symb_decoder(16#2b#)) OR
 					(reg_q2112 AND symb_decoder(16#cf#)) OR
 					(reg_q2112 AND symb_decoder(16#9b#)) OR
 					(reg_q2112 AND symb_decoder(16#cc#)) OR
 					(reg_q2112 AND symb_decoder(16#79#)) OR
 					(reg_q2112 AND symb_decoder(16#43#)) OR
 					(reg_q2112 AND symb_decoder(16#9c#)) OR
 					(reg_q2112 AND symb_decoder(16#3d#)) OR
 					(reg_q2112 AND symb_decoder(16#c5#)) OR
 					(reg_q2112 AND symb_decoder(16#d3#)) OR
 					(reg_q2112 AND symb_decoder(16#6b#)) OR
 					(reg_q2112 AND symb_decoder(16#7d#)) OR
 					(reg_q2112 AND symb_decoder(16#e2#)) OR
 					(reg_q2112 AND symb_decoder(16#73#)) OR
 					(reg_q2112 AND symb_decoder(16#4d#)) OR
 					(reg_q2112 AND symb_decoder(16#56#)) OR
 					(reg_q2112 AND symb_decoder(16#88#)) OR
 					(reg_q2112 AND symb_decoder(16#81#)) OR
 					(reg_q2112 AND symb_decoder(16#ea#)) OR
 					(reg_q2112 AND symb_decoder(16#36#)) OR
 					(reg_q2112 AND symb_decoder(16#10#)) OR
 					(reg_q2112 AND symb_decoder(16#1c#)) OR
 					(reg_q2112 AND symb_decoder(16#20#)) OR
 					(reg_q2112 AND symb_decoder(16#69#)) OR
 					(reg_q2112 AND symb_decoder(16#76#)) OR
 					(reg_q2112 AND symb_decoder(16#3e#)) OR
 					(reg_q2112 AND symb_decoder(16#51#)) OR
 					(reg_q2112 AND symb_decoder(16#01#)) OR
 					(reg_q2112 AND symb_decoder(16#ca#)) OR
 					(reg_q2112 AND symb_decoder(16#84#)) OR
 					(reg_q2112 AND symb_decoder(16#f3#)) OR
 					(reg_q2112 AND symb_decoder(16#fd#)) OR
 					(reg_q2112 AND symb_decoder(16#26#)) OR
 					(reg_q2112 AND symb_decoder(16#f8#)) OR
 					(reg_q2112 AND symb_decoder(16#7c#)) OR
 					(reg_q2112 AND symb_decoder(16#b3#)) OR
 					(reg_q2112 AND symb_decoder(16#9e#)) OR
 					(reg_q2112 AND symb_decoder(16#c0#)) OR
 					(reg_q2112 AND symb_decoder(16#66#)) OR
 					(reg_q2112 AND symb_decoder(16#12#)) OR
 					(reg_q2112 AND symb_decoder(16#49#)) OR
 					(reg_q2112 AND symb_decoder(16#b9#)) OR
 					(reg_q2112 AND symb_decoder(16#13#)) OR
 					(reg_q2112 AND symb_decoder(16#97#)) OR
 					(reg_q2112 AND symb_decoder(16#72#)) OR
 					(reg_q2112 AND symb_decoder(16#5e#)) OR
 					(reg_q2112 AND symb_decoder(16#db#)) OR
 					(reg_q2112 AND symb_decoder(16#bb#)) OR
 					(reg_q2112 AND symb_decoder(16#d5#)) OR
 					(reg_q2112 AND symb_decoder(16#05#)) OR
 					(reg_q2112 AND symb_decoder(16#d8#)) OR
 					(reg_q2112 AND symb_decoder(16#6a#)) OR
 					(reg_q2112 AND symb_decoder(16#bc#)) OR
 					(reg_q2112 AND symb_decoder(16#06#)) OR
 					(reg_q2112 AND symb_decoder(16#d1#)) OR
 					(reg_q2112 AND symb_decoder(16#9d#)) OR
 					(reg_q2112 AND symb_decoder(16#8f#)) OR
 					(reg_q2112 AND symb_decoder(16#67#)) OR
 					(reg_q2112 AND symb_decoder(16#fc#)) OR
 					(reg_q2112 AND symb_decoder(16#38#)) OR
 					(reg_q2112 AND symb_decoder(16#dc#)) OR
 					(reg_q2112 AND symb_decoder(16#a8#)) OR
 					(reg_q2112 AND symb_decoder(16#30#)) OR
 					(reg_q2112 AND symb_decoder(16#83#));
reg_q546_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q545 AND symb_decoder(16#0d#)) OR
 					(reg_q545 AND symb_decoder(16#0a#));
reg_q592_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q591 AND symb_decoder(16#73#)) OR
 					(reg_q591 AND symb_decoder(16#53#));
reg_fullgraph42_init <= "00";

reg_fullgraph42_sel <= "0" & reg_q592_in & reg_q546_in & reg_q2218_in;

	--coder fullgraph42
with reg_fullgraph42_sel select
reg_fullgraph42_in <=
	"01" when "0001",
	"10" when "0010",
	"11" when "0100",
	"00" when others;
 --end coder

	p_reg_fullgraph42: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph42 <= reg_fullgraph42_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph42 <= reg_fullgraph42_init;
        else
          reg_fullgraph42 <= reg_fullgraph42_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph42

		reg_q2218 <= '1' when reg_fullgraph42 = "01" else '0'; 
		reg_q546 <= '1' when reg_fullgraph42 = "10" else '0'; 
		reg_q592 <= '1' when reg_fullgraph42 = "11" else '0'; 
--end decoder 

reg_q2056_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q2056 AND symb_decoder(16#f9#)) OR
 					(reg_q2056 AND symb_decoder(16#f3#)) OR
 					(reg_q2056 AND symb_decoder(16#34#)) OR
 					(reg_q2056 AND symb_decoder(16#e3#)) OR
 					(reg_q2056 AND symb_decoder(16#24#)) OR
 					(reg_q2056 AND symb_decoder(16#dd#)) OR
 					(reg_q2056 AND symb_decoder(16#91#)) OR
 					(reg_q2056 AND symb_decoder(16#e2#)) OR
 					(reg_q2056 AND symb_decoder(16#57#)) OR
 					(reg_q2056 AND symb_decoder(16#55#)) OR
 					(reg_q2056 AND symb_decoder(16#87#)) OR
 					(reg_q2056 AND symb_decoder(16#08#)) OR
 					(reg_q2056 AND symb_decoder(16#a7#)) OR
 					(reg_q2056 AND symb_decoder(16#59#)) OR
 					(reg_q2056 AND symb_decoder(16#93#)) OR
 					(reg_q2056 AND symb_decoder(16#7d#)) OR
 					(reg_q2056 AND symb_decoder(16#01#)) OR
 					(reg_q2056 AND symb_decoder(16#8e#)) OR
 					(reg_q2056 AND symb_decoder(16#36#)) OR
 					(reg_q2056 AND symb_decoder(16#b3#)) OR
 					(reg_q2056 AND symb_decoder(16#5b#)) OR
 					(reg_q2056 AND symb_decoder(16#33#)) OR
 					(reg_q2056 AND symb_decoder(16#b9#)) OR
 					(reg_q2056 AND symb_decoder(16#86#)) OR
 					(reg_q2056 AND symb_decoder(16#d0#)) OR
 					(reg_q2056 AND symb_decoder(16#db#)) OR
 					(reg_q2056 AND symb_decoder(16#2a#)) OR
 					(reg_q2056 AND symb_decoder(16#aa#)) OR
 					(reg_q2056 AND symb_decoder(16#e4#)) OR
 					(reg_q2056 AND symb_decoder(16#ca#)) OR
 					(reg_q2056 AND symb_decoder(16#40#)) OR
 					(reg_q2056 AND symb_decoder(16#da#)) OR
 					(reg_q2056 AND symb_decoder(16#65#)) OR
 					(reg_q2056 AND symb_decoder(16#03#)) OR
 					(reg_q2056 AND symb_decoder(16#60#)) OR
 					(reg_q2056 AND symb_decoder(16#53#)) OR
 					(reg_q2056 AND symb_decoder(16#02#)) OR
 					(reg_q2056 AND symb_decoder(16#6c#)) OR
 					(reg_q2056 AND symb_decoder(16#eb#)) OR
 					(reg_q2056 AND symb_decoder(16#f8#)) OR
 					(reg_q2056 AND symb_decoder(16#9c#)) OR
 					(reg_q2056 AND symb_decoder(16#09#)) OR
 					(reg_q2056 AND symb_decoder(16#17#)) OR
 					(reg_q2056 AND symb_decoder(16#d1#)) OR
 					(reg_q2056 AND symb_decoder(16#8b#)) OR
 					(reg_q2056 AND symb_decoder(16#7c#)) OR
 					(reg_q2056 AND symb_decoder(16#7f#)) OR
 					(reg_q2056 AND symb_decoder(16#d5#)) OR
 					(reg_q2056 AND symb_decoder(16#89#)) OR
 					(reg_q2056 AND symb_decoder(16#f1#)) OR
 					(reg_q2056 AND symb_decoder(16#bb#)) OR
 					(reg_q2056 AND symb_decoder(16#07#)) OR
 					(reg_q2056 AND symb_decoder(16#a4#)) OR
 					(reg_q2056 AND symb_decoder(16#30#)) OR
 					(reg_q2056 AND symb_decoder(16#0c#)) OR
 					(reg_q2056 AND symb_decoder(16#6d#)) OR
 					(reg_q2056 AND symb_decoder(16#c0#)) OR
 					(reg_q2056 AND symb_decoder(16#7e#)) OR
 					(reg_q2056 AND symb_decoder(16#54#)) OR
 					(reg_q2056 AND symb_decoder(16#85#)) OR
 					(reg_q2056 AND symb_decoder(16#00#)) OR
 					(reg_q2056 AND symb_decoder(16#66#)) OR
 					(reg_q2056 AND symb_decoder(16#83#)) OR
 					(reg_q2056 AND symb_decoder(16#96#)) OR
 					(reg_q2056 AND symb_decoder(16#88#)) OR
 					(reg_q2056 AND symb_decoder(16#cf#)) OR
 					(reg_q2056 AND symb_decoder(16#5d#)) OR
 					(reg_q2056 AND symb_decoder(16#16#)) OR
 					(reg_q2056 AND symb_decoder(16#6a#)) OR
 					(reg_q2056 AND symb_decoder(16#3f#)) OR
 					(reg_q2056 AND symb_decoder(16#62#)) OR
 					(reg_q2056 AND symb_decoder(16#a0#)) OR
 					(reg_q2056 AND symb_decoder(16#ac#)) OR
 					(reg_q2056 AND symb_decoder(16#71#)) OR
 					(reg_q2056 AND symb_decoder(16#c9#)) OR
 					(reg_q2056 AND symb_decoder(16#44#)) OR
 					(reg_q2056 AND symb_decoder(16#29#)) OR
 					(reg_q2056 AND symb_decoder(16#31#)) OR
 					(reg_q2056 AND symb_decoder(16#7b#)) OR
 					(reg_q2056 AND symb_decoder(16#a5#)) OR
 					(reg_q2056 AND symb_decoder(16#3c#)) OR
 					(reg_q2056 AND symb_decoder(16#f6#)) OR
 					(reg_q2056 AND symb_decoder(16#2f#)) OR
 					(reg_q2056 AND symb_decoder(16#e6#)) OR
 					(reg_q2056 AND symb_decoder(16#43#)) OR
 					(reg_q2056 AND symb_decoder(16#a8#)) OR
 					(reg_q2056 AND symb_decoder(16#c8#)) OR
 					(reg_q2056 AND symb_decoder(16#48#)) OR
 					(reg_q2056 AND symb_decoder(16#98#)) OR
 					(reg_q2056 AND symb_decoder(16#a6#)) OR
 					(reg_q2056 AND symb_decoder(16#10#)) OR
 					(reg_q2056 AND symb_decoder(16#13#)) OR
 					(reg_q2056 AND symb_decoder(16#80#)) OR
 					(reg_q2056 AND symb_decoder(16#22#)) OR
 					(reg_q2056 AND symb_decoder(16#d7#)) OR
 					(reg_q2056 AND symb_decoder(16#72#)) OR
 					(reg_q2056 AND symb_decoder(16#bf#)) OR
 					(reg_q2056 AND symb_decoder(16#ab#)) OR
 					(reg_q2056 AND symb_decoder(16#d2#)) OR
 					(reg_q2056 AND symb_decoder(16#52#)) OR
 					(reg_q2056 AND symb_decoder(16#b6#)) OR
 					(reg_q2056 AND symb_decoder(16#e7#)) OR
 					(reg_q2056 AND symb_decoder(16#8a#)) OR
 					(reg_q2056 AND symb_decoder(16#6b#)) OR
 					(reg_q2056 AND symb_decoder(16#8d#)) OR
 					(reg_q2056 AND symb_decoder(16#95#)) OR
 					(reg_q2056 AND symb_decoder(16#41#)) OR
 					(reg_q2056 AND symb_decoder(16#38#)) OR
 					(reg_q2056 AND symb_decoder(16#e5#)) OR
 					(reg_q2056 AND symb_decoder(16#25#)) OR
 					(reg_q2056 AND symb_decoder(16#4e#)) OR
 					(reg_q2056 AND symb_decoder(16#47#)) OR
 					(reg_q2056 AND symb_decoder(16#c2#)) OR
 					(reg_q2056 AND symb_decoder(16#45#)) OR
 					(reg_q2056 AND symb_decoder(16#b7#)) OR
 					(reg_q2056 AND symb_decoder(16#73#)) OR
 					(reg_q2056 AND symb_decoder(16#79#)) OR
 					(reg_q2056 AND symb_decoder(16#1f#)) OR
 					(reg_q2056 AND symb_decoder(16#d9#)) OR
 					(reg_q2056 AND symb_decoder(16#70#)) OR
 					(reg_q2056 AND symb_decoder(16#e1#)) OR
 					(reg_q2056 AND symb_decoder(16#c5#)) OR
 					(reg_q2056 AND symb_decoder(16#bc#)) OR
 					(reg_q2056 AND symb_decoder(16#c7#)) OR
 					(reg_q2056 AND symb_decoder(16#bd#)) OR
 					(reg_q2056 AND symb_decoder(16#0b#)) OR
 					(reg_q2056 AND symb_decoder(16#9b#)) OR
 					(reg_q2056 AND symb_decoder(16#2e#)) OR
 					(reg_q2056 AND symb_decoder(16#fd#)) OR
 					(reg_q2056 AND symb_decoder(16#d6#)) OR
 					(reg_q2056 AND symb_decoder(16#28#)) OR
 					(reg_q2056 AND symb_decoder(16#9e#)) OR
 					(reg_q2056 AND symb_decoder(16#12#)) OR
 					(reg_q2056 AND symb_decoder(16#df#)) OR
 					(reg_q2056 AND symb_decoder(16#b2#)) OR
 					(reg_q2056 AND symb_decoder(16#fc#)) OR
 					(reg_q2056 AND symb_decoder(16#dc#)) OR
 					(reg_q2056 AND symb_decoder(16#2b#)) OR
 					(reg_q2056 AND symb_decoder(16#99#)) OR
 					(reg_q2056 AND symb_decoder(16#a9#)) OR
 					(reg_q2056 AND symb_decoder(16#c4#)) OR
 					(reg_q2056 AND symb_decoder(16#39#)) OR
 					(reg_q2056 AND symb_decoder(16#46#)) OR
 					(reg_q2056 AND symb_decoder(16#04#)) OR
 					(reg_q2056 AND symb_decoder(16#ce#)) OR
 					(reg_q2056 AND symb_decoder(16#e8#)) OR
 					(reg_q2056 AND symb_decoder(16#3a#)) OR
 					(reg_q2056 AND symb_decoder(16#ba#)) OR
 					(reg_q2056 AND symb_decoder(16#3b#)) OR
 					(reg_q2056 AND symb_decoder(16#37#)) OR
 					(reg_q2056 AND symb_decoder(16#b8#)) OR
 					(reg_q2056 AND symb_decoder(16#cb#)) OR
 					(reg_q2056 AND symb_decoder(16#0a#)) OR
 					(reg_q2056 AND symb_decoder(16#f5#)) OR
 					(reg_q2056 AND symb_decoder(16#3e#)) OR
 					(reg_q2056 AND symb_decoder(16#ec#)) OR
 					(reg_q2056 AND symb_decoder(16#b5#)) OR
 					(reg_q2056 AND symb_decoder(16#de#)) OR
 					(reg_q2056 AND symb_decoder(16#f7#)) OR
 					(reg_q2056 AND symb_decoder(16#3d#)) OR
 					(reg_q2056 AND symb_decoder(16#56#)) OR
 					(reg_q2056 AND symb_decoder(16#5a#)) OR
 					(reg_q2056 AND symb_decoder(16#5e#)) OR
 					(reg_q2056 AND symb_decoder(16#f4#)) OR
 					(reg_q2056 AND symb_decoder(16#8f#)) OR
 					(reg_q2056 AND symb_decoder(16#ea#)) OR
 					(reg_q2056 AND symb_decoder(16#4c#)) OR
 					(reg_q2056 AND symb_decoder(16#78#)) OR
 					(reg_q2056 AND symb_decoder(16#5c#)) OR
 					(reg_q2056 AND symb_decoder(16#a2#)) OR
 					(reg_q2056 AND symb_decoder(16#e0#)) OR
 					(reg_q2056 AND symb_decoder(16#82#)) OR
 					(reg_q2056 AND symb_decoder(16#fb#)) OR
 					(reg_q2056 AND symb_decoder(16#6e#)) OR
 					(reg_q2056 AND symb_decoder(16#21#)) OR
 					(reg_q2056 AND symb_decoder(16#2d#)) OR
 					(reg_q2056 AND symb_decoder(16#81#)) OR
 					(reg_q2056 AND symb_decoder(16#5f#)) OR
 					(reg_q2056 AND symb_decoder(16#06#)) OR
 					(reg_q2056 AND symb_decoder(16#11#)) OR
 					(reg_q2056 AND symb_decoder(16#0f#)) OR
 					(reg_q2056 AND symb_decoder(16#cd#)) OR
 					(reg_q2056 AND symb_decoder(16#0e#)) OR
 					(reg_q2056 AND symb_decoder(16#74#)) OR
 					(reg_q2056 AND symb_decoder(16#97#)) OR
 					(reg_q2056 AND symb_decoder(16#58#)) OR
 					(reg_q2056 AND symb_decoder(16#4a#)) OR
 					(reg_q2056 AND symb_decoder(16#8c#)) OR
 					(reg_q2056 AND symb_decoder(16#1b#)) OR
 					(reg_q2056 AND symb_decoder(16#1d#)) OR
 					(reg_q2056 AND symb_decoder(16#76#)) OR
 					(reg_q2056 AND symb_decoder(16#a3#)) OR
 					(reg_q2056 AND symb_decoder(16#61#)) OR
 					(reg_q2056 AND symb_decoder(16#9a#)) OR
 					(reg_q2056 AND symb_decoder(16#9d#)) OR
 					(reg_q2056 AND symb_decoder(16#77#)) OR
 					(reg_q2056 AND symb_decoder(16#15#)) OR
 					(reg_q2056 AND symb_decoder(16#20#)) OR
 					(reg_q2056 AND symb_decoder(16#27#)) OR
 					(reg_q2056 AND symb_decoder(16#32#)) OR
 					(reg_q2056 AND symb_decoder(16#75#)) OR
 					(reg_q2056 AND symb_decoder(16#c6#)) OR
 					(reg_q2056 AND symb_decoder(16#67#)) OR
 					(reg_q2056 AND symb_decoder(16#18#)) OR
 					(reg_q2056 AND symb_decoder(16#ed#)) OR
 					(reg_q2056 AND symb_decoder(16#68#)) OR
 					(reg_q2056 AND symb_decoder(16#05#)) OR
 					(reg_q2056 AND symb_decoder(16#e9#)) OR
 					(reg_q2056 AND symb_decoder(16#f0#)) OR
 					(reg_q2056 AND symb_decoder(16#ee#)) OR
 					(reg_q2056 AND symb_decoder(16#b4#)) OR
 					(reg_q2056 AND symb_decoder(16#be#)) OR
 					(reg_q2056 AND symb_decoder(16#2c#)) OR
 					(reg_q2056 AND symb_decoder(16#b1#)) OR
 					(reg_q2056 AND symb_decoder(16#69#)) OR
 					(reg_q2056 AND symb_decoder(16#0d#)) OR
 					(reg_q2056 AND symb_decoder(16#4f#)) OR
 					(reg_q2056 AND symb_decoder(16#ad#)) OR
 					(reg_q2056 AND symb_decoder(16#d3#)) OR
 					(reg_q2056 AND symb_decoder(16#9f#)) OR
 					(reg_q2056 AND symb_decoder(16#4d#)) OR
 					(reg_q2056 AND symb_decoder(16#af#)) OR
 					(reg_q2056 AND symb_decoder(16#94#)) OR
 					(reg_q2056 AND symb_decoder(16#90#)) OR
 					(reg_q2056 AND symb_decoder(16#1e#)) OR
 					(reg_q2056 AND symb_decoder(16#f2#)) OR
 					(reg_q2056 AND symb_decoder(16#ae#)) OR
 					(reg_q2056 AND symb_decoder(16#50#)) OR
 					(reg_q2056 AND symb_decoder(16#d8#)) OR
 					(reg_q2056 AND symb_decoder(16#d4#)) OR
 					(reg_q2056 AND symb_decoder(16#b0#)) OR
 					(reg_q2056 AND symb_decoder(16#fa#)) OR
 					(reg_q2056 AND symb_decoder(16#fe#)) OR
 					(reg_q2056 AND symb_decoder(16#19#)) OR
 					(reg_q2056 AND symb_decoder(16#ff#)) OR
 					(reg_q2056 AND symb_decoder(16#84#)) OR
 					(reg_q2056 AND symb_decoder(16#49#)) OR
 					(reg_q2056 AND symb_decoder(16#26#)) OR
 					(reg_q2056 AND symb_decoder(16#7a#)) OR
 					(reg_q2056 AND symb_decoder(16#42#)) OR
 					(reg_q2056 AND symb_decoder(16#63#)) OR
 					(reg_q2056 AND symb_decoder(16#1a#)) OR
 					(reg_q2056 AND symb_decoder(16#35#)) OR
 					(reg_q2056 AND symb_decoder(16#14#)) OR
 					(reg_q2056 AND symb_decoder(16#92#)) OR
 					(reg_q2056 AND symb_decoder(16#c3#)) OR
 					(reg_q2056 AND symb_decoder(16#51#)) OR
 					(reg_q2056 AND symb_decoder(16#64#)) OR
 					(reg_q2056 AND symb_decoder(16#ef#)) OR
 					(reg_q2056 AND symb_decoder(16#23#)) OR
 					(reg_q2056 AND symb_decoder(16#4b#)) OR
 					(reg_q2056 AND symb_decoder(16#6f#)) OR
 					(reg_q2056 AND symb_decoder(16#c1#)) OR
 					(reg_q2056 AND symb_decoder(16#a1#)) OR
 					(reg_q2056 AND symb_decoder(16#cc#)) OR
 					(reg_q2056 AND symb_decoder(16#1c#));
reg_q2056_init <= '0' ;
	p_reg_q2056: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2056 <= reg_q2056_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2056 <= reg_q2056_init;
        else
          reg_q2056 <= reg_q2056_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1393_in <= (reg_q1393 AND symb_decoder(16#72#)) OR
 					(reg_q1393 AND symb_decoder(16#94#)) OR
 					(reg_q1393 AND symb_decoder(16#43#)) OR
 					(reg_q1393 AND symb_decoder(16#4e#)) OR
 					(reg_q1393 AND symb_decoder(16#9c#)) OR
 					(reg_q1393 AND symb_decoder(16#dc#)) OR
 					(reg_q1393 AND symb_decoder(16#58#)) OR
 					(reg_q1393 AND symb_decoder(16#1c#)) OR
 					(reg_q1393 AND symb_decoder(16#2c#)) OR
 					(reg_q1393 AND symb_decoder(16#a7#)) OR
 					(reg_q1393 AND symb_decoder(16#d4#)) OR
 					(reg_q1393 AND symb_decoder(16#1b#)) OR
 					(reg_q1393 AND symb_decoder(16#fa#)) OR
 					(reg_q1393 AND symb_decoder(16#7c#)) OR
 					(reg_q1393 AND symb_decoder(16#91#)) OR
 					(reg_q1393 AND symb_decoder(16#61#)) OR
 					(reg_q1393 AND symb_decoder(16#a9#)) OR
 					(reg_q1393 AND symb_decoder(16#15#)) OR
 					(reg_q1393 AND symb_decoder(16#fb#)) OR
 					(reg_q1393 AND symb_decoder(16#b7#)) OR
 					(reg_q1393 AND symb_decoder(16#53#)) OR
 					(reg_q1393 AND symb_decoder(16#ca#)) OR
 					(reg_q1393 AND symb_decoder(16#c5#)) OR
 					(reg_q1393 AND symb_decoder(16#87#)) OR
 					(reg_q1393 AND symb_decoder(16#56#)) OR
 					(reg_q1393 AND symb_decoder(16#ae#)) OR
 					(reg_q1393 AND symb_decoder(16#f5#)) OR
 					(reg_q1393 AND symb_decoder(16#f3#)) OR
 					(reg_q1393 AND symb_decoder(16#b2#)) OR
 					(reg_q1393 AND symb_decoder(16#0c#)) OR
 					(reg_q1393 AND symb_decoder(16#06#)) OR
 					(reg_q1393 AND symb_decoder(16#ee#)) OR
 					(reg_q1393 AND symb_decoder(16#c9#)) OR
 					(reg_q1393 AND symb_decoder(16#ba#)) OR
 					(reg_q1393 AND symb_decoder(16#af#)) OR
 					(reg_q1393 AND symb_decoder(16#ea#)) OR
 					(reg_q1393 AND symb_decoder(16#aa#)) OR
 					(reg_q1393 AND symb_decoder(16#d3#)) OR
 					(reg_q1393 AND symb_decoder(16#64#)) OR
 					(reg_q1393 AND symb_decoder(16#5f#)) OR
 					(reg_q1393 AND symb_decoder(16#a6#)) OR
 					(reg_q1393 AND symb_decoder(16#8a#)) OR
 					(reg_q1393 AND symb_decoder(16#ff#)) OR
 					(reg_q1393 AND symb_decoder(16#62#)) OR
 					(reg_q1393 AND symb_decoder(16#66#)) OR
 					(reg_q1393 AND symb_decoder(16#03#)) OR
 					(reg_q1393 AND symb_decoder(16#00#)) OR
 					(reg_q1393 AND symb_decoder(16#96#)) OR
 					(reg_q1393 AND symb_decoder(16#31#)) OR
 					(reg_q1393 AND symb_decoder(16#11#)) OR
 					(reg_q1393 AND symb_decoder(16#73#)) OR
 					(reg_q1393 AND symb_decoder(16#0e#)) OR
 					(reg_q1393 AND symb_decoder(16#f0#)) OR
 					(reg_q1393 AND symb_decoder(16#89#)) OR
 					(reg_q1393 AND symb_decoder(16#17#)) OR
 					(reg_q1393 AND symb_decoder(16#7f#)) OR
 					(reg_q1393 AND symb_decoder(16#ad#)) OR
 					(reg_q1393 AND symb_decoder(16#7b#)) OR
 					(reg_q1393 AND symb_decoder(16#be#)) OR
 					(reg_q1393 AND symb_decoder(16#0d#)) OR
 					(reg_q1393 AND symb_decoder(16#c6#)) OR
 					(reg_q1393 AND symb_decoder(16#d2#)) OR
 					(reg_q1393 AND symb_decoder(16#09#)) OR
 					(reg_q1393 AND symb_decoder(16#71#)) OR
 					(reg_q1393 AND symb_decoder(16#6a#)) OR
 					(reg_q1393 AND symb_decoder(16#d8#)) OR
 					(reg_q1393 AND symb_decoder(16#78#)) OR
 					(reg_q1393 AND symb_decoder(16#8c#)) OR
 					(reg_q1393 AND symb_decoder(16#84#)) OR
 					(reg_q1393 AND symb_decoder(16#1d#)) OR
 					(reg_q1393 AND symb_decoder(16#dd#)) OR
 					(reg_q1393 AND symb_decoder(16#db#)) OR
 					(reg_q1393 AND symb_decoder(16#c3#)) OR
 					(reg_q1393 AND symb_decoder(16#93#)) OR
 					(reg_q1393 AND symb_decoder(16#47#)) OR
 					(reg_q1393 AND symb_decoder(16#f2#)) OR
 					(reg_q1393 AND symb_decoder(16#cf#)) OR
 					(reg_q1393 AND symb_decoder(16#30#)) OR
 					(reg_q1393 AND symb_decoder(16#e5#)) OR
 					(reg_q1393 AND symb_decoder(16#69#)) OR
 					(reg_q1393 AND symb_decoder(16#27#)) OR
 					(reg_q1393 AND symb_decoder(16#44#)) OR
 					(reg_q1393 AND symb_decoder(16#a8#)) OR
 					(reg_q1393 AND symb_decoder(16#2a#)) OR
 					(reg_q1393 AND symb_decoder(16#98#)) OR
 					(reg_q1393 AND symb_decoder(16#48#)) OR
 					(reg_q1393 AND symb_decoder(16#05#)) OR
 					(reg_q1393 AND symb_decoder(16#20#)) OR
 					(reg_q1393 AND symb_decoder(16#a4#)) OR
 					(reg_q1393 AND symb_decoder(16#33#)) OR
 					(reg_q1393 AND symb_decoder(16#70#)) OR
 					(reg_q1393 AND symb_decoder(16#60#)) OR
 					(reg_q1393 AND symb_decoder(16#6f#)) OR
 					(reg_q1393 AND symb_decoder(16#28#)) OR
 					(reg_q1393 AND symb_decoder(16#55#)) OR
 					(reg_q1393 AND symb_decoder(16#b3#)) OR
 					(reg_q1393 AND symb_decoder(16#99#)) OR
 					(reg_q1393 AND symb_decoder(16#81#)) OR
 					(reg_q1393 AND symb_decoder(16#3c#)) OR
 					(reg_q1393 AND symb_decoder(16#7d#)) OR
 					(reg_q1393 AND symb_decoder(16#df#)) OR
 					(reg_q1393 AND symb_decoder(16#51#)) OR
 					(reg_q1393 AND symb_decoder(16#b5#)) OR
 					(reg_q1393 AND symb_decoder(16#3e#)) OR
 					(reg_q1393 AND symb_decoder(16#83#)) OR
 					(reg_q1393 AND symb_decoder(16#3a#)) OR
 					(reg_q1393 AND symb_decoder(16#76#)) OR
 					(reg_q1393 AND symb_decoder(16#b1#)) OR
 					(reg_q1393 AND symb_decoder(16#92#)) OR
 					(reg_q1393 AND symb_decoder(16#22#)) OR
 					(reg_q1393 AND symb_decoder(16#90#)) OR
 					(reg_q1393 AND symb_decoder(16#50#)) OR
 					(reg_q1393 AND symb_decoder(16#57#)) OR
 					(reg_q1393 AND symb_decoder(16#da#)) OR
 					(reg_q1393 AND symb_decoder(16#02#)) OR
 					(reg_q1393 AND symb_decoder(16#e2#)) OR
 					(reg_q1393 AND symb_decoder(16#a1#)) OR
 					(reg_q1393 AND symb_decoder(16#d9#)) OR
 					(reg_q1393 AND symb_decoder(16#e3#)) OR
 					(reg_q1393 AND symb_decoder(16#d6#)) OR
 					(reg_q1393 AND symb_decoder(16#32#)) OR
 					(reg_q1393 AND symb_decoder(16#42#)) OR
 					(reg_q1393 AND symb_decoder(16#a3#)) OR
 					(reg_q1393 AND symb_decoder(16#37#)) OR
 					(reg_q1393 AND symb_decoder(16#80#)) OR
 					(reg_q1393 AND symb_decoder(16#e8#)) OR
 					(reg_q1393 AND symb_decoder(16#7a#)) OR
 					(reg_q1393 AND symb_decoder(16#b8#)) OR
 					(reg_q1393 AND symb_decoder(16#cc#)) OR
 					(reg_q1393 AND symb_decoder(16#e1#)) OR
 					(reg_q1393 AND symb_decoder(16#8b#)) OR
 					(reg_q1393 AND symb_decoder(16#ec#)) OR
 					(reg_q1393 AND symb_decoder(16#5a#)) OR
 					(reg_q1393 AND symb_decoder(16#c7#)) OR
 					(reg_q1393 AND symb_decoder(16#35#)) OR
 					(reg_q1393 AND symb_decoder(16#5b#)) OR
 					(reg_q1393 AND symb_decoder(16#9d#)) OR
 					(reg_q1393 AND symb_decoder(16#4a#)) OR
 					(reg_q1393 AND symb_decoder(16#9f#)) OR
 					(reg_q1393 AND symb_decoder(16#ab#)) OR
 					(reg_q1393 AND symb_decoder(16#5c#)) OR
 					(reg_q1393 AND symb_decoder(16#ed#)) OR
 					(reg_q1393 AND symb_decoder(16#75#)) OR
 					(reg_q1393 AND symb_decoder(16#65#)) OR
 					(reg_q1393 AND symb_decoder(16#79#)) OR
 					(reg_q1393 AND symb_decoder(16#f1#)) OR
 					(reg_q1393 AND symb_decoder(16#8d#)) OR
 					(reg_q1393 AND symb_decoder(16#b6#)) OR
 					(reg_q1393 AND symb_decoder(16#8e#)) OR
 					(reg_q1393 AND symb_decoder(16#21#)) OR
 					(reg_q1393 AND symb_decoder(16#12#)) OR
 					(reg_q1393 AND symb_decoder(16#36#)) OR
 					(reg_q1393 AND symb_decoder(16#3f#)) OR
 					(reg_q1393 AND symb_decoder(16#f9#)) OR
 					(reg_q1393 AND symb_decoder(16#16#)) OR
 					(reg_q1393 AND symb_decoder(16#a0#)) OR
 					(reg_q1393 AND symb_decoder(16#0b#)) OR
 					(reg_q1393 AND symb_decoder(16#82#)) OR
 					(reg_q1393 AND symb_decoder(16#0f#)) OR
 					(reg_q1393 AND symb_decoder(16#2b#)) OR
 					(reg_q1393 AND symb_decoder(16#e4#)) OR
 					(reg_q1393 AND symb_decoder(16#de#)) OR
 					(reg_q1393 AND symb_decoder(16#5d#)) OR
 					(reg_q1393 AND symb_decoder(16#39#)) OR
 					(reg_q1393 AND symb_decoder(16#85#)) OR
 					(reg_q1393 AND symb_decoder(16#13#)) OR
 					(reg_q1393 AND symb_decoder(16#fc#)) OR
 					(reg_q1393 AND symb_decoder(16#18#)) OR
 					(reg_q1393 AND symb_decoder(16#ef#)) OR
 					(reg_q1393 AND symb_decoder(16#29#)) OR
 					(reg_q1393 AND symb_decoder(16#59#)) OR
 					(reg_q1393 AND symb_decoder(16#c4#)) OR
 					(reg_q1393 AND symb_decoder(16#d5#)) OR
 					(reg_q1393 AND symb_decoder(16#1f#)) OR
 					(reg_q1393 AND symb_decoder(16#cb#)) OR
 					(reg_q1393 AND symb_decoder(16#cd#)) OR
 					(reg_q1393 AND symb_decoder(16#e0#)) OR
 					(reg_q1393 AND symb_decoder(16#bc#)) OR
 					(reg_q1393 AND symb_decoder(16#74#)) OR
 					(reg_q1393 AND symb_decoder(16#40#)) OR
 					(reg_q1393 AND symb_decoder(16#a2#)) OR
 					(reg_q1393 AND symb_decoder(16#46#)) OR
 					(reg_q1393 AND symb_decoder(16#24#)) OR
 					(reg_q1393 AND symb_decoder(16#7e#)) OR
 					(reg_q1393 AND symb_decoder(16#bd#)) OR
 					(reg_q1393 AND symb_decoder(16#e9#)) OR
 					(reg_q1393 AND symb_decoder(16#77#)) OR
 					(reg_q1393 AND symb_decoder(16#38#)) OR
 					(reg_q1393 AND symb_decoder(16#68#)) OR
 					(reg_q1393 AND symb_decoder(16#bf#)) OR
 					(reg_q1393 AND symb_decoder(16#45#)) OR
 					(reg_q1393 AND symb_decoder(16#2e#)) OR
 					(reg_q1393 AND symb_decoder(16#8f#)) OR
 					(reg_q1393 AND symb_decoder(16#c8#)) OR
 					(reg_q1393 AND symb_decoder(16#08#)) OR
 					(reg_q1393 AND symb_decoder(16#c1#)) OR
 					(reg_q1393 AND symb_decoder(16#34#)) OR
 					(reg_q1393 AND symb_decoder(16#b9#)) OR
 					(reg_q1393 AND symb_decoder(16#1a#)) OR
 					(reg_q1393 AND symb_decoder(16#23#)) OR
 					(reg_q1393 AND symb_decoder(16#6d#)) OR
 					(reg_q1393 AND symb_decoder(16#63#)) OR
 					(reg_q1393 AND symb_decoder(16#9e#)) OR
 					(reg_q1393 AND symb_decoder(16#9b#)) OR
 					(reg_q1393 AND symb_decoder(16#f7#)) OR
 					(reg_q1393 AND symb_decoder(16#4b#)) OR
 					(reg_q1393 AND symb_decoder(16#04#)) OR
 					(reg_q1393 AND symb_decoder(16#d1#)) OR
 					(reg_q1393 AND symb_decoder(16#a5#)) OR
 					(reg_q1393 AND symb_decoder(16#95#)) OR
 					(reg_q1393 AND symb_decoder(16#fd#)) OR
 					(reg_q1393 AND symb_decoder(16#9a#)) OR
 					(reg_q1393 AND symb_decoder(16#f4#)) OR
 					(reg_q1393 AND symb_decoder(16#41#)) OR
 					(reg_q1393 AND symb_decoder(16#eb#)) OR
 					(reg_q1393 AND symb_decoder(16#88#)) OR
 					(reg_q1393 AND symb_decoder(16#1e#)) OR
 					(reg_q1393 AND symb_decoder(16#bb#)) OR
 					(reg_q1393 AND symb_decoder(16#d0#)) OR
 					(reg_q1393 AND symb_decoder(16#6e#)) OR
 					(reg_q1393 AND symb_decoder(16#10#)) OR
 					(reg_q1393 AND symb_decoder(16#25#)) OR
 					(reg_q1393 AND symb_decoder(16#2f#)) OR
 					(reg_q1393 AND symb_decoder(16#ce#)) OR
 					(reg_q1393 AND symb_decoder(16#c2#)) OR
 					(reg_q1393 AND symb_decoder(16#3b#)) OR
 					(reg_q1393 AND symb_decoder(16#67#)) OR
 					(reg_q1393 AND symb_decoder(16#14#)) OR
 					(reg_q1393 AND symb_decoder(16#4d#)) OR
 					(reg_q1393 AND symb_decoder(16#86#)) OR
 					(reg_q1393 AND symb_decoder(16#0a#)) OR
 					(reg_q1393 AND symb_decoder(16#f6#)) OR
 					(reg_q1393 AND symb_decoder(16#e6#)) OR
 					(reg_q1393 AND symb_decoder(16#e7#)) OR
 					(reg_q1393 AND symb_decoder(16#49#)) OR
 					(reg_q1393 AND symb_decoder(16#2d#)) OR
 					(reg_q1393 AND symb_decoder(16#ac#)) OR
 					(reg_q1393 AND symb_decoder(16#4c#)) OR
 					(reg_q1393 AND symb_decoder(16#6b#)) OR
 					(reg_q1393 AND symb_decoder(16#54#)) OR
 					(reg_q1393 AND symb_decoder(16#f8#)) OR
 					(reg_q1393 AND symb_decoder(16#52#)) OR
 					(reg_q1393 AND symb_decoder(16#26#)) OR
 					(reg_q1393 AND symb_decoder(16#4f#)) OR
 					(reg_q1393 AND symb_decoder(16#c0#)) OR
 					(reg_q1393 AND symb_decoder(16#19#)) OR
 					(reg_q1393 AND symb_decoder(16#b0#)) OR
 					(reg_q1393 AND symb_decoder(16#07#)) OR
 					(reg_q1393 AND symb_decoder(16#5e#)) OR
 					(reg_q1393 AND symb_decoder(16#6c#)) OR
 					(reg_q1393 AND symb_decoder(16#b4#)) OR
 					(reg_q1393 AND symb_decoder(16#01#)) OR
 					(reg_q1393 AND symb_decoder(16#3d#)) OR
 					(reg_q1393 AND symb_decoder(16#fe#)) OR
 					(reg_q1393 AND symb_decoder(16#d7#)) OR
 					(reg_q1393 AND symb_decoder(16#97#)) OR
 					(reg_q1357 AND symb_decoder(16#78#)) OR
 					(reg_q1357 AND symb_decoder(16#41#)) OR
 					(reg_q1357 AND symb_decoder(16#36#)) OR
 					(reg_q1357 AND symb_decoder(16#c4#)) OR
 					(reg_q1357 AND symb_decoder(16#a1#)) OR
 					(reg_q1357 AND symb_decoder(16#ed#)) OR
 					(reg_q1357 AND symb_decoder(16#d3#)) OR
 					(reg_q1357 AND symb_decoder(16#07#)) OR
 					(reg_q1357 AND symb_decoder(16#b1#)) OR
 					(reg_q1357 AND symb_decoder(16#7b#)) OR
 					(reg_q1357 AND symb_decoder(16#d1#)) OR
 					(reg_q1357 AND symb_decoder(16#7d#)) OR
 					(reg_q1357 AND symb_decoder(16#93#)) OR
 					(reg_q1357 AND symb_decoder(16#50#)) OR
 					(reg_q1357 AND symb_decoder(16#10#)) OR
 					(reg_q1357 AND symb_decoder(16#82#)) OR
 					(reg_q1357 AND symb_decoder(16#8e#)) OR
 					(reg_q1357 AND symb_decoder(16#8f#)) OR
 					(reg_q1357 AND symb_decoder(16#86#)) OR
 					(reg_q1357 AND symb_decoder(16#89#)) OR
 					(reg_q1357 AND symb_decoder(16#72#)) OR
 					(reg_q1357 AND symb_decoder(16#13#)) OR
 					(reg_q1357 AND symb_decoder(16#bb#)) OR
 					(reg_q1357 AND symb_decoder(16#f2#)) OR
 					(reg_q1357 AND symb_decoder(16#c2#)) OR
 					(reg_q1357 AND symb_decoder(16#e1#)) OR
 					(reg_q1357 AND symb_decoder(16#96#)) OR
 					(reg_q1357 AND symb_decoder(16#2f#)) OR
 					(reg_q1357 AND symb_decoder(16#f4#)) OR
 					(reg_q1357 AND symb_decoder(16#47#)) OR
 					(reg_q1357 AND symb_decoder(16#46#)) OR
 					(reg_q1357 AND symb_decoder(16#3a#)) OR
 					(reg_q1357 AND symb_decoder(16#24#)) OR
 					(reg_q1357 AND symb_decoder(16#69#)) OR
 					(reg_q1357 AND symb_decoder(16#d6#)) OR
 					(reg_q1357 AND symb_decoder(16#6d#)) OR
 					(reg_q1357 AND symb_decoder(16#45#)) OR
 					(reg_q1357 AND symb_decoder(16#ec#)) OR
 					(reg_q1357 AND symb_decoder(16#e5#)) OR
 					(reg_q1357 AND symb_decoder(16#d4#)) OR
 					(reg_q1357 AND symb_decoder(16#8c#)) OR
 					(reg_q1357 AND symb_decoder(16#0c#)) OR
 					(reg_q1357 AND symb_decoder(16#1a#)) OR
 					(reg_q1357 AND symb_decoder(16#c1#)) OR
 					(reg_q1357 AND symb_decoder(16#a5#)) OR
 					(reg_q1357 AND symb_decoder(16#34#)) OR
 					(reg_q1357 AND symb_decoder(16#20#)) OR
 					(reg_q1357 AND symb_decoder(16#7a#)) OR
 					(reg_q1357 AND symb_decoder(16#8a#)) OR
 					(reg_q1357 AND symb_decoder(16#76#)) OR
 					(reg_q1357 AND symb_decoder(16#62#)) OR
 					(reg_q1357 AND symb_decoder(16#71#)) OR
 					(reg_q1357 AND symb_decoder(16#68#)) OR
 					(reg_q1357 AND symb_decoder(16#a9#)) OR
 					(reg_q1357 AND symb_decoder(16#2c#)) OR
 					(reg_q1357 AND symb_decoder(16#f1#)) OR
 					(reg_q1357 AND symb_decoder(16#a0#)) OR
 					(reg_q1357 AND symb_decoder(16#2a#)) OR
 					(reg_q1357 AND symb_decoder(16#35#)) OR
 					(reg_q1357 AND symb_decoder(16#6b#)) OR
 					(reg_q1357 AND symb_decoder(16#a8#)) OR
 					(reg_q1357 AND symb_decoder(16#4b#)) OR
 					(reg_q1357 AND symb_decoder(16#b2#)) OR
 					(reg_q1357 AND symb_decoder(16#d0#)) OR
 					(reg_q1357 AND symb_decoder(16#9f#)) OR
 					(reg_q1357 AND symb_decoder(16#6c#)) OR
 					(reg_q1357 AND symb_decoder(16#cc#)) OR
 					(reg_q1357 AND symb_decoder(16#9a#)) OR
 					(reg_q1357 AND symb_decoder(16#dd#)) OR
 					(reg_q1357 AND symb_decoder(16#30#)) OR
 					(reg_q1357 AND symb_decoder(16#da#)) OR
 					(reg_q1357 AND symb_decoder(16#7c#)) OR
 					(reg_q1357 AND symb_decoder(16#f9#)) OR
 					(reg_q1357 AND symb_decoder(16#09#)) OR
 					(reg_q1357 AND symb_decoder(16#26#)) OR
 					(reg_q1357 AND symb_decoder(16#3c#)) OR
 					(reg_q1357 AND symb_decoder(16#b5#)) OR
 					(reg_q1357 AND symb_decoder(16#18#)) OR
 					(reg_q1357 AND symb_decoder(16#e6#)) OR
 					(reg_q1357 AND symb_decoder(16#81#)) OR
 					(reg_q1357 AND symb_decoder(16#cf#)) OR
 					(reg_q1357 AND symb_decoder(16#91#)) OR
 					(reg_q1357 AND symb_decoder(16#a7#)) OR
 					(reg_q1357 AND symb_decoder(16#5b#)) OR
 					(reg_q1357 AND symb_decoder(16#c9#)) OR
 					(reg_q1357 AND symb_decoder(16#b6#)) OR
 					(reg_q1357 AND symb_decoder(16#23#)) OR
 					(reg_q1357 AND symb_decoder(16#6f#)) OR
 					(reg_q1357 AND symb_decoder(16#e4#)) OR
 					(reg_q1357 AND symb_decoder(16#f0#)) OR
 					(reg_q1357 AND symb_decoder(16#ff#)) OR
 					(reg_q1357 AND symb_decoder(16#33#)) OR
 					(reg_q1357 AND symb_decoder(16#d9#)) OR
 					(reg_q1357 AND symb_decoder(16#61#)) OR
 					(reg_q1357 AND symb_decoder(16#51#)) OR
 					(reg_q1357 AND symb_decoder(16#2d#)) OR
 					(reg_q1357 AND symb_decoder(16#39#)) OR
 					(reg_q1357 AND symb_decoder(16#75#)) OR
 					(reg_q1357 AND symb_decoder(16#1e#)) OR
 					(reg_q1357 AND symb_decoder(16#44#)) OR
 					(reg_q1357 AND symb_decoder(16#83#)) OR
 					(reg_q1357 AND symb_decoder(16#f8#)) OR
 					(reg_q1357 AND symb_decoder(16#54#)) OR
 					(reg_q1357 AND symb_decoder(16#a2#)) OR
 					(reg_q1357 AND symb_decoder(16#48#)) OR
 					(reg_q1357 AND symb_decoder(16#5a#)) OR
 					(reg_q1357 AND symb_decoder(16#5f#)) OR
 					(reg_q1357 AND symb_decoder(16#0a#)) OR
 					(reg_q1357 AND symb_decoder(16#3b#)) OR
 					(reg_q1357 AND symb_decoder(16#03#)) OR
 					(reg_q1357 AND symb_decoder(16#7e#)) OR
 					(reg_q1357 AND symb_decoder(16#6a#)) OR
 					(reg_q1357 AND symb_decoder(16#65#)) OR
 					(reg_q1357 AND symb_decoder(16#3e#)) OR
 					(reg_q1357 AND symb_decoder(16#f3#)) OR
 					(reg_q1357 AND symb_decoder(16#cd#)) OR
 					(reg_q1357 AND symb_decoder(16#e7#)) OR
 					(reg_q1357 AND symb_decoder(16#57#)) OR
 					(reg_q1357 AND symb_decoder(16#d2#)) OR
 					(reg_q1357 AND symb_decoder(16#aa#)) OR
 					(reg_q1357 AND symb_decoder(16#08#)) OR
 					(reg_q1357 AND symb_decoder(16#0b#)) OR
 					(reg_q1357 AND symb_decoder(16#59#)) OR
 					(reg_q1357 AND symb_decoder(16#ad#)) OR
 					(reg_q1357 AND symb_decoder(16#0f#)) OR
 					(reg_q1357 AND symb_decoder(16#be#)) OR
 					(reg_q1357 AND symb_decoder(16#64#)) OR
 					(reg_q1357 AND symb_decoder(16#87#)) OR
 					(reg_q1357 AND symb_decoder(16#db#)) OR
 					(reg_q1357 AND symb_decoder(16#97#)) OR
 					(reg_q1357 AND symb_decoder(16#a4#)) OR
 					(reg_q1357 AND symb_decoder(16#6e#)) OR
 					(reg_q1357 AND symb_decoder(16#05#)) OR
 					(reg_q1357 AND symb_decoder(16#84#)) OR
 					(reg_q1357 AND symb_decoder(16#19#)) OR
 					(reg_q1357 AND symb_decoder(16#37#)) OR
 					(reg_q1357 AND symb_decoder(16#29#)) OR
 					(reg_q1357 AND symb_decoder(16#9c#)) OR
 					(reg_q1357 AND symb_decoder(16#15#)) OR
 					(reg_q1357 AND symb_decoder(16#17#)) OR
 					(reg_q1357 AND symb_decoder(16#fa#)) OR
 					(reg_q1357 AND symb_decoder(16#8d#)) OR
 					(reg_q1357 AND symb_decoder(16#60#)) OR
 					(reg_q1357 AND symb_decoder(16#02#)) OR
 					(reg_q1357 AND symb_decoder(16#eb#)) OR
 					(reg_q1357 AND symb_decoder(16#ab#)) OR
 					(reg_q1357 AND symb_decoder(16#4c#)) OR
 					(reg_q1357 AND symb_decoder(16#92#)) OR
 					(reg_q1357 AND symb_decoder(16#e8#)) OR
 					(reg_q1357 AND symb_decoder(16#42#)) OR
 					(reg_q1357 AND symb_decoder(16#66#)) OR
 					(reg_q1357 AND symb_decoder(16#5e#)) OR
 					(reg_q1357 AND symb_decoder(16#e0#)) OR
 					(reg_q1357 AND symb_decoder(16#a3#)) OR
 					(reg_q1357 AND symb_decoder(16#1f#)) OR
 					(reg_q1357 AND symb_decoder(16#1b#)) OR
 					(reg_q1357 AND symb_decoder(16#ae#)) OR
 					(reg_q1357 AND symb_decoder(16#0d#)) OR
 					(reg_q1357 AND symb_decoder(16#dc#)) OR
 					(reg_q1357 AND symb_decoder(16#ce#)) OR
 					(reg_q1357 AND symb_decoder(16#d7#)) OR
 					(reg_q1357 AND symb_decoder(16#28#)) OR
 					(reg_q1357 AND symb_decoder(16#ee#)) OR
 					(reg_q1357 AND symb_decoder(16#52#)) OR
 					(reg_q1357 AND symb_decoder(16#af#)) OR
 					(reg_q1357 AND symb_decoder(16#63#)) OR
 					(reg_q1357 AND symb_decoder(16#c8#)) OR
 					(reg_q1357 AND symb_decoder(16#4d#)) OR
 					(reg_q1357 AND symb_decoder(16#4a#)) OR
 					(reg_q1357 AND symb_decoder(16#3d#)) OR
 					(reg_q1357 AND symb_decoder(16#ca#)) OR
 					(reg_q1357 AND symb_decoder(16#73#)) OR
 					(reg_q1357 AND symb_decoder(16#f6#)) OR
 					(reg_q1357 AND symb_decoder(16#04#)) OR
 					(reg_q1357 AND symb_decoder(16#c6#)) OR
 					(reg_q1357 AND symb_decoder(16#14#)) OR
 					(reg_q1357 AND symb_decoder(16#2b#)) OR
 					(reg_q1357 AND symb_decoder(16#de#)) OR
 					(reg_q1357 AND symb_decoder(16#31#)) OR
 					(reg_q1357 AND symb_decoder(16#95#)) OR
 					(reg_q1357 AND symb_decoder(16#01#)) OR
 					(reg_q1357 AND symb_decoder(16#a6#)) OR
 					(reg_q1357 AND symb_decoder(16#b3#)) OR
 					(reg_q1357 AND symb_decoder(16#4f#)) OR
 					(reg_q1357 AND symb_decoder(16#85#)) OR
 					(reg_q1357 AND symb_decoder(16#fd#)) OR
 					(reg_q1357 AND symb_decoder(16#c7#)) OR
 					(reg_q1357 AND symb_decoder(16#bf#)) OR
 					(reg_q1357 AND symb_decoder(16#74#)) OR
 					(reg_q1357 AND symb_decoder(16#4e#)) OR
 					(reg_q1357 AND symb_decoder(16#58#)) OR
 					(reg_q1357 AND symb_decoder(16#06#)) OR
 					(reg_q1357 AND symb_decoder(16#5c#)) OR
 					(reg_q1357 AND symb_decoder(16#f7#)) OR
 					(reg_q1357 AND symb_decoder(16#bd#)) OR
 					(reg_q1357 AND symb_decoder(16#22#)) OR
 					(reg_q1357 AND symb_decoder(16#1c#)) OR
 					(reg_q1357 AND symb_decoder(16#98#)) OR
 					(reg_q1357 AND symb_decoder(16#2e#)) OR
 					(reg_q1357 AND symb_decoder(16#27#)) OR
 					(reg_q1357 AND symb_decoder(16#ea#)) OR
 					(reg_q1357 AND symb_decoder(16#3f#)) OR
 					(reg_q1357 AND symb_decoder(16#53#)) OR
 					(reg_q1357 AND symb_decoder(16#32#)) OR
 					(reg_q1357 AND symb_decoder(16#fc#)) OR
 					(reg_q1357 AND symb_decoder(16#ef#)) OR
 					(reg_q1357 AND symb_decoder(16#67#)) OR
 					(reg_q1357 AND symb_decoder(16#b4#)) OR
 					(reg_q1357 AND symb_decoder(16#55#)) OR
 					(reg_q1357 AND symb_decoder(16#38#)) OR
 					(reg_q1357 AND symb_decoder(16#b8#)) OR
 					(reg_q1357 AND symb_decoder(16#0e#)) OR
 					(reg_q1357 AND symb_decoder(16#90#)) OR
 					(reg_q1357 AND symb_decoder(16#56#)) OR
 					(reg_q1357 AND symb_decoder(16#e3#)) OR
 					(reg_q1357 AND symb_decoder(16#43#)) OR
 					(reg_q1357 AND symb_decoder(16#c5#)) OR
 					(reg_q1357 AND symb_decoder(16#94#)) OR
 					(reg_q1357 AND symb_decoder(16#b0#)) OR
 					(reg_q1357 AND symb_decoder(16#9e#)) OR
 					(reg_q1357 AND symb_decoder(16#25#)) OR
 					(reg_q1357 AND symb_decoder(16#7f#)) OR
 					(reg_q1357 AND symb_decoder(16#df#)) OR
 					(reg_q1357 AND symb_decoder(16#80#)) OR
 					(reg_q1357 AND symb_decoder(16#1d#)) OR
 					(reg_q1357 AND symb_decoder(16#c3#)) OR
 					(reg_q1357 AND symb_decoder(16#9d#)) OR
 					(reg_q1357 AND symb_decoder(16#d5#)) OR
 					(reg_q1357 AND symb_decoder(16#ac#)) OR
 					(reg_q1357 AND symb_decoder(16#e9#)) OR
 					(reg_q1357 AND symb_decoder(16#fb#)) OR
 					(reg_q1357 AND symb_decoder(16#cb#)) OR
 					(reg_q1357 AND symb_decoder(16#8b#)) OR
 					(reg_q1357 AND symb_decoder(16#c0#)) OR
 					(reg_q1357 AND symb_decoder(16#e2#)) OR
 					(reg_q1357 AND symb_decoder(16#70#)) OR
 					(reg_q1357 AND symb_decoder(16#f5#)) OR
 					(reg_q1357 AND symb_decoder(16#fe#)) OR
 					(reg_q1357 AND symb_decoder(16#99#)) OR
 					(reg_q1357 AND symb_decoder(16#77#)) OR
 					(reg_q1357 AND symb_decoder(16#12#)) OR
 					(reg_q1357 AND symb_decoder(16#21#)) OR
 					(reg_q1357 AND symb_decoder(16#11#)) OR
 					(reg_q1357 AND symb_decoder(16#40#)) OR
 					(reg_q1357 AND symb_decoder(16#79#)) OR
 					(reg_q1357 AND symb_decoder(16#ba#)) OR
 					(reg_q1357 AND symb_decoder(16#b7#)) OR
 					(reg_q1357 AND symb_decoder(16#88#)) OR
 					(reg_q1357 AND symb_decoder(16#49#)) OR
 					(reg_q1357 AND symb_decoder(16#bc#)) OR
 					(reg_q1357 AND symb_decoder(16#00#)) OR
 					(reg_q1357 AND symb_decoder(16#b9#)) OR
 					(reg_q1357 AND symb_decoder(16#16#)) OR
 					(reg_q1357 AND symb_decoder(16#d8#)) OR
 					(reg_q1357 AND symb_decoder(16#5d#)) OR
 					(reg_q1357 AND symb_decoder(16#9b#));
reg_q1393_init <= '0' ;
	p_reg_q1393: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1393 <= reg_q1393_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1393 <= reg_q1393_init;
        else
          reg_q1393 <= reg_q1393_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1685_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1685 AND symb_decoder(16#7c#)) OR
 					(reg_q1685 AND symb_decoder(16#83#)) OR
 					(reg_q1685 AND symb_decoder(16#4f#)) OR
 					(reg_q1685 AND symb_decoder(16#00#)) OR
 					(reg_q1685 AND symb_decoder(16#03#)) OR
 					(reg_q1685 AND symb_decoder(16#a5#)) OR
 					(reg_q1685 AND symb_decoder(16#cb#)) OR
 					(reg_q1685 AND symb_decoder(16#6d#)) OR
 					(reg_q1685 AND symb_decoder(16#76#)) OR
 					(reg_q1685 AND symb_decoder(16#be#)) OR
 					(reg_q1685 AND symb_decoder(16#cc#)) OR
 					(reg_q1685 AND symb_decoder(16#da#)) OR
 					(reg_q1685 AND symb_decoder(16#8a#)) OR
 					(reg_q1685 AND symb_decoder(16#22#)) OR
 					(reg_q1685 AND symb_decoder(16#d5#)) OR
 					(reg_q1685 AND symb_decoder(16#df#)) OR
 					(reg_q1685 AND symb_decoder(16#eb#)) OR
 					(reg_q1685 AND symb_decoder(16#9b#)) OR
 					(reg_q1685 AND symb_decoder(16#a7#)) OR
 					(reg_q1685 AND symb_decoder(16#0d#)) OR
 					(reg_q1685 AND symb_decoder(16#de#)) OR
 					(reg_q1685 AND symb_decoder(16#8e#)) OR
 					(reg_q1685 AND symb_decoder(16#54#)) OR
 					(reg_q1685 AND symb_decoder(16#06#)) OR
 					(reg_q1685 AND symb_decoder(16#50#)) OR
 					(reg_q1685 AND symb_decoder(16#90#)) OR
 					(reg_q1685 AND symb_decoder(16#ac#)) OR
 					(reg_q1685 AND symb_decoder(16#a3#)) OR
 					(reg_q1685 AND symb_decoder(16#5c#)) OR
 					(reg_q1685 AND symb_decoder(16#f0#)) OR
 					(reg_q1685 AND symb_decoder(16#2a#)) OR
 					(reg_q1685 AND symb_decoder(16#ce#)) OR
 					(reg_q1685 AND symb_decoder(16#5d#)) OR
 					(reg_q1685 AND symb_decoder(16#f9#)) OR
 					(reg_q1685 AND symb_decoder(16#f4#)) OR
 					(reg_q1685 AND symb_decoder(16#9e#)) OR
 					(reg_q1685 AND symb_decoder(16#3c#)) OR
 					(reg_q1685 AND symb_decoder(16#2c#)) OR
 					(reg_q1685 AND symb_decoder(16#f2#)) OR
 					(reg_q1685 AND symb_decoder(16#71#)) OR
 					(reg_q1685 AND symb_decoder(16#27#)) OR
 					(reg_q1685 AND symb_decoder(16#0e#)) OR
 					(reg_q1685 AND symb_decoder(16#73#)) OR
 					(reg_q1685 AND symb_decoder(16#36#)) OR
 					(reg_q1685 AND symb_decoder(16#5a#)) OR
 					(reg_q1685 AND symb_decoder(16#43#)) OR
 					(reg_q1685 AND symb_decoder(16#6c#)) OR
 					(reg_q1685 AND symb_decoder(16#1a#)) OR
 					(reg_q1685 AND symb_decoder(16#2b#)) OR
 					(reg_q1685 AND symb_decoder(16#59#)) OR
 					(reg_q1685 AND symb_decoder(16#93#)) OR
 					(reg_q1685 AND symb_decoder(16#d2#)) OR
 					(reg_q1685 AND symb_decoder(16#40#)) OR
 					(reg_q1685 AND symb_decoder(16#4a#)) OR
 					(reg_q1685 AND symb_decoder(16#86#)) OR
 					(reg_q1685 AND symb_decoder(16#25#)) OR
 					(reg_q1685 AND symb_decoder(16#ef#)) OR
 					(reg_q1685 AND symb_decoder(16#c2#)) OR
 					(reg_q1685 AND symb_decoder(16#b9#)) OR
 					(reg_q1685 AND symb_decoder(16#ea#)) OR
 					(reg_q1685 AND symb_decoder(16#e0#)) OR
 					(reg_q1685 AND symb_decoder(16#81#)) OR
 					(reg_q1685 AND symb_decoder(16#61#)) OR
 					(reg_q1685 AND symb_decoder(16#1c#)) OR
 					(reg_q1685 AND symb_decoder(16#19#)) OR
 					(reg_q1685 AND symb_decoder(16#e2#)) OR
 					(reg_q1685 AND symb_decoder(16#87#)) OR
 					(reg_q1685 AND symb_decoder(16#d8#)) OR
 					(reg_q1685 AND symb_decoder(16#8d#)) OR
 					(reg_q1685 AND symb_decoder(16#e6#)) OR
 					(reg_q1685 AND symb_decoder(16#6b#)) OR
 					(reg_q1685 AND symb_decoder(16#21#)) OR
 					(reg_q1685 AND symb_decoder(16#fd#)) OR
 					(reg_q1685 AND symb_decoder(16#ae#)) OR
 					(reg_q1685 AND symb_decoder(16#6e#)) OR
 					(reg_q1685 AND symb_decoder(16#12#)) OR
 					(reg_q1685 AND symb_decoder(16#f7#)) OR
 					(reg_q1685 AND symb_decoder(16#99#)) OR
 					(reg_q1685 AND symb_decoder(16#3b#)) OR
 					(reg_q1685 AND symb_decoder(16#94#)) OR
 					(reg_q1685 AND symb_decoder(16#7a#)) OR
 					(reg_q1685 AND symb_decoder(16#41#)) OR
 					(reg_q1685 AND symb_decoder(16#e9#)) OR
 					(reg_q1685 AND symb_decoder(16#1b#)) OR
 					(reg_q1685 AND symb_decoder(16#4e#)) OR
 					(reg_q1685 AND symb_decoder(16#6f#)) OR
 					(reg_q1685 AND symb_decoder(16#ab#)) OR
 					(reg_q1685 AND symb_decoder(16#e3#)) OR
 					(reg_q1685 AND symb_decoder(16#b8#)) OR
 					(reg_q1685 AND symb_decoder(16#c6#)) OR
 					(reg_q1685 AND symb_decoder(16#52#)) OR
 					(reg_q1685 AND symb_decoder(16#5b#)) OR
 					(reg_q1685 AND symb_decoder(16#01#)) OR
 					(reg_q1685 AND symb_decoder(16#35#)) OR
 					(reg_q1685 AND symb_decoder(16#60#)) OR
 					(reg_q1685 AND symb_decoder(16#b6#)) OR
 					(reg_q1685 AND symb_decoder(16#ff#)) OR
 					(reg_q1685 AND symb_decoder(16#18#)) OR
 					(reg_q1685 AND symb_decoder(16#a8#)) OR
 					(reg_q1685 AND symb_decoder(16#62#)) OR
 					(reg_q1685 AND symb_decoder(16#dd#)) OR
 					(reg_q1685 AND symb_decoder(16#32#)) OR
 					(reg_q1685 AND symb_decoder(16#04#)) OR
 					(reg_q1685 AND symb_decoder(16#3d#)) OR
 					(reg_q1685 AND symb_decoder(16#1e#)) OR
 					(reg_q1685 AND symb_decoder(16#58#)) OR
 					(reg_q1685 AND symb_decoder(16#49#)) OR
 					(reg_q1685 AND symb_decoder(16#ec#)) OR
 					(reg_q1685 AND symb_decoder(16#5e#)) OR
 					(reg_q1685 AND symb_decoder(16#cf#)) OR
 					(reg_q1685 AND symb_decoder(16#66#)) OR
 					(reg_q1685 AND symb_decoder(16#ee#)) OR
 					(reg_q1685 AND symb_decoder(16#77#)) OR
 					(reg_q1685 AND symb_decoder(16#7d#)) OR
 					(reg_q1685 AND symb_decoder(16#64#)) OR
 					(reg_q1685 AND symb_decoder(16#13#)) OR
 					(reg_q1685 AND symb_decoder(16#29#)) OR
 					(reg_q1685 AND symb_decoder(16#37#)) OR
 					(reg_q1685 AND symb_decoder(16#57#)) OR
 					(reg_q1685 AND symb_decoder(16#70#)) OR
 					(reg_q1685 AND symb_decoder(16#92#)) OR
 					(reg_q1685 AND symb_decoder(16#af#)) OR
 					(reg_q1685 AND symb_decoder(16#bd#)) OR
 					(reg_q1685 AND symb_decoder(16#4c#)) OR
 					(reg_q1685 AND symb_decoder(16#14#)) OR
 					(reg_q1685 AND symb_decoder(16#a9#)) OR
 					(reg_q1685 AND symb_decoder(16#db#)) OR
 					(reg_q1685 AND symb_decoder(16#79#)) OR
 					(reg_q1685 AND symb_decoder(16#82#)) OR
 					(reg_q1685 AND symb_decoder(16#d9#)) OR
 					(reg_q1685 AND symb_decoder(16#4d#)) OR
 					(reg_q1685 AND symb_decoder(16#bb#)) OR
 					(reg_q1685 AND symb_decoder(16#63#)) OR
 					(reg_q1685 AND symb_decoder(16#dc#)) OR
 					(reg_q1685 AND symb_decoder(16#fb#)) OR
 					(reg_q1685 AND symb_decoder(16#97#)) OR
 					(reg_q1685 AND symb_decoder(16#47#)) OR
 					(reg_q1685 AND symb_decoder(16#d6#)) OR
 					(reg_q1685 AND symb_decoder(16#3f#)) OR
 					(reg_q1685 AND symb_decoder(16#48#)) OR
 					(reg_q1685 AND symb_decoder(16#69#)) OR
 					(reg_q1685 AND symb_decoder(16#89#)) OR
 					(reg_q1685 AND symb_decoder(16#55#)) OR
 					(reg_q1685 AND symb_decoder(16#56#)) OR
 					(reg_q1685 AND symb_decoder(16#15#)) OR
 					(reg_q1685 AND symb_decoder(16#05#)) OR
 					(reg_q1685 AND symb_decoder(16#98#)) OR
 					(reg_q1685 AND symb_decoder(16#c5#)) OR
 					(reg_q1685 AND symb_decoder(16#b0#)) OR
 					(reg_q1685 AND symb_decoder(16#95#)) OR
 					(reg_q1685 AND symb_decoder(16#f3#)) OR
 					(reg_q1685 AND symb_decoder(16#b5#)) OR
 					(reg_q1685 AND symb_decoder(16#24#)) OR
 					(reg_q1685 AND symb_decoder(16#72#)) OR
 					(reg_q1685 AND symb_decoder(16#bc#)) OR
 					(reg_q1685 AND symb_decoder(16#0c#)) OR
 					(reg_q1685 AND symb_decoder(16#33#)) OR
 					(reg_q1685 AND symb_decoder(16#c0#)) OR
 					(reg_q1685 AND symb_decoder(16#07#)) OR
 					(reg_q1685 AND symb_decoder(16#0b#)) OR
 					(reg_q1685 AND symb_decoder(16#e8#)) OR
 					(reg_q1685 AND symb_decoder(16#26#)) OR
 					(reg_q1685 AND symb_decoder(16#fa#)) OR
 					(reg_q1685 AND symb_decoder(16#67#)) OR
 					(reg_q1685 AND symb_decoder(16#ba#)) OR
 					(reg_q1685 AND symb_decoder(16#b7#)) OR
 					(reg_q1685 AND symb_decoder(16#b1#)) OR
 					(reg_q1685 AND symb_decoder(16#3e#)) OR
 					(reg_q1685 AND symb_decoder(16#8b#)) OR
 					(reg_q1685 AND symb_decoder(16#e5#)) OR
 					(reg_q1685 AND symb_decoder(16#f5#)) OR
 					(reg_q1685 AND symb_decoder(16#9a#)) OR
 					(reg_q1685 AND symb_decoder(16#11#)) OR
 					(reg_q1685 AND symb_decoder(16#e4#)) OR
 					(reg_q1685 AND symb_decoder(16#aa#)) OR
 					(reg_q1685 AND symb_decoder(16#96#)) OR
 					(reg_q1685 AND symb_decoder(16#ca#)) OR
 					(reg_q1685 AND symb_decoder(16#b4#)) OR
 					(reg_q1685 AND symb_decoder(16#91#)) OR
 					(reg_q1685 AND symb_decoder(16#2e#)) OR
 					(reg_q1685 AND symb_decoder(16#a6#)) OR
 					(reg_q1685 AND symb_decoder(16#53#)) OR
 					(reg_q1685 AND symb_decoder(16#08#)) OR
 					(reg_q1685 AND symb_decoder(16#d4#)) OR
 					(reg_q1685 AND symb_decoder(16#0a#)) OR
 					(reg_q1685 AND symb_decoder(16#f6#)) OR
 					(reg_q1685 AND symb_decoder(16#39#)) OR
 					(reg_q1685 AND symb_decoder(16#38#)) OR
 					(reg_q1685 AND symb_decoder(16#c3#)) OR
 					(reg_q1685 AND symb_decoder(16#1f#)) OR
 					(reg_q1685 AND symb_decoder(16#78#)) OR
 					(reg_q1685 AND symb_decoder(16#45#)) OR
 					(reg_q1685 AND symb_decoder(16#02#)) OR
 					(reg_q1685 AND symb_decoder(16#c8#)) OR
 					(reg_q1685 AND symb_decoder(16#c1#)) OR
 					(reg_q1685 AND symb_decoder(16#e1#)) OR
 					(reg_q1685 AND symb_decoder(16#31#)) OR
 					(reg_q1685 AND symb_decoder(16#9f#)) OR
 					(reg_q1685 AND symb_decoder(16#17#)) OR
 					(reg_q1685 AND symb_decoder(16#f8#)) OR
 					(reg_q1685 AND symb_decoder(16#b2#)) OR
 					(reg_q1685 AND symb_decoder(16#2d#)) OR
 					(reg_q1685 AND symb_decoder(16#2f#)) OR
 					(reg_q1685 AND symb_decoder(16#cd#)) OR
 					(reg_q1685 AND symb_decoder(16#65#)) OR
 					(reg_q1685 AND symb_decoder(16#51#)) OR
 					(reg_q1685 AND symb_decoder(16#c4#)) OR
 					(reg_q1685 AND symb_decoder(16#ad#)) OR
 					(reg_q1685 AND symb_decoder(16#f1#)) OR
 					(reg_q1685 AND symb_decoder(16#9c#)) OR
 					(reg_q1685 AND symb_decoder(16#d7#)) OR
 					(reg_q1685 AND symb_decoder(16#c7#)) OR
 					(reg_q1685 AND symb_decoder(16#8c#)) OR
 					(reg_q1685 AND symb_decoder(16#fe#)) OR
 					(reg_q1685 AND symb_decoder(16#85#)) OR
 					(reg_q1685 AND symb_decoder(16#23#)) OR
 					(reg_q1685 AND symb_decoder(16#4b#)) OR
 					(reg_q1685 AND symb_decoder(16#80#)) OR
 					(reg_q1685 AND symb_decoder(16#d0#)) OR
 					(reg_q1685 AND symb_decoder(16#75#)) OR
 					(reg_q1685 AND symb_decoder(16#10#)) OR
 					(reg_q1685 AND symb_decoder(16#d1#)) OR
 					(reg_q1685 AND symb_decoder(16#84#)) OR
 					(reg_q1685 AND symb_decoder(16#68#)) OR
 					(reg_q1685 AND symb_decoder(16#3a#)) OR
 					(reg_q1685 AND symb_decoder(16#8f#)) OR
 					(reg_q1685 AND symb_decoder(16#88#)) OR
 					(reg_q1685 AND symb_decoder(16#7e#)) OR
 					(reg_q1685 AND symb_decoder(16#09#)) OR
 					(reg_q1685 AND symb_decoder(16#74#)) OR
 					(reg_q1685 AND symb_decoder(16#b3#)) OR
 					(reg_q1685 AND symb_decoder(16#42#)) OR
 					(reg_q1685 AND symb_decoder(16#c9#)) OR
 					(reg_q1685 AND symb_decoder(16#7b#)) OR
 					(reg_q1685 AND symb_decoder(16#28#)) OR
 					(reg_q1685 AND symb_decoder(16#5f#)) OR
 					(reg_q1685 AND symb_decoder(16#30#)) OR
 					(reg_q1685 AND symb_decoder(16#16#)) OR
 					(reg_q1685 AND symb_decoder(16#44#)) OR
 					(reg_q1685 AND symb_decoder(16#0f#)) OR
 					(reg_q1685 AND symb_decoder(16#20#)) OR
 					(reg_q1685 AND symb_decoder(16#6a#)) OR
 					(reg_q1685 AND symb_decoder(16#34#)) OR
 					(reg_q1685 AND symb_decoder(16#a4#)) OR
 					(reg_q1685 AND symb_decoder(16#a0#)) OR
 					(reg_q1685 AND symb_decoder(16#fc#)) OR
 					(reg_q1685 AND symb_decoder(16#e7#)) OR
 					(reg_q1685 AND symb_decoder(16#d3#)) OR
 					(reg_q1685 AND symb_decoder(16#bf#)) OR
 					(reg_q1685 AND symb_decoder(16#a1#)) OR
 					(reg_q1685 AND symb_decoder(16#ed#)) OR
 					(reg_q1685 AND symb_decoder(16#a2#)) OR
 					(reg_q1685 AND symb_decoder(16#9d#)) OR
 					(reg_q1685 AND symb_decoder(16#7f#)) OR
 					(reg_q1685 AND symb_decoder(16#46#)) OR
 					(reg_q1685 AND symb_decoder(16#1d#));
reg_q1685_init <= '0' ;
	p_reg_q1685: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1685 <= reg_q1685_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1685 <= reg_q1685_init;
        else
          reg_q1685 <= reg_q1685_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2633_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q2633 AND symb_decoder(16#3c#)) OR
 					(reg_q2633 AND symb_decoder(16#16#)) OR
 					(reg_q2633 AND symb_decoder(16#be#)) OR
 					(reg_q2633 AND symb_decoder(16#13#)) OR
 					(reg_q2633 AND symb_decoder(16#20#)) OR
 					(reg_q2633 AND symb_decoder(16#e6#)) OR
 					(reg_q2633 AND symb_decoder(16#a1#)) OR
 					(reg_q2633 AND symb_decoder(16#9d#)) OR
 					(reg_q2633 AND symb_decoder(16#f6#)) OR
 					(reg_q2633 AND symb_decoder(16#0a#)) OR
 					(reg_q2633 AND symb_decoder(16#c5#)) OR
 					(reg_q2633 AND symb_decoder(16#11#)) OR
 					(reg_q2633 AND symb_decoder(16#4f#)) OR
 					(reg_q2633 AND symb_decoder(16#61#)) OR
 					(reg_q2633 AND symb_decoder(16#50#)) OR
 					(reg_q2633 AND symb_decoder(16#33#)) OR
 					(reg_q2633 AND symb_decoder(16#b5#)) OR
 					(reg_q2633 AND symb_decoder(16#91#)) OR
 					(reg_q2633 AND symb_decoder(16#a2#)) OR
 					(reg_q2633 AND symb_decoder(16#66#)) OR
 					(reg_q2633 AND symb_decoder(16#72#)) OR
 					(reg_q2633 AND symb_decoder(16#53#)) OR
 					(reg_q2633 AND symb_decoder(16#1c#)) OR
 					(reg_q2633 AND symb_decoder(16#03#)) OR
 					(reg_q2633 AND symb_decoder(16#c4#)) OR
 					(reg_q2633 AND symb_decoder(16#34#)) OR
 					(reg_q2633 AND symb_decoder(16#48#)) OR
 					(reg_q2633 AND symb_decoder(16#f2#)) OR
 					(reg_q2633 AND symb_decoder(16#9a#)) OR
 					(reg_q2633 AND symb_decoder(16#98#)) OR
 					(reg_q2633 AND symb_decoder(16#01#)) OR
 					(reg_q2633 AND symb_decoder(16#c1#)) OR
 					(reg_q2633 AND symb_decoder(16#8a#)) OR
 					(reg_q2633 AND symb_decoder(16#ed#)) OR
 					(reg_q2633 AND symb_decoder(16#55#)) OR
 					(reg_q2633 AND symb_decoder(16#09#)) OR
 					(reg_q2633 AND symb_decoder(16#7c#)) OR
 					(reg_q2633 AND symb_decoder(16#c8#)) OR
 					(reg_q2633 AND symb_decoder(16#2c#)) OR
 					(reg_q2633 AND symb_decoder(16#7e#)) OR
 					(reg_q2633 AND symb_decoder(16#d0#)) OR
 					(reg_q2633 AND symb_decoder(16#e4#)) OR
 					(reg_q2633 AND symb_decoder(16#64#)) OR
 					(reg_q2633 AND symb_decoder(16#04#)) OR
 					(reg_q2633 AND symb_decoder(16#ab#)) OR
 					(reg_q2633 AND symb_decoder(16#a6#)) OR
 					(reg_q2633 AND symb_decoder(16#22#)) OR
 					(reg_q2633 AND symb_decoder(16#39#)) OR
 					(reg_q2633 AND symb_decoder(16#63#)) OR
 					(reg_q2633 AND symb_decoder(16#82#)) OR
 					(reg_q2633 AND symb_decoder(16#1e#)) OR
 					(reg_q2633 AND symb_decoder(16#ff#)) OR
 					(reg_q2633 AND symb_decoder(16#17#)) OR
 					(reg_q2633 AND symb_decoder(16#41#)) OR
 					(reg_q2633 AND symb_decoder(16#a4#)) OR
 					(reg_q2633 AND symb_decoder(16#cb#)) OR
 					(reg_q2633 AND symb_decoder(16#5d#)) OR
 					(reg_q2633 AND symb_decoder(16#fd#)) OR
 					(reg_q2633 AND symb_decoder(16#54#)) OR
 					(reg_q2633 AND symb_decoder(16#30#)) OR
 					(reg_q2633 AND symb_decoder(16#2d#)) OR
 					(reg_q2633 AND symb_decoder(16#d3#)) OR
 					(reg_q2633 AND symb_decoder(16#9c#)) OR
 					(reg_q2633 AND symb_decoder(16#86#)) OR
 					(reg_q2633 AND symb_decoder(16#e7#)) OR
 					(reg_q2633 AND symb_decoder(16#fe#)) OR
 					(reg_q2633 AND symb_decoder(16#7f#)) OR
 					(reg_q2633 AND symb_decoder(16#8b#)) OR
 					(reg_q2633 AND symb_decoder(16#dd#)) OR
 					(reg_q2633 AND symb_decoder(16#3a#)) OR
 					(reg_q2633 AND symb_decoder(16#b3#)) OR
 					(reg_q2633 AND symb_decoder(16#71#)) OR
 					(reg_q2633 AND symb_decoder(16#4d#)) OR
 					(reg_q2633 AND symb_decoder(16#a9#)) OR
 					(reg_q2633 AND symb_decoder(16#70#)) OR
 					(reg_q2633 AND symb_decoder(16#aa#)) OR
 					(reg_q2633 AND symb_decoder(16#ee#)) OR
 					(reg_q2633 AND symb_decoder(16#2e#)) OR
 					(reg_q2633 AND symb_decoder(16#bb#)) OR
 					(reg_q2633 AND symb_decoder(16#c2#)) OR
 					(reg_q2633 AND symb_decoder(16#3e#)) OR
 					(reg_q2633 AND symb_decoder(16#6d#)) OR
 					(reg_q2633 AND symb_decoder(16#6b#)) OR
 					(reg_q2633 AND symb_decoder(16#83#)) OR
 					(reg_q2633 AND symb_decoder(16#4b#)) OR
 					(reg_q2633 AND symb_decoder(16#1a#)) OR
 					(reg_q2633 AND symb_decoder(16#87#)) OR
 					(reg_q2633 AND symb_decoder(16#b7#)) OR
 					(reg_q2633 AND symb_decoder(16#e5#)) OR
 					(reg_q2633 AND symb_decoder(16#ad#)) OR
 					(reg_q2633 AND symb_decoder(16#5a#)) OR
 					(reg_q2633 AND symb_decoder(16#c7#)) OR
 					(reg_q2633 AND symb_decoder(16#24#)) OR
 					(reg_q2633 AND symb_decoder(16#57#)) OR
 					(reg_q2633 AND symb_decoder(16#b9#)) OR
 					(reg_q2633 AND symb_decoder(16#d9#)) OR
 					(reg_q2633 AND symb_decoder(16#0e#)) OR
 					(reg_q2633 AND symb_decoder(16#3d#)) OR
 					(reg_q2633 AND symb_decoder(16#a8#)) OR
 					(reg_q2633 AND symb_decoder(16#b8#)) OR
 					(reg_q2633 AND symb_decoder(16#05#)) OR
 					(reg_q2633 AND symb_decoder(16#e1#)) OR
 					(reg_q2633 AND symb_decoder(16#37#)) OR
 					(reg_q2633 AND symb_decoder(16#1b#)) OR
 					(reg_q2633 AND symb_decoder(16#db#)) OR
 					(reg_q2633 AND symb_decoder(16#f1#)) OR
 					(reg_q2633 AND symb_decoder(16#d8#)) OR
 					(reg_q2633 AND symb_decoder(16#d6#)) OR
 					(reg_q2633 AND symb_decoder(16#47#)) OR
 					(reg_q2633 AND symb_decoder(16#81#)) OR
 					(reg_q2633 AND symb_decoder(16#b0#)) OR
 					(reg_q2633 AND symb_decoder(16#a5#)) OR
 					(reg_q2633 AND symb_decoder(16#d5#)) OR
 					(reg_q2633 AND symb_decoder(16#15#)) OR
 					(reg_q2633 AND symb_decoder(16#31#)) OR
 					(reg_q2633 AND symb_decoder(16#e9#)) OR
 					(reg_q2633 AND symb_decoder(16#52#)) OR
 					(reg_q2633 AND symb_decoder(16#d1#)) OR
 					(reg_q2633 AND symb_decoder(16#9e#)) OR
 					(reg_q2633 AND symb_decoder(16#0c#)) OR
 					(reg_q2633 AND symb_decoder(16#6a#)) OR
 					(reg_q2633 AND symb_decoder(16#ec#)) OR
 					(reg_q2633 AND symb_decoder(16#40#)) OR
 					(reg_q2633 AND symb_decoder(16#56#)) OR
 					(reg_q2633 AND symb_decoder(16#a7#)) OR
 					(reg_q2633 AND symb_decoder(16#1f#)) OR
 					(reg_q2633 AND symb_decoder(16#2b#)) OR
 					(reg_q2633 AND symb_decoder(16#74#)) OR
 					(reg_q2633 AND symb_decoder(16#28#)) OR
 					(reg_q2633 AND symb_decoder(16#79#)) OR
 					(reg_q2633 AND symb_decoder(16#df#)) OR
 					(reg_q2633 AND symb_decoder(16#d7#)) OR
 					(reg_q2633 AND symb_decoder(16#80#)) OR
 					(reg_q2633 AND symb_decoder(16#3b#)) OR
 					(reg_q2633 AND symb_decoder(16#f7#)) OR
 					(reg_q2633 AND symb_decoder(16#2f#)) OR
 					(reg_q2633 AND symb_decoder(16#95#)) OR
 					(reg_q2633 AND symb_decoder(16#49#)) OR
 					(reg_q2633 AND symb_decoder(16#4a#)) OR
 					(reg_q2633 AND symb_decoder(16#ea#)) OR
 					(reg_q2633 AND symb_decoder(16#60#)) OR
 					(reg_q2633 AND symb_decoder(16#ac#)) OR
 					(reg_q2633 AND symb_decoder(16#8e#)) OR
 					(reg_q2633 AND symb_decoder(16#3f#)) OR
 					(reg_q2633 AND symb_decoder(16#0b#)) OR
 					(reg_q2633 AND symb_decoder(16#8d#)) OR
 					(reg_q2633 AND symb_decoder(16#21#)) OR
 					(reg_q2633 AND symb_decoder(16#32#)) OR
 					(reg_q2633 AND symb_decoder(16#94#)) OR
 					(reg_q2633 AND symb_decoder(16#bf#)) OR
 					(reg_q2633 AND symb_decoder(16#fc#)) OR
 					(reg_q2633 AND symb_decoder(16#84#)) OR
 					(reg_q2633 AND symb_decoder(16#77#)) OR
 					(reg_q2633 AND symb_decoder(16#14#)) OR
 					(reg_q2633 AND symb_decoder(16#23#)) OR
 					(reg_q2633 AND symb_decoder(16#69#)) OR
 					(reg_q2633 AND symb_decoder(16#f4#)) OR
 					(reg_q2633 AND symb_decoder(16#a3#)) OR
 					(reg_q2633 AND symb_decoder(16#2a#)) OR
 					(reg_q2633 AND symb_decoder(16#38#)) OR
 					(reg_q2633 AND symb_decoder(16#89#)) OR
 					(reg_q2633 AND symb_decoder(16#c0#)) OR
 					(reg_q2633 AND symb_decoder(16#78#)) OR
 					(reg_q2633 AND symb_decoder(16#76#)) OR
 					(reg_q2633 AND symb_decoder(16#7a#)) OR
 					(reg_q2633 AND symb_decoder(16#b4#)) OR
 					(reg_q2633 AND symb_decoder(16#36#)) OR
 					(reg_q2633 AND symb_decoder(16#07#)) OR
 					(reg_q2633 AND symb_decoder(16#9b#)) OR
 					(reg_q2633 AND symb_decoder(16#7b#)) OR
 					(reg_q2633 AND symb_decoder(16#58#)) OR
 					(reg_q2633 AND symb_decoder(16#45#)) OR
 					(reg_q2633 AND symb_decoder(16#f8#)) OR
 					(reg_q2633 AND symb_decoder(16#8f#)) OR
 					(reg_q2633 AND symb_decoder(16#1d#)) OR
 					(reg_q2633 AND symb_decoder(16#12#)) OR
 					(reg_q2633 AND symb_decoder(16#fa#)) OR
 					(reg_q2633 AND symb_decoder(16#96#)) OR
 					(reg_q2633 AND symb_decoder(16#75#)) OR
 					(reg_q2633 AND symb_decoder(16#dc#)) OR
 					(reg_q2633 AND symb_decoder(16#e8#)) OR
 					(reg_q2633 AND symb_decoder(16#51#)) OR
 					(reg_q2633 AND symb_decoder(16#02#)) OR
 					(reg_q2633 AND symb_decoder(16#cf#)) OR
 					(reg_q2633 AND symb_decoder(16#85#)) OR
 					(reg_q2633 AND symb_decoder(16#ba#)) OR
 					(reg_q2633 AND symb_decoder(16#88#)) OR
 					(reg_q2633 AND symb_decoder(16#65#)) OR
 					(reg_q2633 AND symb_decoder(16#ef#)) OR
 					(reg_q2633 AND symb_decoder(16#cc#)) OR
 					(reg_q2633 AND symb_decoder(16#73#)) OR
 					(reg_q2633 AND symb_decoder(16#99#)) OR
 					(reg_q2633 AND symb_decoder(16#29#)) OR
 					(reg_q2633 AND symb_decoder(16#c3#)) OR
 					(reg_q2633 AND symb_decoder(16#a0#)) OR
 					(reg_q2633 AND symb_decoder(16#6c#)) OR
 					(reg_q2633 AND symb_decoder(16#6e#)) OR
 					(reg_q2633 AND symb_decoder(16#5f#)) OR
 					(reg_q2633 AND symb_decoder(16#cd#)) OR
 					(reg_q2633 AND symb_decoder(16#af#)) OR
 					(reg_q2633 AND symb_decoder(16#c6#)) OR
 					(reg_q2633 AND symb_decoder(16#c9#)) OR
 					(reg_q2633 AND symb_decoder(16#42#)) OR
 					(reg_q2633 AND symb_decoder(16#5e#)) OR
 					(reg_q2633 AND symb_decoder(16#92#)) OR
 					(reg_q2633 AND symb_decoder(16#27#)) OR
 					(reg_q2633 AND symb_decoder(16#5b#)) OR
 					(reg_q2633 AND symb_decoder(16#97#)) OR
 					(reg_q2633 AND symb_decoder(16#ce#)) OR
 					(reg_q2633 AND symb_decoder(16#0f#)) OR
 					(reg_q2633 AND symb_decoder(16#e3#)) OR
 					(reg_q2633 AND symb_decoder(16#4e#)) OR
 					(reg_q2633 AND symb_decoder(16#e0#)) OR
 					(reg_q2633 AND symb_decoder(16#35#)) OR
 					(reg_q2633 AND symb_decoder(16#26#)) OR
 					(reg_q2633 AND symb_decoder(16#f9#)) OR
 					(reg_q2633 AND symb_decoder(16#bc#)) OR
 					(reg_q2633 AND symb_decoder(16#8c#)) OR
 					(reg_q2633 AND symb_decoder(16#00#)) OR
 					(reg_q2633 AND symb_decoder(16#e2#)) OR
 					(reg_q2633 AND symb_decoder(16#f5#)) OR
 					(reg_q2633 AND symb_decoder(16#18#)) OR
 					(reg_q2633 AND symb_decoder(16#67#)) OR
 					(reg_q2633 AND symb_decoder(16#d4#)) OR
 					(reg_q2633 AND symb_decoder(16#0d#)) OR
 					(reg_q2633 AND symb_decoder(16#46#)) OR
 					(reg_q2633 AND symb_decoder(16#b6#)) OR
 					(reg_q2633 AND symb_decoder(16#93#)) OR
 					(reg_q2633 AND symb_decoder(16#9f#)) OR
 					(reg_q2633 AND symb_decoder(16#ca#)) OR
 					(reg_q2633 AND symb_decoder(16#4c#)) OR
 					(reg_q2633 AND symb_decoder(16#62#)) OR
 					(reg_q2633 AND symb_decoder(16#90#)) OR
 					(reg_q2633 AND symb_decoder(16#d2#)) OR
 					(reg_q2633 AND symb_decoder(16#6f#)) OR
 					(reg_q2633 AND symb_decoder(16#b2#)) OR
 					(reg_q2633 AND symb_decoder(16#fb#)) OR
 					(reg_q2633 AND symb_decoder(16#7d#)) OR
 					(reg_q2633 AND symb_decoder(16#ae#)) OR
 					(reg_q2633 AND symb_decoder(16#bd#)) OR
 					(reg_q2633 AND symb_decoder(16#06#)) OR
 					(reg_q2633 AND symb_decoder(16#44#)) OR
 					(reg_q2633 AND symb_decoder(16#68#)) OR
 					(reg_q2633 AND symb_decoder(16#da#)) OR
 					(reg_q2633 AND symb_decoder(16#eb#)) OR
 					(reg_q2633 AND symb_decoder(16#5c#)) OR
 					(reg_q2633 AND symb_decoder(16#59#)) OR
 					(reg_q2633 AND symb_decoder(16#08#)) OR
 					(reg_q2633 AND symb_decoder(16#10#)) OR
 					(reg_q2633 AND symb_decoder(16#b1#)) OR
 					(reg_q2633 AND symb_decoder(16#f0#)) OR
 					(reg_q2633 AND symb_decoder(16#19#)) OR
 					(reg_q2633 AND symb_decoder(16#de#)) OR
 					(reg_q2633 AND symb_decoder(16#25#)) OR
 					(reg_q2633 AND symb_decoder(16#f3#)) OR
 					(reg_q2633 AND symb_decoder(16#43#));
reg_q2633_init <= '0' ;
	p_reg_q2633: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2633 <= reg_q2633_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2633 <= reg_q2633_init;
        else
          reg_q2633 <= reg_q2633_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1395_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1395 AND symb_decoder(16#56#)) OR
 					(reg_q1395 AND symb_decoder(16#b4#)) OR
 					(reg_q1395 AND symb_decoder(16#b3#)) OR
 					(reg_q1395 AND symb_decoder(16#5b#)) OR
 					(reg_q1395 AND symb_decoder(16#35#)) OR
 					(reg_q1395 AND symb_decoder(16#93#)) OR
 					(reg_q1395 AND symb_decoder(16#19#)) OR
 					(reg_q1395 AND symb_decoder(16#ca#)) OR
 					(reg_q1395 AND symb_decoder(16#3f#)) OR
 					(reg_q1395 AND symb_decoder(16#b0#)) OR
 					(reg_q1395 AND symb_decoder(16#01#)) OR
 					(reg_q1395 AND symb_decoder(16#ac#)) OR
 					(reg_q1395 AND symb_decoder(16#ee#)) OR
 					(reg_q1395 AND symb_decoder(16#f7#)) OR
 					(reg_q1395 AND symb_decoder(16#dd#)) OR
 					(reg_q1395 AND symb_decoder(16#ae#)) OR
 					(reg_q1395 AND symb_decoder(16#8d#)) OR
 					(reg_q1395 AND symb_decoder(16#88#)) OR
 					(reg_q1395 AND symb_decoder(16#39#)) OR
 					(reg_q1395 AND symb_decoder(16#2e#)) OR
 					(reg_q1395 AND symb_decoder(16#c1#)) OR
 					(reg_q1395 AND symb_decoder(16#58#)) OR
 					(reg_q1395 AND symb_decoder(16#85#)) OR
 					(reg_q1395 AND symb_decoder(16#2a#)) OR
 					(reg_q1395 AND symb_decoder(16#32#)) OR
 					(reg_q1395 AND symb_decoder(16#d7#)) OR
 					(reg_q1395 AND symb_decoder(16#71#)) OR
 					(reg_q1395 AND symb_decoder(16#57#)) OR
 					(reg_q1395 AND symb_decoder(16#34#)) OR
 					(reg_q1395 AND symb_decoder(16#90#)) OR
 					(reg_q1395 AND symb_decoder(16#bf#)) OR
 					(reg_q1395 AND symb_decoder(16#25#)) OR
 					(reg_q1395 AND symb_decoder(16#a4#)) OR
 					(reg_q1395 AND symb_decoder(16#16#)) OR
 					(reg_q1395 AND symb_decoder(16#3b#)) OR
 					(reg_q1395 AND symb_decoder(16#50#)) OR
 					(reg_q1395 AND symb_decoder(16#fa#)) OR
 					(reg_q1395 AND symb_decoder(16#c5#)) OR
 					(reg_q1395 AND symb_decoder(16#0b#)) OR
 					(reg_q1395 AND symb_decoder(16#4e#)) OR
 					(reg_q1395 AND symb_decoder(16#08#)) OR
 					(reg_q1395 AND symb_decoder(16#74#)) OR
 					(reg_q1395 AND symb_decoder(16#31#)) OR
 					(reg_q1395 AND symb_decoder(16#67#)) OR
 					(reg_q1395 AND symb_decoder(16#f0#)) OR
 					(reg_q1395 AND symb_decoder(16#f2#)) OR
 					(reg_q1395 AND symb_decoder(16#3d#)) OR
 					(reg_q1395 AND symb_decoder(16#84#)) OR
 					(reg_q1395 AND symb_decoder(16#f1#)) OR
 					(reg_q1395 AND symb_decoder(16#86#)) OR
 					(reg_q1395 AND symb_decoder(16#79#)) OR
 					(reg_q1395 AND symb_decoder(16#1d#)) OR
 					(reg_q1395 AND symb_decoder(16#60#)) OR
 					(reg_q1395 AND symb_decoder(16#7a#)) OR
 					(reg_q1395 AND symb_decoder(16#d0#)) OR
 					(reg_q1395 AND symb_decoder(16#d4#)) OR
 					(reg_q1395 AND symb_decoder(16#ba#)) OR
 					(reg_q1395 AND symb_decoder(16#be#)) OR
 					(reg_q1395 AND symb_decoder(16#ff#)) OR
 					(reg_q1395 AND symb_decoder(16#af#)) OR
 					(reg_q1395 AND symb_decoder(16#61#)) OR
 					(reg_q1395 AND symb_decoder(16#ad#)) OR
 					(reg_q1395 AND symb_decoder(16#87#)) OR
 					(reg_q1395 AND symb_decoder(16#e4#)) OR
 					(reg_q1395 AND symb_decoder(16#06#)) OR
 					(reg_q1395 AND symb_decoder(16#3e#)) OR
 					(reg_q1395 AND symb_decoder(16#b8#)) OR
 					(reg_q1395 AND symb_decoder(16#44#)) OR
 					(reg_q1395 AND symb_decoder(16#13#)) OR
 					(reg_q1395 AND symb_decoder(16#a2#)) OR
 					(reg_q1395 AND symb_decoder(16#e6#)) OR
 					(reg_q1395 AND symb_decoder(16#d8#)) OR
 					(reg_q1395 AND symb_decoder(16#db#)) OR
 					(reg_q1395 AND symb_decoder(16#ef#)) OR
 					(reg_q1395 AND symb_decoder(16#05#)) OR
 					(reg_q1395 AND symb_decoder(16#72#)) OR
 					(reg_q1395 AND symb_decoder(16#8f#)) OR
 					(reg_q1395 AND symb_decoder(16#dc#)) OR
 					(reg_q1395 AND symb_decoder(16#e3#)) OR
 					(reg_q1395 AND symb_decoder(16#2d#)) OR
 					(reg_q1395 AND symb_decoder(16#c3#)) OR
 					(reg_q1395 AND symb_decoder(16#96#)) OR
 					(reg_q1395 AND symb_decoder(16#62#)) OR
 					(reg_q1395 AND symb_decoder(16#c4#)) OR
 					(reg_q1395 AND symb_decoder(16#e0#)) OR
 					(reg_q1395 AND symb_decoder(16#fb#)) OR
 					(reg_q1395 AND symb_decoder(16#b5#)) OR
 					(reg_q1395 AND symb_decoder(16#68#)) OR
 					(reg_q1395 AND symb_decoder(16#aa#)) OR
 					(reg_q1395 AND symb_decoder(16#fe#)) OR
 					(reg_q1395 AND symb_decoder(16#23#)) OR
 					(reg_q1395 AND symb_decoder(16#b9#)) OR
 					(reg_q1395 AND symb_decoder(16#da#)) OR
 					(reg_q1395 AND symb_decoder(16#4f#)) OR
 					(reg_q1395 AND symb_decoder(16#f8#)) OR
 					(reg_q1395 AND symb_decoder(16#e5#)) OR
 					(reg_q1395 AND symb_decoder(16#e1#)) OR
 					(reg_q1395 AND symb_decoder(16#a3#)) OR
 					(reg_q1395 AND symb_decoder(16#c9#)) OR
 					(reg_q1395 AND symb_decoder(16#8e#)) OR
 					(reg_q1395 AND symb_decoder(16#65#)) OR
 					(reg_q1395 AND symb_decoder(16#99#)) OR
 					(reg_q1395 AND symb_decoder(16#20#)) OR
 					(reg_q1395 AND symb_decoder(16#5e#)) OR
 					(reg_q1395 AND symb_decoder(16#36#)) OR
 					(reg_q1395 AND symb_decoder(16#75#)) OR
 					(reg_q1395 AND symb_decoder(16#a1#)) OR
 					(reg_q1395 AND symb_decoder(16#46#)) OR
 					(reg_q1395 AND symb_decoder(16#7f#)) OR
 					(reg_q1395 AND symb_decoder(16#6f#)) OR
 					(reg_q1395 AND symb_decoder(16#00#)) OR
 					(reg_q1395 AND symb_decoder(16#e9#)) OR
 					(reg_q1395 AND symb_decoder(16#c0#)) OR
 					(reg_q1395 AND symb_decoder(16#cc#)) OR
 					(reg_q1395 AND symb_decoder(16#5a#)) OR
 					(reg_q1395 AND symb_decoder(16#47#)) OR
 					(reg_q1395 AND symb_decoder(16#98#)) OR
 					(reg_q1395 AND symb_decoder(16#df#)) OR
 					(reg_q1395 AND symb_decoder(16#78#)) OR
 					(reg_q1395 AND symb_decoder(16#10#)) OR
 					(reg_q1395 AND symb_decoder(16#17#)) OR
 					(reg_q1395 AND symb_decoder(16#30#)) OR
 					(reg_q1395 AND symb_decoder(16#6b#)) OR
 					(reg_q1395 AND symb_decoder(16#3a#)) OR
 					(reg_q1395 AND symb_decoder(16#bc#)) OR
 					(reg_q1395 AND symb_decoder(16#43#)) OR
 					(reg_q1395 AND symb_decoder(16#1c#)) OR
 					(reg_q1395 AND symb_decoder(16#63#)) OR
 					(reg_q1395 AND symb_decoder(16#a8#)) OR
 					(reg_q1395 AND symb_decoder(16#73#)) OR
 					(reg_q1395 AND symb_decoder(16#66#)) OR
 					(reg_q1395 AND symb_decoder(16#d3#)) OR
 					(reg_q1395 AND symb_decoder(16#ed#)) OR
 					(reg_q1395 AND symb_decoder(16#02#)) OR
 					(reg_q1395 AND symb_decoder(16#d9#)) OR
 					(reg_q1395 AND symb_decoder(16#bb#)) OR
 					(reg_q1395 AND symb_decoder(16#5f#)) OR
 					(reg_q1395 AND symb_decoder(16#49#)) OR
 					(reg_q1395 AND symb_decoder(16#1b#)) OR
 					(reg_q1395 AND symb_decoder(16#29#)) OR
 					(reg_q1395 AND symb_decoder(16#ab#)) OR
 					(reg_q1395 AND symb_decoder(16#8b#)) OR
 					(reg_q1395 AND symb_decoder(16#9b#)) OR
 					(reg_q1395 AND symb_decoder(16#c6#)) OR
 					(reg_q1395 AND symb_decoder(16#7c#)) OR
 					(reg_q1395 AND symb_decoder(16#c2#)) OR
 					(reg_q1395 AND symb_decoder(16#cb#)) OR
 					(reg_q1395 AND symb_decoder(16#91#)) OR
 					(reg_q1395 AND symb_decoder(16#77#)) OR
 					(reg_q1395 AND symb_decoder(16#a7#)) OR
 					(reg_q1395 AND symb_decoder(16#c8#)) OR
 					(reg_q1395 AND symb_decoder(16#45#)) OR
 					(reg_q1395 AND symb_decoder(16#0c#)) OR
 					(reg_q1395 AND symb_decoder(16#24#)) OR
 					(reg_q1395 AND symb_decoder(16#54#)) OR
 					(reg_q1395 AND symb_decoder(16#33#)) OR
 					(reg_q1395 AND symb_decoder(16#cf#)) OR
 					(reg_q1395 AND symb_decoder(16#7d#)) OR
 					(reg_q1395 AND symb_decoder(16#d2#)) OR
 					(reg_q1395 AND symb_decoder(16#15#)) OR
 					(reg_q1395 AND symb_decoder(16#4d#)) OR
 					(reg_q1395 AND symb_decoder(16#09#)) OR
 					(reg_q1395 AND symb_decoder(16#38#)) OR
 					(reg_q1395 AND symb_decoder(16#bd#)) OR
 					(reg_q1395 AND symb_decoder(16#d1#)) OR
 					(reg_q1395 AND symb_decoder(16#9c#)) OR
 					(reg_q1395 AND symb_decoder(16#04#)) OR
 					(reg_q1395 AND symb_decoder(16#80#)) OR
 					(reg_q1395 AND symb_decoder(16#9d#)) OR
 					(reg_q1395 AND symb_decoder(16#2f#)) OR
 					(reg_q1395 AND symb_decoder(16#ce#)) OR
 					(reg_q1395 AND symb_decoder(16#6e#)) OR
 					(reg_q1395 AND symb_decoder(16#fd#)) OR
 					(reg_q1395 AND symb_decoder(16#e2#)) OR
 					(reg_q1395 AND symb_decoder(16#e7#)) OR
 					(reg_q1395 AND symb_decoder(16#81#)) OR
 					(reg_q1395 AND symb_decoder(16#ec#)) OR
 					(reg_q1395 AND symb_decoder(16#6d#)) OR
 					(reg_q1395 AND symb_decoder(16#03#)) OR
 					(reg_q1395 AND symb_decoder(16#26#)) OR
 					(reg_q1395 AND symb_decoder(16#0f#)) OR
 					(reg_q1395 AND symb_decoder(16#b1#)) OR
 					(reg_q1395 AND symb_decoder(16#2c#)) OR
 					(reg_q1395 AND symb_decoder(16#6a#)) OR
 					(reg_q1395 AND symb_decoder(16#14#)) OR
 					(reg_q1395 AND symb_decoder(16#f6#)) OR
 					(reg_q1395 AND symb_decoder(16#95#)) OR
 					(reg_q1395 AND symb_decoder(16#22#)) OR
 					(reg_q1395 AND symb_decoder(16#cd#)) OR
 					(reg_q1395 AND symb_decoder(16#a6#)) OR
 					(reg_q1395 AND symb_decoder(16#7b#)) OR
 					(reg_q1395 AND symb_decoder(16#ea#)) OR
 					(reg_q1395 AND symb_decoder(16#42#)) OR
 					(reg_q1395 AND symb_decoder(16#f9#)) OR
 					(reg_q1395 AND symb_decoder(16#11#)) OR
 					(reg_q1395 AND symb_decoder(16#b7#)) OR
 					(reg_q1395 AND symb_decoder(16#8c#)) OR
 					(reg_q1395 AND symb_decoder(16#9f#)) OR
 					(reg_q1395 AND symb_decoder(16#51#)) OR
 					(reg_q1395 AND symb_decoder(16#f4#)) OR
 					(reg_q1395 AND symb_decoder(16#fc#)) OR
 					(reg_q1395 AND symb_decoder(16#b6#)) OR
 					(reg_q1395 AND symb_decoder(16#d6#)) OR
 					(reg_q1395 AND symb_decoder(16#de#)) OR
 					(reg_q1395 AND symb_decoder(16#8a#)) OR
 					(reg_q1395 AND symb_decoder(16#a0#)) OR
 					(reg_q1395 AND symb_decoder(16#4a#)) OR
 					(reg_q1395 AND symb_decoder(16#64#)) OR
 					(reg_q1395 AND symb_decoder(16#27#)) OR
 					(reg_q1395 AND symb_decoder(16#5d#)) OR
 					(reg_q1395 AND symb_decoder(16#7e#)) OR
 					(reg_q1395 AND symb_decoder(16#1e#)) OR
 					(reg_q1395 AND symb_decoder(16#1f#)) OR
 					(reg_q1395 AND symb_decoder(16#f5#)) OR
 					(reg_q1395 AND symb_decoder(16#83#)) OR
 					(reg_q1395 AND symb_decoder(16#d5#)) OR
 					(reg_q1395 AND symb_decoder(16#4b#)) OR
 					(reg_q1395 AND symb_decoder(16#12#)) OR
 					(reg_q1395 AND symb_decoder(16#4c#)) OR
 					(reg_q1395 AND symb_decoder(16#1a#)) OR
 					(reg_q1395 AND symb_decoder(16#f3#)) OR
 					(reg_q1395 AND symb_decoder(16#70#)) OR
 					(reg_q1395 AND symb_decoder(16#97#)) OR
 					(reg_q1395 AND symb_decoder(16#2b#)) OR
 					(reg_q1395 AND symb_decoder(16#40#)) OR
 					(reg_q1395 AND symb_decoder(16#9e#)) OR
 					(reg_q1395 AND symb_decoder(16#52#)) OR
 					(reg_q1395 AND symb_decoder(16#53#)) OR
 					(reg_q1395 AND symb_decoder(16#5c#)) OR
 					(reg_q1395 AND symb_decoder(16#3c#)) OR
 					(reg_q1395 AND symb_decoder(16#89#)) OR
 					(reg_q1395 AND symb_decoder(16#6c#)) OR
 					(reg_q1395 AND symb_decoder(16#37#)) OR
 					(reg_q1395 AND symb_decoder(16#c7#)) OR
 					(reg_q1395 AND symb_decoder(16#18#)) OR
 					(reg_q1395 AND symb_decoder(16#e8#)) OR
 					(reg_q1395 AND symb_decoder(16#0d#)) OR
 					(reg_q1395 AND symb_decoder(16#94#)) OR
 					(reg_q1395 AND symb_decoder(16#0a#)) OR
 					(reg_q1395 AND symb_decoder(16#07#)) OR
 					(reg_q1395 AND symb_decoder(16#eb#)) OR
 					(reg_q1395 AND symb_decoder(16#69#)) OR
 					(reg_q1395 AND symb_decoder(16#59#)) OR
 					(reg_q1395 AND symb_decoder(16#b2#)) OR
 					(reg_q1395 AND symb_decoder(16#55#)) OR
 					(reg_q1395 AND symb_decoder(16#a9#)) OR
 					(reg_q1395 AND symb_decoder(16#a5#)) OR
 					(reg_q1395 AND symb_decoder(16#82#)) OR
 					(reg_q1395 AND symb_decoder(16#92#)) OR
 					(reg_q1395 AND symb_decoder(16#28#)) OR
 					(reg_q1395 AND symb_decoder(16#21#)) OR
 					(reg_q1395 AND symb_decoder(16#9a#)) OR
 					(reg_q1395 AND symb_decoder(16#41#)) OR
 					(reg_q1395 AND symb_decoder(16#0e#)) OR
 					(reg_q1395 AND symb_decoder(16#48#)) OR
 					(reg_q1395 AND symb_decoder(16#76#));
reg_q1395_init <= '0' ;
	p_reg_q1395: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1395 <= reg_q1395_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1395 <= reg_q1395_init;
        else
          reg_q1395 <= reg_q1395_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q516_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q516 AND symb_decoder(16#e7#)) OR
 					(reg_q516 AND symb_decoder(16#09#)) OR
 					(reg_q516 AND symb_decoder(16#88#)) OR
 					(reg_q516 AND symb_decoder(16#61#)) OR
 					(reg_q516 AND symb_decoder(16#46#)) OR
 					(reg_q516 AND symb_decoder(16#10#)) OR
 					(reg_q516 AND symb_decoder(16#fc#)) OR
 					(reg_q516 AND symb_decoder(16#e9#)) OR
 					(reg_q516 AND symb_decoder(16#08#)) OR
 					(reg_q516 AND symb_decoder(16#ca#)) OR
 					(reg_q516 AND symb_decoder(16#3c#)) OR
 					(reg_q516 AND symb_decoder(16#b8#)) OR
 					(reg_q516 AND symb_decoder(16#b9#)) OR
 					(reg_q516 AND symb_decoder(16#a0#)) OR
 					(reg_q516 AND symb_decoder(16#59#)) OR
 					(reg_q516 AND symb_decoder(16#2e#)) OR
 					(reg_q516 AND symb_decoder(16#e4#)) OR
 					(reg_q516 AND symb_decoder(16#11#)) OR
 					(reg_q516 AND symb_decoder(16#ac#)) OR
 					(reg_q516 AND symb_decoder(16#7b#)) OR
 					(reg_q516 AND symb_decoder(16#9d#)) OR
 					(reg_q516 AND symb_decoder(16#00#)) OR
 					(reg_q516 AND symb_decoder(16#49#)) OR
 					(reg_q516 AND symb_decoder(16#8e#)) OR
 					(reg_q516 AND symb_decoder(16#b4#)) OR
 					(reg_q516 AND symb_decoder(16#97#)) OR
 					(reg_q516 AND symb_decoder(16#04#)) OR
 					(reg_q516 AND symb_decoder(16#54#)) OR
 					(reg_q516 AND symb_decoder(16#b7#)) OR
 					(reg_q516 AND symb_decoder(16#bb#)) OR
 					(reg_q516 AND symb_decoder(16#a5#)) OR
 					(reg_q516 AND symb_decoder(16#c2#)) OR
 					(reg_q516 AND symb_decoder(16#f1#)) OR
 					(reg_q516 AND symb_decoder(16#78#)) OR
 					(reg_q516 AND symb_decoder(16#e8#)) OR
 					(reg_q516 AND symb_decoder(16#b1#)) OR
 					(reg_q516 AND symb_decoder(16#e1#)) OR
 					(reg_q516 AND symb_decoder(16#f2#)) OR
 					(reg_q516 AND symb_decoder(16#f6#)) OR
 					(reg_q516 AND symb_decoder(16#4b#)) OR
 					(reg_q516 AND symb_decoder(16#5d#)) OR
 					(reg_q516 AND symb_decoder(16#79#)) OR
 					(reg_q516 AND symb_decoder(16#ea#)) OR
 					(reg_q516 AND symb_decoder(16#72#)) OR
 					(reg_q516 AND symb_decoder(16#c8#)) OR
 					(reg_q516 AND symb_decoder(16#75#)) OR
 					(reg_q516 AND symb_decoder(16#48#)) OR
 					(reg_q516 AND symb_decoder(16#86#)) OR
 					(reg_q516 AND symb_decoder(16#67#)) OR
 					(reg_q516 AND symb_decoder(16#6a#)) OR
 					(reg_q516 AND symb_decoder(16#f3#)) OR
 					(reg_q516 AND symb_decoder(16#95#)) OR
 					(reg_q516 AND symb_decoder(16#65#)) OR
 					(reg_q516 AND symb_decoder(16#df#)) OR
 					(reg_q516 AND symb_decoder(16#29#)) OR
 					(reg_q516 AND symb_decoder(16#f5#)) OR
 					(reg_q516 AND symb_decoder(16#1f#)) OR
 					(reg_q516 AND symb_decoder(16#40#)) OR
 					(reg_q516 AND symb_decoder(16#36#)) OR
 					(reg_q516 AND symb_decoder(16#63#)) OR
 					(reg_q516 AND symb_decoder(16#bd#)) OR
 					(reg_q516 AND symb_decoder(16#ef#)) OR
 					(reg_q516 AND symb_decoder(16#2f#)) OR
 					(reg_q516 AND symb_decoder(16#e0#)) OR
 					(reg_q516 AND symb_decoder(16#de#)) OR
 					(reg_q516 AND symb_decoder(16#8b#)) OR
 					(reg_q516 AND symb_decoder(16#83#)) OR
 					(reg_q516 AND symb_decoder(16#2a#)) OR
 					(reg_q516 AND symb_decoder(16#da#)) OR
 					(reg_q516 AND symb_decoder(16#1e#)) OR
 					(reg_q516 AND symb_decoder(16#c0#)) OR
 					(reg_q516 AND symb_decoder(16#fe#)) OR
 					(reg_q516 AND symb_decoder(16#c4#)) OR
 					(reg_q516 AND symb_decoder(16#55#)) OR
 					(reg_q516 AND symb_decoder(16#fb#)) OR
 					(reg_q516 AND symb_decoder(16#b5#)) OR
 					(reg_q516 AND symb_decoder(16#16#)) OR
 					(reg_q516 AND symb_decoder(16#c5#)) OR
 					(reg_q516 AND symb_decoder(16#51#)) OR
 					(reg_q516 AND symb_decoder(16#42#)) OR
 					(reg_q516 AND symb_decoder(16#db#)) OR
 					(reg_q516 AND symb_decoder(16#06#)) OR
 					(reg_q516 AND symb_decoder(16#23#)) OR
 					(reg_q516 AND symb_decoder(16#ff#)) OR
 					(reg_q516 AND symb_decoder(16#1a#)) OR
 					(reg_q516 AND symb_decoder(16#2b#)) OR
 					(reg_q516 AND symb_decoder(16#3a#)) OR
 					(reg_q516 AND symb_decoder(16#7a#)) OR
 					(reg_q516 AND symb_decoder(16#76#)) OR
 					(reg_q516 AND symb_decoder(16#f0#)) OR
 					(reg_q516 AND symb_decoder(16#d9#)) OR
 					(reg_q516 AND symb_decoder(16#0a#)) OR
 					(reg_q516 AND symb_decoder(16#1b#)) OR
 					(reg_q516 AND symb_decoder(16#5b#)) OR
 					(reg_q516 AND symb_decoder(16#6f#)) OR
 					(reg_q516 AND symb_decoder(16#fa#)) OR
 					(reg_q516 AND symb_decoder(16#b2#)) OR
 					(reg_q516 AND symb_decoder(16#f4#)) OR
 					(reg_q516 AND symb_decoder(16#0b#)) OR
 					(reg_q516 AND symb_decoder(16#58#)) OR
 					(reg_q516 AND symb_decoder(16#57#)) OR
 					(reg_q516 AND symb_decoder(16#0d#)) OR
 					(reg_q516 AND symb_decoder(16#96#)) OR
 					(reg_q516 AND symb_decoder(16#94#)) OR
 					(reg_q516 AND symb_decoder(16#4c#)) OR
 					(reg_q516 AND symb_decoder(16#b6#)) OR
 					(reg_q516 AND symb_decoder(16#25#)) OR
 					(reg_q516 AND symb_decoder(16#66#)) OR
 					(reg_q516 AND symb_decoder(16#a4#)) OR
 					(reg_q516 AND symb_decoder(16#6c#)) OR
 					(reg_q516 AND symb_decoder(16#53#)) OR
 					(reg_q516 AND symb_decoder(16#ee#)) OR
 					(reg_q516 AND symb_decoder(16#b0#)) OR
 					(reg_q516 AND symb_decoder(16#50#)) OR
 					(reg_q516 AND symb_decoder(16#27#)) OR
 					(reg_q516 AND symb_decoder(16#8a#)) OR
 					(reg_q516 AND symb_decoder(16#5e#)) OR
 					(reg_q516 AND symb_decoder(16#d8#)) OR
 					(reg_q516 AND symb_decoder(16#99#)) OR
 					(reg_q516 AND symb_decoder(16#68#)) OR
 					(reg_q516 AND symb_decoder(16#ab#)) OR
 					(reg_q516 AND symb_decoder(16#85#)) OR
 					(reg_q516 AND symb_decoder(16#a7#)) OR
 					(reg_q516 AND symb_decoder(16#03#)) OR
 					(reg_q516 AND symb_decoder(16#ad#)) OR
 					(reg_q516 AND symb_decoder(16#ec#)) OR
 					(reg_q516 AND symb_decoder(16#74#)) OR
 					(reg_q516 AND symb_decoder(16#22#)) OR
 					(reg_q516 AND symb_decoder(16#ba#)) OR
 					(reg_q516 AND symb_decoder(16#8d#)) OR
 					(reg_q516 AND symb_decoder(16#ae#)) OR
 					(reg_q516 AND symb_decoder(16#a3#)) OR
 					(reg_q516 AND symb_decoder(16#93#)) OR
 					(reg_q516 AND symb_decoder(16#e3#)) OR
 					(reg_q516 AND symb_decoder(16#cc#)) OR
 					(reg_q516 AND symb_decoder(16#9c#)) OR
 					(reg_q516 AND symb_decoder(16#c7#)) OR
 					(reg_q516 AND symb_decoder(16#3b#)) OR
 					(reg_q516 AND symb_decoder(16#bc#)) OR
 					(reg_q516 AND symb_decoder(16#3f#)) OR
 					(reg_q516 AND symb_decoder(16#37#)) OR
 					(reg_q516 AND symb_decoder(16#77#)) OR
 					(reg_q516 AND symb_decoder(16#7f#)) OR
 					(reg_q516 AND symb_decoder(16#47#)) OR
 					(reg_q516 AND symb_decoder(16#e2#)) OR
 					(reg_q516 AND symb_decoder(16#bf#)) OR
 					(reg_q516 AND symb_decoder(16#9a#)) OR
 					(reg_q516 AND symb_decoder(16#80#)) OR
 					(reg_q516 AND symb_decoder(16#a9#)) OR
 					(reg_q516 AND symb_decoder(16#45#)) OR
 					(reg_q516 AND symb_decoder(16#5c#)) OR
 					(reg_q516 AND symb_decoder(16#71#)) OR
 					(reg_q516 AND symb_decoder(16#fd#)) OR
 					(reg_q516 AND symb_decoder(16#6e#)) OR
 					(reg_q516 AND symb_decoder(16#81#)) OR
 					(reg_q516 AND symb_decoder(16#dd#)) OR
 					(reg_q516 AND symb_decoder(16#6d#)) OR
 					(reg_q516 AND symb_decoder(16#64#)) OR
 					(reg_q516 AND symb_decoder(16#4e#)) OR
 					(reg_q516 AND symb_decoder(16#d0#)) OR
 					(reg_q516 AND symb_decoder(16#af#)) OR
 					(reg_q516 AND symb_decoder(16#f7#)) OR
 					(reg_q516 AND symb_decoder(16#17#)) OR
 					(reg_q516 AND symb_decoder(16#90#)) OR
 					(reg_q516 AND symb_decoder(16#8c#)) OR
 					(reg_q516 AND symb_decoder(16#31#)) OR
 					(reg_q516 AND symb_decoder(16#0e#)) OR
 					(reg_q516 AND symb_decoder(16#92#)) OR
 					(reg_q516 AND symb_decoder(16#26#)) OR
 					(reg_q516 AND symb_decoder(16#d3#)) OR
 					(reg_q516 AND symb_decoder(16#d5#)) OR
 					(reg_q516 AND symb_decoder(16#d1#)) OR
 					(reg_q516 AND symb_decoder(16#a2#)) OR
 					(reg_q516 AND symb_decoder(16#a8#)) OR
 					(reg_q516 AND symb_decoder(16#84#)) OR
 					(reg_q516 AND symb_decoder(16#be#)) OR
 					(reg_q516 AND symb_decoder(16#1d#)) OR
 					(reg_q516 AND symb_decoder(16#4d#)) OR
 					(reg_q516 AND symb_decoder(16#33#)) OR
 					(reg_q516 AND symb_decoder(16#d7#)) OR
 					(reg_q516 AND symb_decoder(16#56#)) OR
 					(reg_q516 AND symb_decoder(16#05#)) OR
 					(reg_q516 AND symb_decoder(16#5a#)) OR
 					(reg_q516 AND symb_decoder(16#20#)) OR
 					(reg_q516 AND symb_decoder(16#f9#)) OR
 					(reg_q516 AND symb_decoder(16#02#)) OR
 					(reg_q516 AND symb_decoder(16#98#)) OR
 					(reg_q516 AND symb_decoder(16#44#)) OR
 					(reg_q516 AND symb_decoder(16#a6#)) OR
 					(reg_q516 AND symb_decoder(16#43#)) OR
 					(reg_q516 AND symb_decoder(16#dc#)) OR
 					(reg_q516 AND symb_decoder(16#39#)) OR
 					(reg_q516 AND symb_decoder(16#2c#)) OR
 					(reg_q516 AND symb_decoder(16#28#)) OR
 					(reg_q516 AND symb_decoder(16#62#)) OR
 					(reg_q516 AND symb_decoder(16#18#)) OR
 					(reg_q516 AND symb_decoder(16#c9#)) OR
 					(reg_q516 AND symb_decoder(16#ce#)) OR
 					(reg_q516 AND symb_decoder(16#9b#)) OR
 					(reg_q516 AND symb_decoder(16#3e#)) OR
 					(reg_q516 AND symb_decoder(16#aa#)) OR
 					(reg_q516 AND symb_decoder(16#eb#)) OR
 					(reg_q516 AND symb_decoder(16#cd#)) OR
 					(reg_q516 AND symb_decoder(16#cf#)) OR
 					(reg_q516 AND symb_decoder(16#87#)) OR
 					(reg_q516 AND symb_decoder(16#e5#)) OR
 					(reg_q516 AND symb_decoder(16#5f#)) OR
 					(reg_q516 AND symb_decoder(16#52#)) OR
 					(reg_q516 AND symb_decoder(16#69#)) OR
 					(reg_q516 AND symb_decoder(16#4a#)) OR
 					(reg_q516 AND symb_decoder(16#3d#)) OR
 					(reg_q516 AND symb_decoder(16#01#)) OR
 					(reg_q516 AND symb_decoder(16#4f#)) OR
 					(reg_q516 AND symb_decoder(16#7d#)) OR
 					(reg_q516 AND symb_decoder(16#21#)) OR
 					(reg_q516 AND symb_decoder(16#d4#)) OR
 					(reg_q516 AND symb_decoder(16#15#)) OR
 					(reg_q516 AND symb_decoder(16#a1#)) OR
 					(reg_q516 AND symb_decoder(16#35#)) OR
 					(reg_q516 AND symb_decoder(16#19#)) OR
 					(reg_q516 AND symb_decoder(16#9f#)) OR
 					(reg_q516 AND symb_decoder(16#cb#)) OR
 					(reg_q516 AND symb_decoder(16#89#)) OR
 					(reg_q516 AND symb_decoder(16#d6#)) OR
 					(reg_q516 AND symb_decoder(16#14#)) OR
 					(reg_q516 AND symb_decoder(16#32#)) OR
 					(reg_q516 AND symb_decoder(16#70#)) OR
 					(reg_q516 AND symb_decoder(16#f8#)) OR
 					(reg_q516 AND symb_decoder(16#2d#)) OR
 					(reg_q516 AND symb_decoder(16#c6#)) OR
 					(reg_q516 AND symb_decoder(16#8f#)) OR
 					(reg_q516 AND symb_decoder(16#0c#)) OR
 					(reg_q516 AND symb_decoder(16#d2#)) OR
 					(reg_q516 AND symb_decoder(16#0f#)) OR
 					(reg_q516 AND symb_decoder(16#13#)) OR
 					(reg_q516 AND symb_decoder(16#c3#)) OR
 					(reg_q516 AND symb_decoder(16#12#)) OR
 					(reg_q516 AND symb_decoder(16#7e#)) OR
 					(reg_q516 AND symb_decoder(16#34#)) OR
 					(reg_q516 AND symb_decoder(16#60#)) OR
 					(reg_q516 AND symb_decoder(16#82#)) OR
 					(reg_q516 AND symb_decoder(16#30#)) OR
 					(reg_q516 AND symb_decoder(16#41#)) OR
 					(reg_q516 AND symb_decoder(16#38#)) OR
 					(reg_q516 AND symb_decoder(16#07#)) OR
 					(reg_q516 AND symb_decoder(16#91#)) OR
 					(reg_q516 AND symb_decoder(16#c1#)) OR
 					(reg_q516 AND symb_decoder(16#73#)) OR
 					(reg_q516 AND symb_decoder(16#7c#)) OR
 					(reg_q516 AND symb_decoder(16#6b#)) OR
 					(reg_q516 AND symb_decoder(16#24#)) OR
 					(reg_q516 AND symb_decoder(16#ed#)) OR
 					(reg_q516 AND symb_decoder(16#e6#)) OR
 					(reg_q516 AND symb_decoder(16#9e#)) OR
 					(reg_q516 AND symb_decoder(16#b3#)) OR
 					(reg_q516 AND symb_decoder(16#1c#));
reg_q516_init <= '0' ;
	p_reg_q516: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q516 <= reg_q516_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q516 <= reg_q516_init;
        else
          reg_q516 <= reg_q516_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1 AND symb_decoder(16#7b#)) OR
 					(reg_q1 AND symb_decoder(16#ed#)) OR
 					(reg_q1 AND symb_decoder(16#c2#)) OR
 					(reg_q1 AND symb_decoder(16#b1#)) OR
 					(reg_q1 AND symb_decoder(16#32#)) OR
 					(reg_q1 AND symb_decoder(16#11#)) OR
 					(reg_q1 AND symb_decoder(16#51#)) OR
 					(reg_q1 AND symb_decoder(16#d5#)) OR
 					(reg_q1 AND symb_decoder(16#e2#)) OR
 					(reg_q1 AND symb_decoder(16#bf#)) OR
 					(reg_q1 AND symb_decoder(16#cc#)) OR
 					(reg_q1 AND symb_decoder(16#34#)) OR
 					(reg_q1 AND symb_decoder(16#77#)) OR
 					(reg_q1 AND symb_decoder(16#4d#)) OR
 					(reg_q1 AND symb_decoder(16#29#)) OR
 					(reg_q1 AND symb_decoder(16#c7#)) OR
 					(reg_q1 AND symb_decoder(16#ef#)) OR
 					(reg_q1 AND symb_decoder(16#93#)) OR
 					(reg_q1 AND symb_decoder(16#d7#)) OR
 					(reg_q1 AND symb_decoder(16#91#)) OR
 					(reg_q1 AND symb_decoder(16#8a#)) OR
 					(reg_q1 AND symb_decoder(16#57#)) OR
 					(reg_q1 AND symb_decoder(16#c6#)) OR
 					(reg_q1 AND symb_decoder(16#88#)) OR
 					(reg_q1 AND symb_decoder(16#e1#)) OR
 					(reg_q1 AND symb_decoder(16#7e#)) OR
 					(reg_q1 AND symb_decoder(16#66#)) OR
 					(reg_q1 AND symb_decoder(16#e6#)) OR
 					(reg_q1 AND symb_decoder(16#f7#)) OR
 					(reg_q1 AND symb_decoder(16#d0#)) OR
 					(reg_q1 AND symb_decoder(16#40#)) OR
 					(reg_q1 AND symb_decoder(16#b2#)) OR
 					(reg_q1 AND symb_decoder(16#52#)) OR
 					(reg_q1 AND symb_decoder(16#24#)) OR
 					(reg_q1 AND symb_decoder(16#6b#)) OR
 					(reg_q1 AND symb_decoder(16#cf#)) OR
 					(reg_q1 AND symb_decoder(16#75#)) OR
 					(reg_q1 AND symb_decoder(16#37#)) OR
 					(reg_q1 AND symb_decoder(16#06#)) OR
 					(reg_q1 AND symb_decoder(16#b8#)) OR
 					(reg_q1 AND symb_decoder(16#4f#)) OR
 					(reg_q1 AND symb_decoder(16#85#)) OR
 					(reg_q1 AND symb_decoder(16#1f#)) OR
 					(reg_q1 AND symb_decoder(16#ec#)) OR
 					(reg_q1 AND symb_decoder(16#5b#)) OR
 					(reg_q1 AND symb_decoder(16#13#)) OR
 					(reg_q1 AND symb_decoder(16#6a#)) OR
 					(reg_q1 AND symb_decoder(16#17#)) OR
 					(reg_q1 AND symb_decoder(16#a0#)) OR
 					(reg_q1 AND symb_decoder(16#eb#)) OR
 					(reg_q1 AND symb_decoder(16#36#)) OR
 					(reg_q1 AND symb_decoder(16#9c#)) OR
 					(reg_q1 AND symb_decoder(16#15#)) OR
 					(reg_q1 AND symb_decoder(16#61#)) OR
 					(reg_q1 AND symb_decoder(16#78#)) OR
 					(reg_q1 AND symb_decoder(16#79#)) OR
 					(reg_q1 AND symb_decoder(16#2d#)) OR
 					(reg_q1 AND symb_decoder(16#42#)) OR
 					(reg_q1 AND symb_decoder(16#71#)) OR
 					(reg_q1 AND symb_decoder(16#e8#)) OR
 					(reg_q1 AND symb_decoder(16#82#)) OR
 					(reg_q1 AND symb_decoder(16#74#)) OR
 					(reg_q1 AND symb_decoder(16#0d#)) OR
 					(reg_q1 AND symb_decoder(16#02#)) OR
 					(reg_q1 AND symb_decoder(16#5c#)) OR
 					(reg_q1 AND symb_decoder(16#bb#)) OR
 					(reg_q1 AND symb_decoder(16#8e#)) OR
 					(reg_q1 AND symb_decoder(16#10#)) OR
 					(reg_q1 AND symb_decoder(16#5f#)) OR
 					(reg_q1 AND symb_decoder(16#f3#)) OR
 					(reg_q1 AND symb_decoder(16#d4#)) OR
 					(reg_q1 AND symb_decoder(16#1d#)) OR
 					(reg_q1 AND symb_decoder(16#4e#)) OR
 					(reg_q1 AND symb_decoder(16#ba#)) OR
 					(reg_q1 AND symb_decoder(16#76#)) OR
 					(reg_q1 AND symb_decoder(16#fc#)) OR
 					(reg_q1 AND symb_decoder(16#ee#)) OR
 					(reg_q1 AND symb_decoder(16#0a#)) OR
 					(reg_q1 AND symb_decoder(16#0f#)) OR
 					(reg_q1 AND symb_decoder(16#3f#)) OR
 					(reg_q1 AND symb_decoder(16#7f#)) OR
 					(reg_q1 AND symb_decoder(16#69#)) OR
 					(reg_q1 AND symb_decoder(16#55#)) OR
 					(reg_q1 AND symb_decoder(16#f4#)) OR
 					(reg_q1 AND symb_decoder(16#d8#)) OR
 					(reg_q1 AND symb_decoder(16#14#)) OR
 					(reg_q1 AND symb_decoder(16#4b#)) OR
 					(reg_q1 AND symb_decoder(16#27#)) OR
 					(reg_q1 AND symb_decoder(16#83#)) OR
 					(reg_q1 AND symb_decoder(16#38#)) OR
 					(reg_q1 AND symb_decoder(16#58#)) OR
 					(reg_q1 AND symb_decoder(16#da#)) OR
 					(reg_q1 AND symb_decoder(16#0e#)) OR
 					(reg_q1 AND symb_decoder(16#39#)) OR
 					(reg_q1 AND symb_decoder(16#ac#)) OR
 					(reg_q1 AND symb_decoder(16#2b#)) OR
 					(reg_q1 AND symb_decoder(16#16#)) OR
 					(reg_q1 AND symb_decoder(16#67#)) OR
 					(reg_q1 AND symb_decoder(16#5e#)) OR
 					(reg_q1 AND symb_decoder(16#22#)) OR
 					(reg_q1 AND symb_decoder(16#1b#)) OR
 					(reg_q1 AND symb_decoder(16#95#)) OR
 					(reg_q1 AND symb_decoder(16#df#)) OR
 					(reg_q1 AND symb_decoder(16#8b#)) OR
 					(reg_q1 AND symb_decoder(16#98#)) OR
 					(reg_q1 AND symb_decoder(16#c4#)) OR
 					(reg_q1 AND symb_decoder(16#68#)) OR
 					(reg_q1 AND symb_decoder(16#9f#)) OR
 					(reg_q1 AND symb_decoder(16#9d#)) OR
 					(reg_q1 AND symb_decoder(16#45#)) OR
 					(reg_q1 AND symb_decoder(16#8d#)) OR
 					(reg_q1 AND symb_decoder(16#00#)) OR
 					(reg_q1 AND symb_decoder(16#fe#)) OR
 					(reg_q1 AND symb_decoder(16#b4#)) OR
 					(reg_q1 AND symb_decoder(16#86#)) OR
 					(reg_q1 AND symb_decoder(16#d3#)) OR
 					(reg_q1 AND symb_decoder(16#5d#)) OR
 					(reg_q1 AND symb_decoder(16#43#)) OR
 					(reg_q1 AND symb_decoder(16#fd#)) OR
 					(reg_q1 AND symb_decoder(16#dc#)) OR
 					(reg_q1 AND symb_decoder(16#81#)) OR
 					(reg_q1 AND symb_decoder(16#c1#)) OR
 					(reg_q1 AND symb_decoder(16#c8#)) OR
 					(reg_q1 AND symb_decoder(16#84#)) OR
 					(reg_q1 AND symb_decoder(16#a1#)) OR
 					(reg_q1 AND symb_decoder(16#62#)) OR
 					(reg_q1 AND symb_decoder(16#f2#)) OR
 					(reg_q1 AND symb_decoder(16#09#)) OR
 					(reg_q1 AND symb_decoder(16#a5#)) OR
 					(reg_q1 AND symb_decoder(16#50#)) OR
 					(reg_q1 AND symb_decoder(16#9b#)) OR
 					(reg_q1 AND symb_decoder(16#d1#)) OR
 					(reg_q1 AND symb_decoder(16#0b#)) OR
 					(reg_q1 AND symb_decoder(16#a2#)) OR
 					(reg_q1 AND symb_decoder(16#8f#)) OR
 					(reg_q1 AND symb_decoder(16#97#)) OR
 					(reg_q1 AND symb_decoder(16#ae#)) OR
 					(reg_q1 AND symb_decoder(16#7c#)) OR
 					(reg_q1 AND symb_decoder(16#90#)) OR
 					(reg_q1 AND symb_decoder(16#dd#)) OR
 					(reg_q1 AND symb_decoder(16#7d#)) OR
 					(reg_q1 AND symb_decoder(16#3c#)) OR
 					(reg_q1 AND symb_decoder(16#7a#)) OR
 					(reg_q1 AND symb_decoder(16#f5#)) OR
 					(reg_q1 AND symb_decoder(16#21#)) OR
 					(reg_q1 AND symb_decoder(16#87#)) OR
 					(reg_q1 AND symb_decoder(16#6f#)) OR
 					(reg_q1 AND symb_decoder(16#56#)) OR
 					(reg_q1 AND symb_decoder(16#a7#)) OR
 					(reg_q1 AND symb_decoder(16#12#)) OR
 					(reg_q1 AND symb_decoder(16#23#)) OR
 					(reg_q1 AND symb_decoder(16#fa#)) OR
 					(reg_q1 AND symb_decoder(16#2a#)) OR
 					(reg_q1 AND symb_decoder(16#60#)) OR
 					(reg_q1 AND symb_decoder(16#30#)) OR
 					(reg_q1 AND symb_decoder(16#04#)) OR
 					(reg_q1 AND symb_decoder(16#73#)) OR
 					(reg_q1 AND symb_decoder(16#48#)) OR
 					(reg_q1 AND symb_decoder(16#01#)) OR
 					(reg_q1 AND symb_decoder(16#a9#)) OR
 					(reg_q1 AND symb_decoder(16#33#)) OR
 					(reg_q1 AND symb_decoder(16#2c#)) OR
 					(reg_q1 AND symb_decoder(16#3e#)) OR
 					(reg_q1 AND symb_decoder(16#3b#)) OR
 					(reg_q1 AND symb_decoder(16#4a#)) OR
 					(reg_q1 AND symb_decoder(16#ce#)) OR
 					(reg_q1 AND symb_decoder(16#2e#)) OR
 					(reg_q1 AND symb_decoder(16#f1#)) OR
 					(reg_q1 AND symb_decoder(16#59#)) OR
 					(reg_q1 AND symb_decoder(16#54#)) OR
 					(reg_q1 AND symb_decoder(16#e7#)) OR
 					(reg_q1 AND symb_decoder(16#9a#)) OR
 					(reg_q1 AND symb_decoder(16#e4#)) OR
 					(reg_q1 AND symb_decoder(16#26#)) OR
 					(reg_q1 AND symb_decoder(16#a6#)) OR
 					(reg_q1 AND symb_decoder(16#cd#)) OR
 					(reg_q1 AND symb_decoder(16#63#)) OR
 					(reg_q1 AND symb_decoder(16#89#)) OR
 					(reg_q1 AND symb_decoder(16#3a#)) OR
 					(reg_q1 AND symb_decoder(16#f0#)) OR
 					(reg_q1 AND symb_decoder(16#1e#)) OR
 					(reg_q1 AND symb_decoder(16#a3#)) OR
 					(reg_q1 AND symb_decoder(16#6c#)) OR
 					(reg_q1 AND symb_decoder(16#d2#)) OR
 					(reg_q1 AND symb_decoder(16#b9#)) OR
 					(reg_q1 AND symb_decoder(16#03#)) OR
 					(reg_q1 AND symb_decoder(16#db#)) OR
 					(reg_q1 AND symb_decoder(16#28#)) OR
 					(reg_q1 AND symb_decoder(16#d6#)) OR
 					(reg_q1 AND symb_decoder(16#ff#)) OR
 					(reg_q1 AND symb_decoder(16#af#)) OR
 					(reg_q1 AND symb_decoder(16#5a#)) OR
 					(reg_q1 AND symb_decoder(16#bd#)) OR
 					(reg_q1 AND symb_decoder(16#aa#)) OR
 					(reg_q1 AND symb_decoder(16#99#)) OR
 					(reg_q1 AND symb_decoder(16#c0#)) OR
 					(reg_q1 AND symb_decoder(16#9e#)) OR
 					(reg_q1 AND symb_decoder(16#05#)) OR
 					(reg_q1 AND symb_decoder(16#31#)) OR
 					(reg_q1 AND symb_decoder(16#2f#)) OR
 					(reg_q1 AND symb_decoder(16#19#)) OR
 					(reg_q1 AND symb_decoder(16#ea#)) OR
 					(reg_q1 AND symb_decoder(16#80#)) OR
 					(reg_q1 AND symb_decoder(16#65#)) OR
 					(reg_q1 AND symb_decoder(16#a8#)) OR
 					(reg_q1 AND symb_decoder(16#72#)) OR
 					(reg_q1 AND symb_decoder(16#53#)) OR
 					(reg_q1 AND symb_decoder(16#c5#)) OR
 					(reg_q1 AND symb_decoder(16#94#)) OR
 					(reg_q1 AND symb_decoder(16#25#)) OR
 					(reg_q1 AND symb_decoder(16#be#)) OR
 					(reg_q1 AND symb_decoder(16#6e#)) OR
 					(reg_q1 AND symb_decoder(16#41#)) OR
 					(reg_q1 AND symb_decoder(16#64#)) OR
 					(reg_q1 AND symb_decoder(16#35#)) OR
 					(reg_q1 AND symb_decoder(16#c3#)) OR
 					(reg_q1 AND symb_decoder(16#96#)) OR
 					(reg_q1 AND symb_decoder(16#46#)) OR
 					(reg_q1 AND symb_decoder(16#47#)) OR
 					(reg_q1 AND symb_decoder(16#f8#)) OR
 					(reg_q1 AND symb_decoder(16#44#)) OR
 					(reg_q1 AND symb_decoder(16#f6#)) OR
 					(reg_q1 AND symb_decoder(16#ab#)) OR
 					(reg_q1 AND symb_decoder(16#f9#)) OR
 					(reg_q1 AND symb_decoder(16#b6#)) OR
 					(reg_q1 AND symb_decoder(16#4c#)) OR
 					(reg_q1 AND symb_decoder(16#d9#)) OR
 					(reg_q1 AND symb_decoder(16#b0#)) OR
 					(reg_q1 AND symb_decoder(16#e5#)) OR
 					(reg_q1 AND symb_decoder(16#18#)) OR
 					(reg_q1 AND symb_decoder(16#92#)) OR
 					(reg_q1 AND symb_decoder(16#cb#)) OR
 					(reg_q1 AND symb_decoder(16#07#)) OR
 					(reg_q1 AND symb_decoder(16#e3#)) OR
 					(reg_q1 AND symb_decoder(16#a4#)) OR
 					(reg_q1 AND symb_decoder(16#b5#)) OR
 					(reg_q1 AND symb_decoder(16#70#)) OR
 					(reg_q1 AND symb_decoder(16#c9#)) OR
 					(reg_q1 AND symb_decoder(16#6d#)) OR
 					(reg_q1 AND symb_decoder(16#fb#)) OR
 					(reg_q1 AND symb_decoder(16#49#)) OR
 					(reg_q1 AND symb_decoder(16#e9#)) OR
 					(reg_q1 AND symb_decoder(16#0c#)) OR
 					(reg_q1 AND symb_decoder(16#ca#)) OR
 					(reg_q1 AND symb_decoder(16#e0#)) OR
 					(reg_q1 AND symb_decoder(16#1c#)) OR
 					(reg_q1 AND symb_decoder(16#bc#)) OR
 					(reg_q1 AND symb_decoder(16#08#)) OR
 					(reg_q1 AND symb_decoder(16#b7#)) OR
 					(reg_q1 AND symb_decoder(16#8c#)) OR
 					(reg_q1 AND symb_decoder(16#3d#)) OR
 					(reg_q1 AND symb_decoder(16#20#)) OR
 					(reg_q1 AND symb_decoder(16#ad#)) OR
 					(reg_q1 AND symb_decoder(16#de#)) OR
 					(reg_q1 AND symb_decoder(16#1a#)) OR
 					(reg_q1 AND symb_decoder(16#b3#));
reg_q1_init <= '0' ;
	p_reg_q1: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1 <= reg_q1_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1 <= reg_q1_init;
        else
          reg_q1 <= reg_q1_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2556_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q2556 AND symb_decoder(16#db#)) OR
 					(reg_q2556 AND symb_decoder(16#8c#)) OR
 					(reg_q2556 AND symb_decoder(16#ab#)) OR
 					(reg_q2556 AND symb_decoder(16#e2#)) OR
 					(reg_q2556 AND symb_decoder(16#67#)) OR
 					(reg_q2556 AND symb_decoder(16#09#)) OR
 					(reg_q2556 AND symb_decoder(16#1e#)) OR
 					(reg_q2556 AND symb_decoder(16#11#)) OR
 					(reg_q2556 AND symb_decoder(16#24#)) OR
 					(reg_q2556 AND symb_decoder(16#dd#)) OR
 					(reg_q2556 AND symb_decoder(16#35#)) OR
 					(reg_q2556 AND symb_decoder(16#c0#)) OR
 					(reg_q2556 AND symb_decoder(16#1d#)) OR
 					(reg_q2556 AND symb_decoder(16#5a#)) OR
 					(reg_q2556 AND symb_decoder(16#89#)) OR
 					(reg_q2556 AND symb_decoder(16#29#)) OR
 					(reg_q2556 AND symb_decoder(16#fc#)) OR
 					(reg_q2556 AND symb_decoder(16#5f#)) OR
 					(reg_q2556 AND symb_decoder(16#55#)) OR
 					(reg_q2556 AND symb_decoder(16#0d#)) OR
 					(reg_q2556 AND symb_decoder(16#e4#)) OR
 					(reg_q2556 AND symb_decoder(16#4f#)) OR
 					(reg_q2556 AND symb_decoder(16#1a#)) OR
 					(reg_q2556 AND symb_decoder(16#0b#)) OR
 					(reg_q2556 AND symb_decoder(16#c1#)) OR
 					(reg_q2556 AND symb_decoder(16#0a#)) OR
 					(reg_q2556 AND symb_decoder(16#71#)) OR
 					(reg_q2556 AND symb_decoder(16#b7#)) OR
 					(reg_q2556 AND symb_decoder(16#ce#)) OR
 					(reg_q2556 AND symb_decoder(16#cd#)) OR
 					(reg_q2556 AND symb_decoder(16#f9#)) OR
 					(reg_q2556 AND symb_decoder(16#ff#)) OR
 					(reg_q2556 AND symb_decoder(16#d7#)) OR
 					(reg_q2556 AND symb_decoder(16#82#)) OR
 					(reg_q2556 AND symb_decoder(16#10#)) OR
 					(reg_q2556 AND symb_decoder(16#69#)) OR
 					(reg_q2556 AND symb_decoder(16#0f#)) OR
 					(reg_q2556 AND symb_decoder(16#b5#)) OR
 					(reg_q2556 AND symb_decoder(16#af#)) OR
 					(reg_q2556 AND symb_decoder(16#80#)) OR
 					(reg_q2556 AND symb_decoder(16#bd#)) OR
 					(reg_q2556 AND symb_decoder(16#88#)) OR
 					(reg_q2556 AND symb_decoder(16#53#)) OR
 					(reg_q2556 AND symb_decoder(16#f0#)) OR
 					(reg_q2556 AND symb_decoder(16#31#)) OR
 					(reg_q2556 AND symb_decoder(16#77#)) OR
 					(reg_q2556 AND symb_decoder(16#64#)) OR
 					(reg_q2556 AND symb_decoder(16#02#)) OR
 					(reg_q2556 AND symb_decoder(16#12#)) OR
 					(reg_q2556 AND symb_decoder(16#ac#)) OR
 					(reg_q2556 AND symb_decoder(16#8e#)) OR
 					(reg_q2556 AND symb_decoder(16#aa#)) OR
 					(reg_q2556 AND symb_decoder(16#9c#)) OR
 					(reg_q2556 AND symb_decoder(16#8f#)) OR
 					(reg_q2556 AND symb_decoder(16#59#)) OR
 					(reg_q2556 AND symb_decoder(16#95#)) OR
 					(reg_q2556 AND symb_decoder(16#c9#)) OR
 					(reg_q2556 AND symb_decoder(16#6b#)) OR
 					(reg_q2556 AND symb_decoder(16#cb#)) OR
 					(reg_q2556 AND symb_decoder(16#be#)) OR
 					(reg_q2556 AND symb_decoder(16#c3#)) OR
 					(reg_q2556 AND symb_decoder(16#18#)) OR
 					(reg_q2556 AND symb_decoder(16#e7#)) OR
 					(reg_q2556 AND symb_decoder(16#7f#)) OR
 					(reg_q2556 AND symb_decoder(16#2f#)) OR
 					(reg_q2556 AND symb_decoder(16#e5#)) OR
 					(reg_q2556 AND symb_decoder(16#93#)) OR
 					(reg_q2556 AND symb_decoder(16#5e#)) OR
 					(reg_q2556 AND symb_decoder(16#b2#)) OR
 					(reg_q2556 AND symb_decoder(16#d8#)) OR
 					(reg_q2556 AND symb_decoder(16#3d#)) OR
 					(reg_q2556 AND symb_decoder(16#3a#)) OR
 					(reg_q2556 AND symb_decoder(16#e6#)) OR
 					(reg_q2556 AND symb_decoder(16#4b#)) OR
 					(reg_q2556 AND symb_decoder(16#97#)) OR
 					(reg_q2556 AND symb_decoder(16#6c#)) OR
 					(reg_q2556 AND symb_decoder(16#c2#)) OR
 					(reg_q2556 AND symb_decoder(16#44#)) OR
 					(reg_q2556 AND symb_decoder(16#cf#)) OR
 					(reg_q2556 AND symb_decoder(16#1f#)) OR
 					(reg_q2556 AND symb_decoder(16#cc#)) OR
 					(reg_q2556 AND symb_decoder(16#66#)) OR
 					(reg_q2556 AND symb_decoder(16#01#)) OR
 					(reg_q2556 AND symb_decoder(16#fd#)) OR
 					(reg_q2556 AND symb_decoder(16#8a#)) OR
 					(reg_q2556 AND symb_decoder(16#fb#)) OR
 					(reg_q2556 AND symb_decoder(16#2e#)) OR
 					(reg_q2556 AND symb_decoder(16#98#)) OR
 					(reg_q2556 AND symb_decoder(16#96#)) OR
 					(reg_q2556 AND symb_decoder(16#13#)) OR
 					(reg_q2556 AND symb_decoder(16#3f#)) OR
 					(reg_q2556 AND symb_decoder(16#21#)) OR
 					(reg_q2556 AND symb_decoder(16#d2#)) OR
 					(reg_q2556 AND symb_decoder(16#17#)) OR
 					(reg_q2556 AND symb_decoder(16#bf#)) OR
 					(reg_q2556 AND symb_decoder(16#48#)) OR
 					(reg_q2556 AND symb_decoder(16#81#)) OR
 					(reg_q2556 AND symb_decoder(16#54#)) OR
 					(reg_q2556 AND symb_decoder(16#c8#)) OR
 					(reg_q2556 AND symb_decoder(16#15#)) OR
 					(reg_q2556 AND symb_decoder(16#5b#)) OR
 					(reg_q2556 AND symb_decoder(16#9f#)) OR
 					(reg_q2556 AND symb_decoder(16#b1#)) OR
 					(reg_q2556 AND symb_decoder(16#99#)) OR
 					(reg_q2556 AND symb_decoder(16#26#)) OR
 					(reg_q2556 AND symb_decoder(16#49#)) OR
 					(reg_q2556 AND symb_decoder(16#a0#)) OR
 					(reg_q2556 AND symb_decoder(16#61#)) OR
 					(reg_q2556 AND symb_decoder(16#43#)) OR
 					(reg_q2556 AND symb_decoder(16#a4#)) OR
 					(reg_q2556 AND symb_decoder(16#45#)) OR
 					(reg_q2556 AND symb_decoder(16#6d#)) OR
 					(reg_q2556 AND symb_decoder(16#d3#)) OR
 					(reg_q2556 AND symb_decoder(16#08#)) OR
 					(reg_q2556 AND symb_decoder(16#df#)) OR
 					(reg_q2556 AND symb_decoder(16#68#)) OR
 					(reg_q2556 AND symb_decoder(16#a8#)) OR
 					(reg_q2556 AND symb_decoder(16#e1#)) OR
 					(reg_q2556 AND symb_decoder(16#23#)) OR
 					(reg_q2556 AND symb_decoder(16#47#)) OR
 					(reg_q2556 AND symb_decoder(16#84#)) OR
 					(reg_q2556 AND symb_decoder(16#8d#)) OR
 					(reg_q2556 AND symb_decoder(16#92#)) OR
 					(reg_q2556 AND symb_decoder(16#d9#)) OR
 					(reg_q2556 AND symb_decoder(16#51#)) OR
 					(reg_q2556 AND symb_decoder(16#1b#)) OR
 					(reg_q2556 AND symb_decoder(16#c7#)) OR
 					(reg_q2556 AND symb_decoder(16#d0#)) OR
 					(reg_q2556 AND symb_decoder(16#2b#)) OR
 					(reg_q2556 AND symb_decoder(16#d5#)) OR
 					(reg_q2556 AND symb_decoder(16#c4#)) OR
 					(reg_q2556 AND symb_decoder(16#3b#)) OR
 					(reg_q2556 AND symb_decoder(16#dc#)) OR
 					(reg_q2556 AND symb_decoder(16#28#)) OR
 					(reg_q2556 AND symb_decoder(16#30#)) OR
 					(reg_q2556 AND symb_decoder(16#f6#)) OR
 					(reg_q2556 AND symb_decoder(16#6a#)) OR
 					(reg_q2556 AND symb_decoder(16#7b#)) OR
 					(reg_q2556 AND symb_decoder(16#b3#)) OR
 					(reg_q2556 AND symb_decoder(16#03#)) OR
 					(reg_q2556 AND symb_decoder(16#9a#)) OR
 					(reg_q2556 AND symb_decoder(16#eb#)) OR
 					(reg_q2556 AND symb_decoder(16#32#)) OR
 					(reg_q2556 AND symb_decoder(16#91#)) OR
 					(reg_q2556 AND symb_decoder(16#a3#)) OR
 					(reg_q2556 AND symb_decoder(16#73#)) OR
 					(reg_q2556 AND symb_decoder(16#f1#)) OR
 					(reg_q2556 AND symb_decoder(16#56#)) OR
 					(reg_q2556 AND symb_decoder(16#76#)) OR
 					(reg_q2556 AND symb_decoder(16#7d#)) OR
 					(reg_q2556 AND symb_decoder(16#a5#)) OR
 					(reg_q2556 AND symb_decoder(16#3c#)) OR
 					(reg_q2556 AND symb_decoder(16#06#)) OR
 					(reg_q2556 AND symb_decoder(16#57#)) OR
 					(reg_q2556 AND symb_decoder(16#bb#)) OR
 					(reg_q2556 AND symb_decoder(16#f7#)) OR
 					(reg_q2556 AND symb_decoder(16#7a#)) OR
 					(reg_q2556 AND symb_decoder(16#d6#)) OR
 					(reg_q2556 AND symb_decoder(16#52#)) OR
 					(reg_q2556 AND symb_decoder(16#7e#)) OR
 					(reg_q2556 AND symb_decoder(16#c5#)) OR
 					(reg_q2556 AND symb_decoder(16#ea#)) OR
 					(reg_q2556 AND symb_decoder(16#f3#)) OR
 					(reg_q2556 AND symb_decoder(16#ee#)) OR
 					(reg_q2556 AND symb_decoder(16#62#)) OR
 					(reg_q2556 AND symb_decoder(16#b6#)) OR
 					(reg_q2556 AND symb_decoder(16#ad#)) OR
 					(reg_q2556 AND symb_decoder(16#ef#)) OR
 					(reg_q2556 AND symb_decoder(16#a9#)) OR
 					(reg_q2556 AND symb_decoder(16#a6#)) OR
 					(reg_q2556 AND symb_decoder(16#58#)) OR
 					(reg_q2556 AND symb_decoder(16#b0#)) OR
 					(reg_q2556 AND symb_decoder(16#38#)) OR
 					(reg_q2556 AND symb_decoder(16#f8#)) OR
 					(reg_q2556 AND symb_decoder(16#4a#)) OR
 					(reg_q2556 AND symb_decoder(16#05#)) OR
 					(reg_q2556 AND symb_decoder(16#41#)) OR
 					(reg_q2556 AND symb_decoder(16#40#)) OR
 					(reg_q2556 AND symb_decoder(16#8b#)) OR
 					(reg_q2556 AND symb_decoder(16#50#)) OR
 					(reg_q2556 AND symb_decoder(16#bc#)) OR
 					(reg_q2556 AND symb_decoder(16#c6#)) OR
 					(reg_q2556 AND symb_decoder(16#42#)) OR
 					(reg_q2556 AND symb_decoder(16#f5#)) OR
 					(reg_q2556 AND symb_decoder(16#2a#)) OR
 					(reg_q2556 AND symb_decoder(16#87#)) OR
 					(reg_q2556 AND symb_decoder(16#63#)) OR
 					(reg_q2556 AND symb_decoder(16#70#)) OR
 					(reg_q2556 AND symb_decoder(16#e0#)) OR
 					(reg_q2556 AND symb_decoder(16#4c#)) OR
 					(reg_q2556 AND symb_decoder(16#20#)) OR
 					(reg_q2556 AND symb_decoder(16#b4#)) OR
 					(reg_q2556 AND symb_decoder(16#a1#)) OR
 					(reg_q2556 AND symb_decoder(16#16#)) OR
 					(reg_q2556 AND symb_decoder(16#79#)) OR
 					(reg_q2556 AND symb_decoder(16#3e#)) OR
 					(reg_q2556 AND symb_decoder(16#83#)) OR
 					(reg_q2556 AND symb_decoder(16#ed#)) OR
 					(reg_q2556 AND symb_decoder(16#1c#)) OR
 					(reg_q2556 AND symb_decoder(16#7c#)) OR
 					(reg_q2556 AND symb_decoder(16#74#)) OR
 					(reg_q2556 AND symb_decoder(16#5c#)) OR
 					(reg_q2556 AND symb_decoder(16#d1#)) OR
 					(reg_q2556 AND symb_decoder(16#ae#)) OR
 					(reg_q2556 AND symb_decoder(16#4e#)) OR
 					(reg_q2556 AND symb_decoder(16#ba#)) OR
 					(reg_q2556 AND symb_decoder(16#37#)) OR
 					(reg_q2556 AND symb_decoder(16#14#)) OR
 					(reg_q2556 AND symb_decoder(16#e8#)) OR
 					(reg_q2556 AND symb_decoder(16#ec#)) OR
 					(reg_q2556 AND symb_decoder(16#94#)) OR
 					(reg_q2556 AND symb_decoder(16#b8#)) OR
 					(reg_q2556 AND symb_decoder(16#9d#)) OR
 					(reg_q2556 AND symb_decoder(16#04#)) OR
 					(reg_q2556 AND symb_decoder(16#25#)) OR
 					(reg_q2556 AND symb_decoder(16#36#)) OR
 					(reg_q2556 AND symb_decoder(16#00#)) OR
 					(reg_q2556 AND symb_decoder(16#0c#)) OR
 					(reg_q2556 AND symb_decoder(16#85#)) OR
 					(reg_q2556 AND symb_decoder(16#fe#)) OR
 					(reg_q2556 AND symb_decoder(16#78#)) OR
 					(reg_q2556 AND symb_decoder(16#34#)) OR
 					(reg_q2556 AND symb_decoder(16#4d#)) OR
 					(reg_q2556 AND symb_decoder(16#86#)) OR
 					(reg_q2556 AND symb_decoder(16#72#)) OR
 					(reg_q2556 AND symb_decoder(16#6e#)) OR
 					(reg_q2556 AND symb_decoder(16#ca#)) OR
 					(reg_q2556 AND symb_decoder(16#39#)) OR
 					(reg_q2556 AND symb_decoder(16#19#)) OR
 					(reg_q2556 AND symb_decoder(16#de#)) OR
 					(reg_q2556 AND symb_decoder(16#a7#)) OR
 					(reg_q2556 AND symb_decoder(16#07#)) OR
 					(reg_q2556 AND symb_decoder(16#f4#)) OR
 					(reg_q2556 AND symb_decoder(16#46#)) OR
 					(reg_q2556 AND symb_decoder(16#0e#)) OR
 					(reg_q2556 AND symb_decoder(16#f2#)) OR
 					(reg_q2556 AND symb_decoder(16#a2#)) OR
 					(reg_q2556 AND symb_decoder(16#60#)) OR
 					(reg_q2556 AND symb_decoder(16#27#)) OR
 					(reg_q2556 AND symb_decoder(16#22#)) OR
 					(reg_q2556 AND symb_decoder(16#65#)) OR
 					(reg_q2556 AND symb_decoder(16#90#)) OR
 					(reg_q2556 AND symb_decoder(16#2c#)) OR
 					(reg_q2556 AND symb_decoder(16#2d#)) OR
 					(reg_q2556 AND symb_decoder(16#da#)) OR
 					(reg_q2556 AND symb_decoder(16#b9#)) OR
 					(reg_q2556 AND symb_decoder(16#6f#)) OR
 					(reg_q2556 AND symb_decoder(16#e3#)) OR
 					(reg_q2556 AND symb_decoder(16#33#)) OR
 					(reg_q2556 AND symb_decoder(16#fa#)) OR
 					(reg_q2556 AND symb_decoder(16#9b#)) OR
 					(reg_q2556 AND symb_decoder(16#5d#)) OR
 					(reg_q2556 AND symb_decoder(16#75#)) OR
 					(reg_q2556 AND symb_decoder(16#9e#)) OR
 					(reg_q2556 AND symb_decoder(16#d4#)) OR
 					(reg_q2556 AND symb_decoder(16#e9#));
reg_q2556_init <= '0' ;
	p_reg_q2556: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2556 <= reg_q2556_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2556 <= reg_q2556_init;
        else
          reg_q2556 <= reg_q2556_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q399_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q399 AND symb_decoder(16#08#)) OR
 					(reg_q399 AND symb_decoder(16#00#)) OR
 					(reg_q399 AND symb_decoder(16#a1#)) OR
 					(reg_q399 AND symb_decoder(16#40#)) OR
 					(reg_q399 AND symb_decoder(16#42#)) OR
 					(reg_q399 AND symb_decoder(16#46#)) OR
 					(reg_q399 AND symb_decoder(16#f5#)) OR
 					(reg_q399 AND symb_decoder(16#8c#)) OR
 					(reg_q399 AND symb_decoder(16#c6#)) OR
 					(reg_q399 AND symb_decoder(16#92#)) OR
 					(reg_q399 AND symb_decoder(16#32#)) OR
 					(reg_q399 AND symb_decoder(16#e4#)) OR
 					(reg_q399 AND symb_decoder(16#90#)) OR
 					(reg_q399 AND symb_decoder(16#3f#)) OR
 					(reg_q399 AND symb_decoder(16#7a#)) OR
 					(reg_q399 AND symb_decoder(16#25#)) OR
 					(reg_q399 AND symb_decoder(16#b2#)) OR
 					(reg_q399 AND symb_decoder(16#06#)) OR
 					(reg_q399 AND symb_decoder(16#c5#)) OR
 					(reg_q399 AND symb_decoder(16#8d#)) OR
 					(reg_q399 AND symb_decoder(16#2f#)) OR
 					(reg_q399 AND symb_decoder(16#69#)) OR
 					(reg_q399 AND symb_decoder(16#f4#)) OR
 					(reg_q399 AND symb_decoder(16#7b#)) OR
 					(reg_q399 AND symb_decoder(16#5d#)) OR
 					(reg_q399 AND symb_decoder(16#33#)) OR
 					(reg_q399 AND symb_decoder(16#c3#)) OR
 					(reg_q399 AND symb_decoder(16#6e#)) OR
 					(reg_q399 AND symb_decoder(16#94#)) OR
 					(reg_q399 AND symb_decoder(16#d4#)) OR
 					(reg_q399 AND symb_decoder(16#2c#)) OR
 					(reg_q399 AND symb_decoder(16#57#)) OR
 					(reg_q399 AND symb_decoder(16#56#)) OR
 					(reg_q399 AND symb_decoder(16#96#)) OR
 					(reg_q399 AND symb_decoder(16#91#)) OR
 					(reg_q399 AND symb_decoder(16#a2#)) OR
 					(reg_q399 AND symb_decoder(16#cb#)) OR
 					(reg_q399 AND symb_decoder(16#77#)) OR
 					(reg_q399 AND symb_decoder(16#5c#)) OR
 					(reg_q399 AND symb_decoder(16#80#)) OR
 					(reg_q399 AND symb_decoder(16#6c#)) OR
 					(reg_q399 AND symb_decoder(16#1a#)) OR
 					(reg_q399 AND symb_decoder(16#f9#)) OR
 					(reg_q399 AND symb_decoder(16#b3#)) OR
 					(reg_q399 AND symb_decoder(16#45#)) OR
 					(reg_q399 AND symb_decoder(16#67#)) OR
 					(reg_q399 AND symb_decoder(16#4d#)) OR
 					(reg_q399 AND symb_decoder(16#f8#)) OR
 					(reg_q399 AND symb_decoder(16#1c#)) OR
 					(reg_q399 AND symb_decoder(16#ee#)) OR
 					(reg_q399 AND symb_decoder(16#e2#)) OR
 					(reg_q399 AND symb_decoder(16#20#)) OR
 					(reg_q399 AND symb_decoder(16#75#)) OR
 					(reg_q399 AND symb_decoder(16#ed#)) OR
 					(reg_q399 AND symb_decoder(16#0e#)) OR
 					(reg_q399 AND symb_decoder(16#e5#)) OR
 					(reg_q399 AND symb_decoder(16#ad#)) OR
 					(reg_q399 AND symb_decoder(16#31#)) OR
 					(reg_q399 AND symb_decoder(16#1d#)) OR
 					(reg_q399 AND symb_decoder(16#64#)) OR
 					(reg_q399 AND symb_decoder(16#58#)) OR
 					(reg_q399 AND symb_decoder(16#29#)) OR
 					(reg_q399 AND symb_decoder(16#2b#)) OR
 					(reg_q399 AND symb_decoder(16#cf#)) OR
 					(reg_q399 AND symb_decoder(16#bf#)) OR
 					(reg_q399 AND symb_decoder(16#68#)) OR
 					(reg_q399 AND symb_decoder(16#10#)) OR
 					(reg_q399 AND symb_decoder(16#fe#)) OR
 					(reg_q399 AND symb_decoder(16#53#)) OR
 					(reg_q399 AND symb_decoder(16#b7#)) OR
 					(reg_q399 AND symb_decoder(16#97#)) OR
 					(reg_q399 AND symb_decoder(16#72#)) OR
 					(reg_q399 AND symb_decoder(16#3e#)) OR
 					(reg_q399 AND symb_decoder(16#81#)) OR
 					(reg_q399 AND symb_decoder(16#8a#)) OR
 					(reg_q399 AND symb_decoder(16#a7#)) OR
 					(reg_q399 AND symb_decoder(16#d0#)) OR
 					(reg_q399 AND symb_decoder(16#5e#)) OR
 					(reg_q399 AND symb_decoder(16#d7#)) OR
 					(reg_q399 AND symb_decoder(16#0f#)) OR
 					(reg_q399 AND symb_decoder(16#24#)) OR
 					(reg_q399 AND symb_decoder(16#fd#)) OR
 					(reg_q399 AND symb_decoder(16#22#)) OR
 					(reg_q399 AND symb_decoder(16#39#)) OR
 					(reg_q399 AND symb_decoder(16#ec#)) OR
 					(reg_q399 AND symb_decoder(16#d8#)) OR
 					(reg_q399 AND symb_decoder(16#ce#)) OR
 					(reg_q399 AND symb_decoder(16#3c#)) OR
 					(reg_q399 AND symb_decoder(16#1e#)) OR
 					(reg_q399 AND symb_decoder(16#48#)) OR
 					(reg_q399 AND symb_decoder(16#5b#)) OR
 					(reg_q399 AND symb_decoder(16#82#)) OR
 					(reg_q399 AND symb_decoder(16#8b#)) OR
 					(reg_q399 AND symb_decoder(16#47#)) OR
 					(reg_q399 AND symb_decoder(16#3d#)) OR
 					(reg_q399 AND symb_decoder(16#19#)) OR
 					(reg_q399 AND symb_decoder(16#74#)) OR
 					(reg_q399 AND symb_decoder(16#df#)) OR
 					(reg_q399 AND symb_decoder(16#21#)) OR
 					(reg_q399 AND symb_decoder(16#55#)) OR
 					(reg_q399 AND symb_decoder(16#0b#)) OR
 					(reg_q399 AND symb_decoder(16#65#)) OR
 					(reg_q399 AND symb_decoder(16#99#)) OR
 					(reg_q399 AND symb_decoder(16#84#)) OR
 					(reg_q399 AND symb_decoder(16#93#)) OR
 					(reg_q399 AND symb_decoder(16#27#)) OR
 					(reg_q399 AND symb_decoder(16#de#)) OR
 					(reg_q399 AND symb_decoder(16#4e#)) OR
 					(reg_q399 AND symb_decoder(16#36#)) OR
 					(reg_q399 AND symb_decoder(16#a4#)) OR
 					(reg_q399 AND symb_decoder(16#85#)) OR
 					(reg_q399 AND symb_decoder(16#9c#)) OR
 					(reg_q399 AND symb_decoder(16#ef#)) OR
 					(reg_q399 AND symb_decoder(16#28#)) OR
 					(reg_q399 AND symb_decoder(16#e1#)) OR
 					(reg_q399 AND symb_decoder(16#88#)) OR
 					(reg_q399 AND symb_decoder(16#8e#)) OR
 					(reg_q399 AND symb_decoder(16#5a#)) OR
 					(reg_q399 AND symb_decoder(16#98#)) OR
 					(reg_q399 AND symb_decoder(16#ac#)) OR
 					(reg_q399 AND symb_decoder(16#2a#)) OR
 					(reg_q399 AND symb_decoder(16#60#)) OR
 					(reg_q399 AND symb_decoder(16#ba#)) OR
 					(reg_q399 AND symb_decoder(16#e0#)) OR
 					(reg_q399 AND symb_decoder(16#8f#)) OR
 					(reg_q399 AND symb_decoder(16#0d#)) OR
 					(reg_q399 AND symb_decoder(16#9e#)) OR
 					(reg_q399 AND symb_decoder(16#6a#)) OR
 					(reg_q399 AND symb_decoder(16#bb#)) OR
 					(reg_q399 AND symb_decoder(16#1f#)) OR
 					(reg_q399 AND symb_decoder(16#fb#)) OR
 					(reg_q399 AND symb_decoder(16#d9#)) OR
 					(reg_q399 AND symb_decoder(16#d6#)) OR
 					(reg_q399 AND symb_decoder(16#54#)) OR
 					(reg_q399 AND symb_decoder(16#f0#)) OR
 					(reg_q399 AND symb_decoder(16#5f#)) OR
 					(reg_q399 AND symb_decoder(16#b6#)) OR
 					(reg_q399 AND symb_decoder(16#bd#)) OR
 					(reg_q399 AND symb_decoder(16#c8#)) OR
 					(reg_q399 AND symb_decoder(16#4b#)) OR
 					(reg_q399 AND symb_decoder(16#76#)) OR
 					(reg_q399 AND symb_decoder(16#db#)) OR
 					(reg_q399 AND symb_decoder(16#d1#)) OR
 					(reg_q399 AND symb_decoder(16#2e#)) OR
 					(reg_q399 AND symb_decoder(16#50#)) OR
 					(reg_q399 AND symb_decoder(16#3a#)) OR
 					(reg_q399 AND symb_decoder(16#4c#)) OR
 					(reg_q399 AND symb_decoder(16#62#)) OR
 					(reg_q399 AND symb_decoder(16#f1#)) OR
 					(reg_q399 AND symb_decoder(16#b4#)) OR
 					(reg_q399 AND symb_decoder(16#f7#)) OR
 					(reg_q399 AND symb_decoder(16#c4#)) OR
 					(reg_q399 AND symb_decoder(16#13#)) OR
 					(reg_q399 AND symb_decoder(16#70#)) OR
 					(reg_q399 AND symb_decoder(16#e6#)) OR
 					(reg_q399 AND symb_decoder(16#38#)) OR
 					(reg_q399 AND symb_decoder(16#9b#)) OR
 					(reg_q399 AND symb_decoder(16#03#)) OR
 					(reg_q399 AND symb_decoder(16#e3#)) OR
 					(reg_q399 AND symb_decoder(16#23#)) OR
 					(reg_q399 AND symb_decoder(16#95#)) OR
 					(reg_q399 AND symb_decoder(16#9a#)) OR
 					(reg_q399 AND symb_decoder(16#37#)) OR
 					(reg_q399 AND symb_decoder(16#6b#)) OR
 					(reg_q399 AND symb_decoder(16#61#)) OR
 					(reg_q399 AND symb_decoder(16#a9#)) OR
 					(reg_q399 AND symb_decoder(16#b0#)) OR
 					(reg_q399 AND symb_decoder(16#02#)) OR
 					(reg_q399 AND symb_decoder(16#01#)) OR
 					(reg_q399 AND symb_decoder(16#44#)) OR
 					(reg_q399 AND symb_decoder(16#d5#)) OR
 					(reg_q399 AND symb_decoder(16#41#)) OR
 					(reg_q399 AND symb_decoder(16#07#)) OR
 					(reg_q399 AND symb_decoder(16#eb#)) OR
 					(reg_q399 AND symb_decoder(16#4a#)) OR
 					(reg_q399 AND symb_decoder(16#ae#)) OR
 					(reg_q399 AND symb_decoder(16#dd#)) OR
 					(reg_q399 AND symb_decoder(16#4f#)) OR
 					(reg_q399 AND symb_decoder(16#e8#)) OR
 					(reg_q399 AND symb_decoder(16#43#)) OR
 					(reg_q399 AND symb_decoder(16#fa#)) OR
 					(reg_q399 AND symb_decoder(16#34#)) OR
 					(reg_q399 AND symb_decoder(16#a8#)) OR
 					(reg_q399 AND symb_decoder(16#73#)) OR
 					(reg_q399 AND symb_decoder(16#17#)) OR
 					(reg_q399 AND symb_decoder(16#cd#)) OR
 					(reg_q399 AND symb_decoder(16#d3#)) OR
 					(reg_q399 AND symb_decoder(16#15#)) OR
 					(reg_q399 AND symb_decoder(16#89#)) OR
 					(reg_q399 AND symb_decoder(16#35#)) OR
 					(reg_q399 AND symb_decoder(16#f2#)) OR
 					(reg_q399 AND symb_decoder(16#2d#)) OR
 					(reg_q399 AND symb_decoder(16#b8#)) OR
 					(reg_q399 AND symb_decoder(16#83#)) OR
 					(reg_q399 AND symb_decoder(16#e7#)) OR
 					(reg_q399 AND symb_decoder(16#3b#)) OR
 					(reg_q399 AND symb_decoder(16#aa#)) OR
 					(reg_q399 AND symb_decoder(16#71#)) OR
 					(reg_q399 AND symb_decoder(16#79#)) OR
 					(reg_q399 AND symb_decoder(16#6f#)) OR
 					(reg_q399 AND symb_decoder(16#e9#)) OR
 					(reg_q399 AND symb_decoder(16#59#)) OR
 					(reg_q399 AND symb_decoder(16#f6#)) OR
 					(reg_q399 AND symb_decoder(16#49#)) OR
 					(reg_q399 AND symb_decoder(16#52#)) OR
 					(reg_q399 AND symb_decoder(16#ff#)) OR
 					(reg_q399 AND symb_decoder(16#a5#)) OR
 					(reg_q399 AND symb_decoder(16#86#)) OR
 					(reg_q399 AND symb_decoder(16#05#)) OR
 					(reg_q399 AND symb_decoder(16#ab#)) OR
 					(reg_q399 AND symb_decoder(16#7d#)) OR
 					(reg_q399 AND symb_decoder(16#9d#)) OR
 					(reg_q399 AND symb_decoder(16#fc#)) OR
 					(reg_q399 AND symb_decoder(16#af#)) OR
 					(reg_q399 AND symb_decoder(16#63#)) OR
 					(reg_q399 AND symb_decoder(16#0a#)) OR
 					(reg_q399 AND symb_decoder(16#1b#)) OR
 					(reg_q399 AND symb_decoder(16#a0#)) OR
 					(reg_q399 AND symb_decoder(16#7c#)) OR
 					(reg_q399 AND symb_decoder(16#ea#)) OR
 					(reg_q399 AND symb_decoder(16#51#)) OR
 					(reg_q399 AND symb_decoder(16#87#)) OR
 					(reg_q399 AND symb_decoder(16#6d#)) OR
 					(reg_q399 AND symb_decoder(16#7f#)) OR
 					(reg_q399 AND symb_decoder(16#c0#)) OR
 					(reg_q399 AND symb_decoder(16#30#)) OR
 					(reg_q399 AND symb_decoder(16#78#)) OR
 					(reg_q399 AND symb_decoder(16#b1#)) OR
 					(reg_q399 AND symb_decoder(16#c2#)) OR
 					(reg_q399 AND symb_decoder(16#9f#)) OR
 					(reg_q399 AND symb_decoder(16#c9#)) OR
 					(reg_q399 AND symb_decoder(16#b5#)) OR
 					(reg_q399 AND symb_decoder(16#cc#)) OR
 					(reg_q399 AND symb_decoder(16#a6#)) OR
 					(reg_q399 AND symb_decoder(16#0c#)) OR
 					(reg_q399 AND symb_decoder(16#12#)) OR
 					(reg_q399 AND symb_decoder(16#16#)) OR
 					(reg_q399 AND symb_decoder(16#ca#)) OR
 					(reg_q399 AND symb_decoder(16#d2#)) OR
 					(reg_q399 AND symb_decoder(16#04#)) OR
 					(reg_q399 AND symb_decoder(16#da#)) OR
 					(reg_q399 AND symb_decoder(16#be#)) OR
 					(reg_q399 AND symb_decoder(16#09#)) OR
 					(reg_q399 AND symb_decoder(16#14#)) OR
 					(reg_q399 AND symb_decoder(16#66#)) OR
 					(reg_q399 AND symb_decoder(16#f3#)) OR
 					(reg_q399 AND symb_decoder(16#dc#)) OR
 					(reg_q399 AND symb_decoder(16#26#)) OR
 					(reg_q399 AND symb_decoder(16#a3#)) OR
 					(reg_q399 AND symb_decoder(16#18#)) OR
 					(reg_q399 AND symb_decoder(16#bc#)) OR
 					(reg_q399 AND symb_decoder(16#c1#)) OR
 					(reg_q399 AND symb_decoder(16#b9#)) OR
 					(reg_q399 AND symb_decoder(16#11#)) OR
 					(reg_q399 AND symb_decoder(16#c7#)) OR
 					(reg_q399 AND symb_decoder(16#7e#));
reg_q399_init <= '0' ;
	p_reg_q399: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q399 <= reg_q399_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q399 <= reg_q399_init;
        else
          reg_q399 <= reg_q399_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1628_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1628 AND symb_decoder(16#9c#)) OR
 					(reg_q1628 AND symb_decoder(16#f5#)) OR
 					(reg_q1628 AND symb_decoder(16#4b#)) OR
 					(reg_q1628 AND symb_decoder(16#dd#)) OR
 					(reg_q1628 AND symb_decoder(16#22#)) OR
 					(reg_q1628 AND symb_decoder(16#53#)) OR
 					(reg_q1628 AND symb_decoder(16#50#)) OR
 					(reg_q1628 AND symb_decoder(16#17#)) OR
 					(reg_q1628 AND symb_decoder(16#9e#)) OR
 					(reg_q1628 AND symb_decoder(16#16#)) OR
 					(reg_q1628 AND symb_decoder(16#c9#)) OR
 					(reg_q1628 AND symb_decoder(16#79#)) OR
 					(reg_q1628 AND symb_decoder(16#be#)) OR
 					(reg_q1628 AND symb_decoder(16#d6#)) OR
 					(reg_q1628 AND symb_decoder(16#26#)) OR
 					(reg_q1628 AND symb_decoder(16#4e#)) OR
 					(reg_q1628 AND symb_decoder(16#88#)) OR
 					(reg_q1628 AND symb_decoder(16#21#)) OR
 					(reg_q1628 AND symb_decoder(16#83#)) OR
 					(reg_q1628 AND symb_decoder(16#61#)) OR
 					(reg_q1628 AND symb_decoder(16#48#)) OR
 					(reg_q1628 AND symb_decoder(16#47#)) OR
 					(reg_q1628 AND symb_decoder(16#11#)) OR
 					(reg_q1628 AND symb_decoder(16#5f#)) OR
 					(reg_q1628 AND symb_decoder(16#7e#)) OR
 					(reg_q1628 AND symb_decoder(16#06#)) OR
 					(reg_q1628 AND symb_decoder(16#07#)) OR
 					(reg_q1628 AND symb_decoder(16#ca#)) OR
 					(reg_q1628 AND symb_decoder(16#36#)) OR
 					(reg_q1628 AND symb_decoder(16#27#)) OR
 					(reg_q1628 AND symb_decoder(16#99#)) OR
 					(reg_q1628 AND symb_decoder(16#7b#)) OR
 					(reg_q1628 AND symb_decoder(16#d3#)) OR
 					(reg_q1628 AND symb_decoder(16#20#)) OR
 					(reg_q1628 AND symb_decoder(16#ef#)) OR
 					(reg_q1628 AND symb_decoder(16#72#)) OR
 					(reg_q1628 AND symb_decoder(16#30#)) OR
 					(reg_q1628 AND symb_decoder(16#a1#)) OR
 					(reg_q1628 AND symb_decoder(16#25#)) OR
 					(reg_q1628 AND symb_decoder(16#00#)) OR
 					(reg_q1628 AND symb_decoder(16#fa#)) OR
 					(reg_q1628 AND symb_decoder(16#1e#)) OR
 					(reg_q1628 AND symb_decoder(16#70#)) OR
 					(reg_q1628 AND symb_decoder(16#66#)) OR
 					(reg_q1628 AND symb_decoder(16#1d#)) OR
 					(reg_q1628 AND symb_decoder(16#ba#)) OR
 					(reg_q1628 AND symb_decoder(16#b3#)) OR
 					(reg_q1628 AND symb_decoder(16#3a#)) OR
 					(reg_q1628 AND symb_decoder(16#52#)) OR
 					(reg_q1628 AND symb_decoder(16#f3#)) OR
 					(reg_q1628 AND symb_decoder(16#d1#)) OR
 					(reg_q1628 AND symb_decoder(16#73#)) OR
 					(reg_q1628 AND symb_decoder(16#42#)) OR
 					(reg_q1628 AND symb_decoder(16#4a#)) OR
 					(reg_q1628 AND symb_decoder(16#46#)) OR
 					(reg_q1628 AND symb_decoder(16#7c#)) OR
 					(reg_q1628 AND symb_decoder(16#e7#)) OR
 					(reg_q1628 AND symb_decoder(16#68#)) OR
 					(reg_q1628 AND symb_decoder(16#85#)) OR
 					(reg_q1628 AND symb_decoder(16#55#)) OR
 					(reg_q1628 AND symb_decoder(16#c1#)) OR
 					(reg_q1628 AND symb_decoder(16#f1#)) OR
 					(reg_q1628 AND symb_decoder(16#5a#)) OR
 					(reg_q1628 AND symb_decoder(16#3c#)) OR
 					(reg_q1628 AND symb_decoder(16#8a#)) OR
 					(reg_q1628 AND symb_decoder(16#0b#)) OR
 					(reg_q1628 AND symb_decoder(16#9a#)) OR
 					(reg_q1628 AND symb_decoder(16#bf#)) OR
 					(reg_q1628 AND symb_decoder(16#45#)) OR
 					(reg_q1628 AND symb_decoder(16#78#)) OR
 					(reg_q1628 AND symb_decoder(16#f9#)) OR
 					(reg_q1628 AND symb_decoder(16#d9#)) OR
 					(reg_q1628 AND symb_decoder(16#e4#)) OR
 					(reg_q1628 AND symb_decoder(16#74#)) OR
 					(reg_q1628 AND symb_decoder(16#59#)) OR
 					(reg_q1628 AND symb_decoder(16#aa#)) OR
 					(reg_q1628 AND symb_decoder(16#e6#)) OR
 					(reg_q1628 AND symb_decoder(16#6a#)) OR
 					(reg_q1628 AND symb_decoder(16#e1#)) OR
 					(reg_q1628 AND symb_decoder(16#39#)) OR
 					(reg_q1628 AND symb_decoder(16#08#)) OR
 					(reg_q1628 AND symb_decoder(16#a3#)) OR
 					(reg_q1628 AND symb_decoder(16#0d#)) OR
 					(reg_q1628 AND symb_decoder(16#40#)) OR
 					(reg_q1628 AND symb_decoder(16#da#)) OR
 					(reg_q1628 AND symb_decoder(16#12#)) OR
 					(reg_q1628 AND symb_decoder(16#a8#)) OR
 					(reg_q1628 AND symb_decoder(16#1a#)) OR
 					(reg_q1628 AND symb_decoder(16#e2#)) OR
 					(reg_q1628 AND symb_decoder(16#18#)) OR
 					(reg_q1628 AND symb_decoder(16#cc#)) OR
 					(reg_q1628 AND symb_decoder(16#af#)) OR
 					(reg_q1628 AND symb_decoder(16#c0#)) OR
 					(reg_q1628 AND symb_decoder(16#63#)) OR
 					(reg_q1628 AND symb_decoder(16#ad#)) OR
 					(reg_q1628 AND symb_decoder(16#19#)) OR
 					(reg_q1628 AND symb_decoder(16#ff#)) OR
 					(reg_q1628 AND symb_decoder(16#3d#)) OR
 					(reg_q1628 AND symb_decoder(16#05#)) OR
 					(reg_q1628 AND symb_decoder(16#f8#)) OR
 					(reg_q1628 AND symb_decoder(16#d8#)) OR
 					(reg_q1628 AND symb_decoder(16#bb#)) OR
 					(reg_q1628 AND symb_decoder(16#bd#)) OR
 					(reg_q1628 AND symb_decoder(16#0a#)) OR
 					(reg_q1628 AND symb_decoder(16#f7#)) OR
 					(reg_q1628 AND symb_decoder(16#1b#)) OR
 					(reg_q1628 AND symb_decoder(16#b7#)) OR
 					(reg_q1628 AND symb_decoder(16#94#)) OR
 					(reg_q1628 AND symb_decoder(16#5e#)) OR
 					(reg_q1628 AND symb_decoder(16#96#)) OR
 					(reg_q1628 AND symb_decoder(16#b0#)) OR
 					(reg_q1628 AND symb_decoder(16#fb#)) OR
 					(reg_q1628 AND symb_decoder(16#fc#)) OR
 					(reg_q1628 AND symb_decoder(16#4d#)) OR
 					(reg_q1628 AND symb_decoder(16#6c#)) OR
 					(reg_q1628 AND symb_decoder(16#0c#)) OR
 					(reg_q1628 AND symb_decoder(16#c7#)) OR
 					(reg_q1628 AND symb_decoder(16#95#)) OR
 					(reg_q1628 AND symb_decoder(16#de#)) OR
 					(reg_q1628 AND symb_decoder(16#33#)) OR
 					(reg_q1628 AND symb_decoder(16#fd#)) OR
 					(reg_q1628 AND symb_decoder(16#97#)) OR
 					(reg_q1628 AND symb_decoder(16#ac#)) OR
 					(reg_q1628 AND symb_decoder(16#37#)) OR
 					(reg_q1628 AND symb_decoder(16#41#)) OR
 					(reg_q1628 AND symb_decoder(16#c4#)) OR
 					(reg_q1628 AND symb_decoder(16#3e#)) OR
 					(reg_q1628 AND symb_decoder(16#db#)) OR
 					(reg_q1628 AND symb_decoder(16#7a#)) OR
 					(reg_q1628 AND symb_decoder(16#0e#)) OR
 					(reg_q1628 AND symb_decoder(16#a4#)) OR
 					(reg_q1628 AND symb_decoder(16#4f#)) OR
 					(reg_q1628 AND symb_decoder(16#c3#)) OR
 					(reg_q1628 AND symb_decoder(16#ce#)) OR
 					(reg_q1628 AND symb_decoder(16#5c#)) OR
 					(reg_q1628 AND symb_decoder(16#28#)) OR
 					(reg_q1628 AND symb_decoder(16#3f#)) OR
 					(reg_q1628 AND symb_decoder(16#d0#)) OR
 					(reg_q1628 AND symb_decoder(16#2c#)) OR
 					(reg_q1628 AND symb_decoder(16#ec#)) OR
 					(reg_q1628 AND symb_decoder(16#13#)) OR
 					(reg_q1628 AND symb_decoder(16#14#)) OR
 					(reg_q1628 AND symb_decoder(16#77#)) OR
 					(reg_q1628 AND symb_decoder(16#29#)) OR
 					(reg_q1628 AND symb_decoder(16#e0#)) OR
 					(reg_q1628 AND symb_decoder(16#d4#)) OR
 					(reg_q1628 AND symb_decoder(16#75#)) OR
 					(reg_q1628 AND symb_decoder(16#90#)) OR
 					(reg_q1628 AND symb_decoder(16#02#)) OR
 					(reg_q1628 AND symb_decoder(16#44#)) OR
 					(reg_q1628 AND symb_decoder(16#0f#)) OR
 					(reg_q1628 AND symb_decoder(16#e3#)) OR
 					(reg_q1628 AND symb_decoder(16#65#)) OR
 					(reg_q1628 AND symb_decoder(16#6e#)) OR
 					(reg_q1628 AND symb_decoder(16#b1#)) OR
 					(reg_q1628 AND symb_decoder(16#8d#)) OR
 					(reg_q1628 AND symb_decoder(16#32#)) OR
 					(reg_q1628 AND symb_decoder(16#8f#)) OR
 					(reg_q1628 AND symb_decoder(16#76#)) OR
 					(reg_q1628 AND symb_decoder(16#9f#)) OR
 					(reg_q1628 AND symb_decoder(16#ab#)) OR
 					(reg_q1628 AND symb_decoder(16#04#)) OR
 					(reg_q1628 AND symb_decoder(16#5d#)) OR
 					(reg_q1628 AND symb_decoder(16#81#)) OR
 					(reg_q1628 AND symb_decoder(16#b6#)) OR
 					(reg_q1628 AND symb_decoder(16#5b#)) OR
 					(reg_q1628 AND symb_decoder(16#62#)) OR
 					(reg_q1628 AND symb_decoder(16#ee#)) OR
 					(reg_q1628 AND symb_decoder(16#e8#)) OR
 					(reg_q1628 AND symb_decoder(16#6f#)) OR
 					(reg_q1628 AND symb_decoder(16#34#)) OR
 					(reg_q1628 AND symb_decoder(16#57#)) OR
 					(reg_q1628 AND symb_decoder(16#80#)) OR
 					(reg_q1628 AND symb_decoder(16#a7#)) OR
 					(reg_q1628 AND symb_decoder(16#f6#)) OR
 					(reg_q1628 AND symb_decoder(16#b8#)) OR
 					(reg_q1628 AND symb_decoder(16#2b#)) OR
 					(reg_q1628 AND symb_decoder(16#1c#)) OR
 					(reg_q1628 AND symb_decoder(16#dc#)) OR
 					(reg_q1628 AND symb_decoder(16#cd#)) OR
 					(reg_q1628 AND symb_decoder(16#51#)) OR
 					(reg_q1628 AND symb_decoder(16#e9#)) OR
 					(reg_q1628 AND symb_decoder(16#fe#)) OR
 					(reg_q1628 AND symb_decoder(16#67#)) OR
 					(reg_q1628 AND symb_decoder(16#2f#)) OR
 					(reg_q1628 AND symb_decoder(16#df#)) OR
 					(reg_q1628 AND symb_decoder(16#15#)) OR
 					(reg_q1628 AND symb_decoder(16#89#)) OR
 					(reg_q1628 AND symb_decoder(16#54#)) OR
 					(reg_q1628 AND symb_decoder(16#d5#)) OR
 					(reg_q1628 AND symb_decoder(16#9b#)) OR
 					(reg_q1628 AND symb_decoder(16#eb#)) OR
 					(reg_q1628 AND symb_decoder(16#49#)) OR
 					(reg_q1628 AND symb_decoder(16#c6#)) OR
 					(reg_q1628 AND symb_decoder(16#64#)) OR
 					(reg_q1628 AND symb_decoder(16#58#)) OR
 					(reg_q1628 AND symb_decoder(16#24#)) OR
 					(reg_q1628 AND symb_decoder(16#01#)) OR
 					(reg_q1628 AND symb_decoder(16#35#)) OR
 					(reg_q1628 AND symb_decoder(16#ea#)) OR
 					(reg_q1628 AND symb_decoder(16#f0#)) OR
 					(reg_q1628 AND symb_decoder(16#23#)) OR
 					(reg_q1628 AND symb_decoder(16#10#)) OR
 					(reg_q1628 AND symb_decoder(16#a6#)) OR
 					(reg_q1628 AND symb_decoder(16#2e#)) OR
 					(reg_q1628 AND symb_decoder(16#ae#)) OR
 					(reg_q1628 AND symb_decoder(16#c2#)) OR
 					(reg_q1628 AND symb_decoder(16#6d#)) OR
 					(reg_q1628 AND symb_decoder(16#60#)) OR
 					(reg_q1628 AND symb_decoder(16#b9#)) OR
 					(reg_q1628 AND symb_decoder(16#98#)) OR
 					(reg_q1628 AND symb_decoder(16#c8#)) OR
 					(reg_q1628 AND symb_decoder(16#31#)) OR
 					(reg_q1628 AND symb_decoder(16#84#)) OR
 					(reg_q1628 AND symb_decoder(16#b2#)) OR
 					(reg_q1628 AND symb_decoder(16#4c#)) OR
 					(reg_q1628 AND symb_decoder(16#c5#)) OR
 					(reg_q1628 AND symb_decoder(16#92#)) OR
 					(reg_q1628 AND symb_decoder(16#2d#)) OR
 					(reg_q1628 AND symb_decoder(16#87#)) OR
 					(reg_q1628 AND symb_decoder(16#8c#)) OR
 					(reg_q1628 AND symb_decoder(16#82#)) OR
 					(reg_q1628 AND symb_decoder(16#9d#)) OR
 					(reg_q1628 AND symb_decoder(16#7f#)) OR
 					(reg_q1628 AND symb_decoder(16#91#)) OR
 					(reg_q1628 AND symb_decoder(16#d7#)) OR
 					(reg_q1628 AND symb_decoder(16#a0#)) OR
 					(reg_q1628 AND symb_decoder(16#71#)) OR
 					(reg_q1628 AND symb_decoder(16#2a#)) OR
 					(reg_q1628 AND symb_decoder(16#cf#)) OR
 					(reg_q1628 AND symb_decoder(16#7d#)) OR
 					(reg_q1628 AND symb_decoder(16#b5#)) OR
 					(reg_q1628 AND symb_decoder(16#09#)) OR
 					(reg_q1628 AND symb_decoder(16#86#)) OR
 					(reg_q1628 AND symb_decoder(16#a9#)) OR
 					(reg_q1628 AND symb_decoder(16#1f#)) OR
 					(reg_q1628 AND symb_decoder(16#93#)) OR
 					(reg_q1628 AND symb_decoder(16#a5#)) OR
 					(reg_q1628 AND symb_decoder(16#8b#)) OR
 					(reg_q1628 AND symb_decoder(16#d2#)) OR
 					(reg_q1628 AND symb_decoder(16#b4#)) OR
 					(reg_q1628 AND symb_decoder(16#6b#)) OR
 					(reg_q1628 AND symb_decoder(16#f4#)) OR
 					(reg_q1628 AND symb_decoder(16#bc#)) OR
 					(reg_q1628 AND symb_decoder(16#ed#)) OR
 					(reg_q1628 AND symb_decoder(16#56#)) OR
 					(reg_q1628 AND symb_decoder(16#8e#)) OR
 					(reg_q1628 AND symb_decoder(16#cb#)) OR
 					(reg_q1628 AND symb_decoder(16#43#)) OR
 					(reg_q1628 AND symb_decoder(16#3b#)) OR
 					(reg_q1628 AND symb_decoder(16#38#)) OR
 					(reg_q1628 AND symb_decoder(16#03#)) OR
 					(reg_q1628 AND symb_decoder(16#69#)) OR
 					(reg_q1628 AND symb_decoder(16#a2#)) OR
 					(reg_q1628 AND symb_decoder(16#e5#)) OR
 					(reg_q1628 AND symb_decoder(16#f2#));
reg_q1628_init <= '0' ;
	p_reg_q1628: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1628 <= reg_q1628_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1628 <= reg_q1628_init;
        else
          reg_q1628 <= reg_q1628_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2552_in <= (reg_q2534 AND symb_decoder(16#d0#)) OR
 					(reg_q2534 AND symb_decoder(16#3b#)) OR
 					(reg_q2534 AND symb_decoder(16#c7#)) OR
 					(reg_q2534 AND symb_decoder(16#f7#)) OR
 					(reg_q2534 AND symb_decoder(16#b5#)) OR
 					(reg_q2534 AND symb_decoder(16#44#)) OR
 					(reg_q2534 AND symb_decoder(16#9b#)) OR
 					(reg_q2534 AND symb_decoder(16#83#)) OR
 					(reg_q2534 AND symb_decoder(16#c8#)) OR
 					(reg_q2534 AND symb_decoder(16#bc#)) OR
 					(reg_q2534 AND symb_decoder(16#3a#)) OR
 					(reg_q2534 AND symb_decoder(16#30#)) OR
 					(reg_q2534 AND symb_decoder(16#fb#)) OR
 					(reg_q2534 AND symb_decoder(16#7f#)) OR
 					(reg_q2534 AND symb_decoder(16#6d#)) OR
 					(reg_q2534 AND symb_decoder(16#3d#)) OR
 					(reg_q2534 AND symb_decoder(16#20#)) OR
 					(reg_q2534 AND symb_decoder(16#9a#)) OR
 					(reg_q2534 AND symb_decoder(16#79#)) OR
 					(reg_q2534 AND symb_decoder(16#7c#)) OR
 					(reg_q2534 AND symb_decoder(16#33#)) OR
 					(reg_q2534 AND symb_decoder(16#d4#)) OR
 					(reg_q2534 AND symb_decoder(16#00#)) OR
 					(reg_q2534 AND symb_decoder(16#5c#)) OR
 					(reg_q2534 AND symb_decoder(16#ef#)) OR
 					(reg_q2534 AND symb_decoder(16#11#)) OR
 					(reg_q2534 AND symb_decoder(16#f1#)) OR
 					(reg_q2534 AND symb_decoder(16#94#)) OR
 					(reg_q2534 AND symb_decoder(16#46#)) OR
 					(reg_q2534 AND symb_decoder(16#eb#)) OR
 					(reg_q2534 AND symb_decoder(16#13#)) OR
 					(reg_q2534 AND symb_decoder(16#8a#)) OR
 					(reg_q2534 AND symb_decoder(16#21#)) OR
 					(reg_q2534 AND symb_decoder(16#0b#)) OR
 					(reg_q2534 AND symb_decoder(16#74#)) OR
 					(reg_q2534 AND symb_decoder(16#bb#)) OR
 					(reg_q2534 AND symb_decoder(16#fd#)) OR
 					(reg_q2534 AND symb_decoder(16#97#)) OR
 					(reg_q2534 AND symb_decoder(16#a1#)) OR
 					(reg_q2534 AND symb_decoder(16#ad#)) OR
 					(reg_q2534 AND symb_decoder(16#37#)) OR
 					(reg_q2534 AND symb_decoder(16#2f#)) OR
 					(reg_q2534 AND symb_decoder(16#b9#)) OR
 					(reg_q2534 AND symb_decoder(16#f2#)) OR
 					(reg_q2534 AND symb_decoder(16#fc#)) OR
 					(reg_q2534 AND symb_decoder(16#17#)) OR
 					(reg_q2534 AND symb_decoder(16#0e#)) OR
 					(reg_q2534 AND symb_decoder(16#ca#)) OR
 					(reg_q2534 AND symb_decoder(16#7d#)) OR
 					(reg_q2534 AND symb_decoder(16#2c#)) OR
 					(reg_q2534 AND symb_decoder(16#ae#)) OR
 					(reg_q2534 AND symb_decoder(16#48#)) OR
 					(reg_q2534 AND symb_decoder(16#93#)) OR
 					(reg_q2534 AND symb_decoder(16#aa#)) OR
 					(reg_q2534 AND symb_decoder(16#65#)) OR
 					(reg_q2534 AND symb_decoder(16#a6#)) OR
 					(reg_q2534 AND symb_decoder(16#54#)) OR
 					(reg_q2534 AND symb_decoder(16#ff#)) OR
 					(reg_q2534 AND symb_decoder(16#0d#)) OR
 					(reg_q2534 AND symb_decoder(16#09#)) OR
 					(reg_q2534 AND symb_decoder(16#07#)) OR
 					(reg_q2534 AND symb_decoder(16#ac#)) OR
 					(reg_q2534 AND symb_decoder(16#da#)) OR
 					(reg_q2534 AND symb_decoder(16#95#)) OR
 					(reg_q2534 AND symb_decoder(16#15#)) OR
 					(reg_q2534 AND symb_decoder(16#8b#)) OR
 					(reg_q2534 AND symb_decoder(16#d6#)) OR
 					(reg_q2534 AND symb_decoder(16#de#)) OR
 					(reg_q2534 AND symb_decoder(16#39#)) OR
 					(reg_q2534 AND symb_decoder(16#cd#)) OR
 					(reg_q2534 AND symb_decoder(16#96#)) OR
 					(reg_q2534 AND symb_decoder(16#9c#)) OR
 					(reg_q2534 AND symb_decoder(16#53#)) OR
 					(reg_q2534 AND symb_decoder(16#d8#)) OR
 					(reg_q2534 AND symb_decoder(16#56#)) OR
 					(reg_q2534 AND symb_decoder(16#58#)) OR
 					(reg_q2534 AND symb_decoder(16#f9#)) OR
 					(reg_q2534 AND symb_decoder(16#e2#)) OR
 					(reg_q2534 AND symb_decoder(16#01#)) OR
 					(reg_q2534 AND symb_decoder(16#f3#)) OR
 					(reg_q2534 AND symb_decoder(16#c6#)) OR
 					(reg_q2534 AND symb_decoder(16#f8#)) OR
 					(reg_q2534 AND symb_decoder(16#5b#)) OR
 					(reg_q2534 AND symb_decoder(16#4e#)) OR
 					(reg_q2534 AND symb_decoder(16#26#)) OR
 					(reg_q2534 AND symb_decoder(16#14#)) OR
 					(reg_q2534 AND symb_decoder(16#5e#)) OR
 					(reg_q2534 AND symb_decoder(16#f6#)) OR
 					(reg_q2534 AND symb_decoder(16#b4#)) OR
 					(reg_q2534 AND symb_decoder(16#c4#)) OR
 					(reg_q2534 AND symb_decoder(16#23#)) OR
 					(reg_q2534 AND symb_decoder(16#90#)) OR
 					(reg_q2534 AND symb_decoder(16#f0#)) OR
 					(reg_q2534 AND symb_decoder(16#27#)) OR
 					(reg_q2534 AND symb_decoder(16#4c#)) OR
 					(reg_q2534 AND symb_decoder(16#1a#)) OR
 					(reg_q2534 AND symb_decoder(16#70#)) OR
 					(reg_q2534 AND symb_decoder(16#10#)) OR
 					(reg_q2534 AND symb_decoder(16#59#)) OR
 					(reg_q2534 AND symb_decoder(16#61#)) OR
 					(reg_q2534 AND symb_decoder(16#b0#)) OR
 					(reg_q2534 AND symb_decoder(16#08#)) OR
 					(reg_q2534 AND symb_decoder(16#8e#)) OR
 					(reg_q2534 AND symb_decoder(16#22#)) OR
 					(reg_q2534 AND symb_decoder(16#7e#)) OR
 					(reg_q2534 AND symb_decoder(16#62#)) OR
 					(reg_q2534 AND symb_decoder(16#71#)) OR
 					(reg_q2534 AND symb_decoder(16#a8#)) OR
 					(reg_q2534 AND symb_decoder(16#a7#)) OR
 					(reg_q2534 AND symb_decoder(16#24#)) OR
 					(reg_q2534 AND symb_decoder(16#2e#)) OR
 					(reg_q2534 AND symb_decoder(16#bf#)) OR
 					(reg_q2534 AND symb_decoder(16#6e#)) OR
 					(reg_q2534 AND symb_decoder(16#1b#)) OR
 					(reg_q2534 AND symb_decoder(16#84#)) OR
 					(reg_q2534 AND symb_decoder(16#9f#)) OR
 					(reg_q2534 AND symb_decoder(16#af#)) OR
 					(reg_q2534 AND symb_decoder(16#b6#)) OR
 					(reg_q2534 AND symb_decoder(16#5d#)) OR
 					(reg_q2534 AND symb_decoder(16#1e#)) OR
 					(reg_q2534 AND symb_decoder(16#28#)) OR
 					(reg_q2534 AND symb_decoder(16#e7#)) OR
 					(reg_q2534 AND symb_decoder(16#88#)) OR
 					(reg_q2534 AND symb_decoder(16#6a#)) OR
 					(reg_q2534 AND symb_decoder(16#fa#)) OR
 					(reg_q2534 AND symb_decoder(16#45#)) OR
 					(reg_q2534 AND symb_decoder(16#6b#)) OR
 					(reg_q2534 AND symb_decoder(16#e8#)) OR
 					(reg_q2534 AND symb_decoder(16#49#)) OR
 					(reg_q2534 AND symb_decoder(16#4b#)) OR
 					(reg_q2534 AND symb_decoder(16#e1#)) OR
 					(reg_q2534 AND symb_decoder(16#51#)) OR
 					(reg_q2534 AND symb_decoder(16#b3#)) OR
 					(reg_q2534 AND symb_decoder(16#19#)) OR
 					(reg_q2534 AND symb_decoder(16#32#)) OR
 					(reg_q2534 AND symb_decoder(16#b7#)) OR
 					(reg_q2534 AND symb_decoder(16#2a#)) OR
 					(reg_q2534 AND symb_decoder(16#b1#)) OR
 					(reg_q2534 AND symb_decoder(16#d1#)) OR
 					(reg_q2534 AND symb_decoder(16#c2#)) OR
 					(reg_q2534 AND symb_decoder(16#c9#)) OR
 					(reg_q2534 AND symb_decoder(16#cb#)) OR
 					(reg_q2534 AND symb_decoder(16#63#)) OR
 					(reg_q2534 AND symb_decoder(16#cc#)) OR
 					(reg_q2534 AND symb_decoder(16#8f#)) OR
 					(reg_q2534 AND symb_decoder(16#ed#)) OR
 					(reg_q2534 AND symb_decoder(16#ec#)) OR
 					(reg_q2534 AND symb_decoder(16#36#)) OR
 					(reg_q2534 AND symb_decoder(16#85#)) OR
 					(reg_q2534 AND symb_decoder(16#c3#)) OR
 					(reg_q2534 AND symb_decoder(16#99#)) OR
 					(reg_q2534 AND symb_decoder(16#40#)) OR
 					(reg_q2534 AND symb_decoder(16#c5#)) OR
 					(reg_q2534 AND symb_decoder(16#7b#)) OR
 					(reg_q2534 AND symb_decoder(16#d2#)) OR
 					(reg_q2534 AND symb_decoder(16#e9#)) OR
 					(reg_q2534 AND symb_decoder(16#18#)) OR
 					(reg_q2534 AND symb_decoder(16#9d#)) OR
 					(reg_q2534 AND symb_decoder(16#29#)) OR
 					(reg_q2534 AND symb_decoder(16#47#)) OR
 					(reg_q2534 AND symb_decoder(16#b8#)) OR
 					(reg_q2534 AND symb_decoder(16#5f#)) OR
 					(reg_q2534 AND symb_decoder(16#92#)) OR
 					(reg_q2534 AND symb_decoder(16#ab#)) OR
 					(reg_q2534 AND symb_decoder(16#75#)) OR
 					(reg_q2534 AND symb_decoder(16#50#)) OR
 					(reg_q2534 AND symb_decoder(16#72#)) OR
 					(reg_q2534 AND symb_decoder(16#34#)) OR
 					(reg_q2534 AND symb_decoder(16#60#)) OR
 					(reg_q2534 AND symb_decoder(16#57#)) OR
 					(reg_q2534 AND symb_decoder(16#cf#)) OR
 					(reg_q2534 AND symb_decoder(16#82#)) OR
 					(reg_q2534 AND symb_decoder(16#06#)) OR
 					(reg_q2534 AND symb_decoder(16#0f#)) OR
 					(reg_q2534 AND symb_decoder(16#7a#)) OR
 					(reg_q2534 AND symb_decoder(16#bd#)) OR
 					(reg_q2534 AND symb_decoder(16#db#)) OR
 					(reg_q2534 AND symb_decoder(16#c1#)) OR
 					(reg_q2534 AND symb_decoder(16#df#)) OR
 					(reg_q2534 AND symb_decoder(16#41#)) OR
 					(reg_q2534 AND symb_decoder(16#c0#)) OR
 					(reg_q2534 AND symb_decoder(16#4d#)) OR
 					(reg_q2534 AND symb_decoder(16#0c#)) OR
 					(reg_q2534 AND symb_decoder(16#d5#)) OR
 					(reg_q2534 AND symb_decoder(16#a2#)) OR
 					(reg_q2534 AND symb_decoder(16#03#)) OR
 					(reg_q2534 AND symb_decoder(16#78#)) OR
 					(reg_q2534 AND symb_decoder(16#f5#)) OR
 					(reg_q2534 AND symb_decoder(16#76#)) OR
 					(reg_q2534 AND symb_decoder(16#42#)) OR
 					(reg_q2534 AND symb_decoder(16#6c#)) OR
 					(reg_q2534 AND symb_decoder(16#0a#)) OR
 					(reg_q2534 AND symb_decoder(16#31#)) OR
 					(reg_q2534 AND symb_decoder(16#25#)) OR
 					(reg_q2534 AND symb_decoder(16#04#)) OR
 					(reg_q2534 AND symb_decoder(16#43#)) OR
 					(reg_q2534 AND symb_decoder(16#1c#)) OR
 					(reg_q2534 AND symb_decoder(16#4a#)) OR
 					(reg_q2534 AND symb_decoder(16#55#)) OR
 					(reg_q2534 AND symb_decoder(16#a0#)) OR
 					(reg_q2534 AND symb_decoder(16#86#)) OR
 					(reg_q2534 AND symb_decoder(16#38#)) OR
 					(reg_q2534 AND symb_decoder(16#ee#)) OR
 					(reg_q2534 AND symb_decoder(16#5a#)) OR
 					(reg_q2534 AND symb_decoder(16#4f#)) OR
 					(reg_q2534 AND symb_decoder(16#3f#)) OR
 					(reg_q2534 AND symb_decoder(16#67#)) OR
 					(reg_q2534 AND symb_decoder(16#8d#)) OR
 					(reg_q2534 AND symb_decoder(16#91#)) OR
 					(reg_q2534 AND symb_decoder(16#dd#)) OR
 					(reg_q2534 AND symb_decoder(16#d3#)) OR
 					(reg_q2534 AND symb_decoder(16#d7#)) OR
 					(reg_q2534 AND symb_decoder(16#be#)) OR
 					(reg_q2534 AND symb_decoder(16#1f#)) OR
 					(reg_q2534 AND symb_decoder(16#69#)) OR
 					(reg_q2534 AND symb_decoder(16#dc#)) OR
 					(reg_q2534 AND symb_decoder(16#f4#)) OR
 					(reg_q2534 AND symb_decoder(16#ba#)) OR
 					(reg_q2534 AND symb_decoder(16#e5#)) OR
 					(reg_q2534 AND symb_decoder(16#66#)) OR
 					(reg_q2534 AND symb_decoder(16#89#)) OR
 					(reg_q2534 AND symb_decoder(16#9e#)) OR
 					(reg_q2534 AND symb_decoder(16#8c#)) OR
 					(reg_q2534 AND symb_decoder(16#b2#)) OR
 					(reg_q2534 AND symb_decoder(16#ce#)) OR
 					(reg_q2534 AND symb_decoder(16#77#)) OR
 					(reg_q2534 AND symb_decoder(16#d9#)) OR
 					(reg_q2534 AND symb_decoder(16#e6#)) OR
 					(reg_q2534 AND symb_decoder(16#80#)) OR
 					(reg_q2534 AND symb_decoder(16#e0#)) OR
 					(reg_q2534 AND symb_decoder(16#ea#)) OR
 					(reg_q2534 AND symb_decoder(16#a5#)) OR
 					(reg_q2534 AND symb_decoder(16#6f#)) OR
 					(reg_q2534 AND symb_decoder(16#98#)) OR
 					(reg_q2534 AND symb_decoder(16#12#)) OR
 					(reg_q2534 AND symb_decoder(16#2b#)) OR
 					(reg_q2534 AND symb_decoder(16#02#)) OR
 					(reg_q2534 AND symb_decoder(16#64#)) OR
 					(reg_q2534 AND symb_decoder(16#a3#)) OR
 					(reg_q2534 AND symb_decoder(16#35#)) OR
 					(reg_q2534 AND symb_decoder(16#e4#)) OR
 					(reg_q2534 AND symb_decoder(16#3c#)) OR
 					(reg_q2534 AND symb_decoder(16#a9#)) OR
 					(reg_q2534 AND symb_decoder(16#52#)) OR
 					(reg_q2534 AND symb_decoder(16#05#)) OR
 					(reg_q2534 AND symb_decoder(16#16#)) OR
 					(reg_q2534 AND symb_decoder(16#a4#)) OR
 					(reg_q2534 AND symb_decoder(16#68#)) OR
 					(reg_q2534 AND symb_decoder(16#3e#)) OR
 					(reg_q2534 AND symb_decoder(16#87#)) OR
 					(reg_q2534 AND symb_decoder(16#81#)) OR
 					(reg_q2534 AND symb_decoder(16#2d#)) OR
 					(reg_q2534 AND symb_decoder(16#1d#)) OR
 					(reg_q2534 AND symb_decoder(16#e3#)) OR
 					(reg_q2534 AND symb_decoder(16#fe#)) OR
 					(reg_q2534 AND symb_decoder(16#73#)) OR
 					(reg_q2552 AND symb_decoder(16#c5#)) OR
 					(reg_q2552 AND symb_decoder(16#40#)) OR
 					(reg_q2552 AND symb_decoder(16#93#)) OR
 					(reg_q2552 AND symb_decoder(16#ff#)) OR
 					(reg_q2552 AND symb_decoder(16#f7#)) OR
 					(reg_q2552 AND symb_decoder(16#d1#)) OR
 					(reg_q2552 AND symb_decoder(16#2e#)) OR
 					(reg_q2552 AND symb_decoder(16#9d#)) OR
 					(reg_q2552 AND symb_decoder(16#9b#)) OR
 					(reg_q2552 AND symb_decoder(16#68#)) OR
 					(reg_q2552 AND symb_decoder(16#aa#)) OR
 					(reg_q2552 AND symb_decoder(16#73#)) OR
 					(reg_q2552 AND symb_decoder(16#a0#)) OR
 					(reg_q2552 AND symb_decoder(16#7a#)) OR
 					(reg_q2552 AND symb_decoder(16#2b#)) OR
 					(reg_q2552 AND symb_decoder(16#30#)) OR
 					(reg_q2552 AND symb_decoder(16#6b#)) OR
 					(reg_q2552 AND symb_decoder(16#80#)) OR
 					(reg_q2552 AND symb_decoder(16#6d#)) OR
 					(reg_q2552 AND symb_decoder(16#2d#)) OR
 					(reg_q2552 AND symb_decoder(16#69#)) OR
 					(reg_q2552 AND symb_decoder(16#f2#)) OR
 					(reg_q2552 AND symb_decoder(16#bb#)) OR
 					(reg_q2552 AND symb_decoder(16#c0#)) OR
 					(reg_q2552 AND symb_decoder(16#ab#)) OR
 					(reg_q2552 AND symb_decoder(16#b7#)) OR
 					(reg_q2552 AND symb_decoder(16#7f#)) OR
 					(reg_q2552 AND symb_decoder(16#a6#)) OR
 					(reg_q2552 AND symb_decoder(16#6c#)) OR
 					(reg_q2552 AND symb_decoder(16#88#)) OR
 					(reg_q2552 AND symb_decoder(16#98#)) OR
 					(reg_q2552 AND symb_decoder(16#5c#)) OR
 					(reg_q2552 AND symb_decoder(16#5e#)) OR
 					(reg_q2552 AND symb_decoder(16#dc#)) OR
 					(reg_q2552 AND symb_decoder(16#42#)) OR
 					(reg_q2552 AND symb_decoder(16#be#)) OR
 					(reg_q2552 AND symb_decoder(16#e4#)) OR
 					(reg_q2552 AND symb_decoder(16#ef#)) OR
 					(reg_q2552 AND symb_decoder(16#3b#)) OR
 					(reg_q2552 AND symb_decoder(16#63#)) OR
 					(reg_q2552 AND symb_decoder(16#67#)) OR
 					(reg_q2552 AND symb_decoder(16#66#)) OR
 					(reg_q2552 AND symb_decoder(16#4a#)) OR
 					(reg_q2552 AND symb_decoder(16#14#)) OR
 					(reg_q2552 AND symb_decoder(16#62#)) OR
 					(reg_q2552 AND symb_decoder(16#96#)) OR
 					(reg_q2552 AND symb_decoder(16#f6#)) OR
 					(reg_q2552 AND symb_decoder(16#5f#)) OR
 					(reg_q2552 AND symb_decoder(16#bc#)) OR
 					(reg_q2552 AND symb_decoder(16#a1#)) OR
 					(reg_q2552 AND symb_decoder(16#d9#)) OR
 					(reg_q2552 AND symb_decoder(16#ac#)) OR
 					(reg_q2552 AND symb_decoder(16#bf#)) OR
 					(reg_q2552 AND symb_decoder(16#33#)) OR
 					(reg_q2552 AND symb_decoder(16#28#)) OR
 					(reg_q2552 AND symb_decoder(16#4e#)) OR
 					(reg_q2552 AND symb_decoder(16#7c#)) OR
 					(reg_q2552 AND symb_decoder(16#fe#)) OR
 					(reg_q2552 AND symb_decoder(16#cd#)) OR
 					(reg_q2552 AND symb_decoder(16#08#)) OR
 					(reg_q2552 AND symb_decoder(16#41#)) OR
 					(reg_q2552 AND symb_decoder(16#1e#)) OR
 					(reg_q2552 AND symb_decoder(16#8e#)) OR
 					(reg_q2552 AND symb_decoder(16#10#)) OR
 					(reg_q2552 AND symb_decoder(16#16#)) OR
 					(reg_q2552 AND symb_decoder(16#cf#)) OR
 					(reg_q2552 AND symb_decoder(16#0f#)) OR
 					(reg_q2552 AND symb_decoder(16#0d#)) OR
 					(reg_q2552 AND symb_decoder(16#83#)) OR
 					(reg_q2552 AND symb_decoder(16#64#)) OR
 					(reg_q2552 AND symb_decoder(16#1f#)) OR
 					(reg_q2552 AND symb_decoder(16#48#)) OR
 					(reg_q2552 AND symb_decoder(16#50#)) OR
 					(reg_q2552 AND symb_decoder(16#db#)) OR
 					(reg_q2552 AND symb_decoder(16#8d#)) OR
 					(reg_q2552 AND symb_decoder(16#65#)) OR
 					(reg_q2552 AND symb_decoder(16#43#)) OR
 					(reg_q2552 AND symb_decoder(16#22#)) OR
 					(reg_q2552 AND symb_decoder(16#0e#)) OR
 					(reg_q2552 AND symb_decoder(16#24#)) OR
 					(reg_q2552 AND symb_decoder(16#e2#)) OR
 					(reg_q2552 AND symb_decoder(16#6a#)) OR
 					(reg_q2552 AND symb_decoder(16#32#)) OR
 					(reg_q2552 AND symb_decoder(16#9e#)) OR
 					(reg_q2552 AND symb_decoder(16#d8#)) OR
 					(reg_q2552 AND symb_decoder(16#c3#)) OR
 					(reg_q2552 AND symb_decoder(16#ca#)) OR
 					(reg_q2552 AND symb_decoder(16#9a#)) OR
 					(reg_q2552 AND symb_decoder(16#d4#)) OR
 					(reg_q2552 AND symb_decoder(16#76#)) OR
 					(reg_q2552 AND symb_decoder(16#97#)) OR
 					(reg_q2552 AND symb_decoder(16#46#)) OR
 					(reg_q2552 AND symb_decoder(16#e1#)) OR
 					(reg_q2552 AND symb_decoder(16#75#)) OR
 					(reg_q2552 AND symb_decoder(16#c7#)) OR
 					(reg_q2552 AND symb_decoder(16#f4#)) OR
 					(reg_q2552 AND symb_decoder(16#57#)) OR
 					(reg_q2552 AND symb_decoder(16#85#)) OR
 					(reg_q2552 AND symb_decoder(16#47#)) OR
 					(reg_q2552 AND symb_decoder(16#d2#)) OR
 					(reg_q2552 AND symb_decoder(16#49#)) OR
 					(reg_q2552 AND symb_decoder(16#90#)) OR
 					(reg_q2552 AND symb_decoder(16#af#)) OR
 					(reg_q2552 AND symb_decoder(16#00#)) OR
 					(reg_q2552 AND symb_decoder(16#56#)) OR
 					(reg_q2552 AND symb_decoder(16#70#)) OR
 					(reg_q2552 AND symb_decoder(16#89#)) OR
 					(reg_q2552 AND symb_decoder(16#4f#)) OR
 					(reg_q2552 AND symb_decoder(16#d0#)) OR
 					(reg_q2552 AND symb_decoder(16#d5#)) OR
 					(reg_q2552 AND symb_decoder(16#c8#)) OR
 					(reg_q2552 AND symb_decoder(16#94#)) OR
 					(reg_q2552 AND symb_decoder(16#e0#)) OR
 					(reg_q2552 AND symb_decoder(16#92#)) OR
 					(reg_q2552 AND symb_decoder(16#ee#)) OR
 					(reg_q2552 AND symb_decoder(16#87#)) OR
 					(reg_q2552 AND symb_decoder(16#b2#)) OR
 					(reg_q2552 AND symb_decoder(16#ec#)) OR
 					(reg_q2552 AND symb_decoder(16#4c#)) OR
 					(reg_q2552 AND symb_decoder(16#e9#)) OR
 					(reg_q2552 AND symb_decoder(16#7d#)) OR
 					(reg_q2552 AND symb_decoder(16#c9#)) OR
 					(reg_q2552 AND symb_decoder(16#d6#)) OR
 					(reg_q2552 AND symb_decoder(16#f9#)) OR
 					(reg_q2552 AND symb_decoder(16#72#)) OR
 					(reg_q2552 AND symb_decoder(16#26#)) OR
 					(reg_q2552 AND symb_decoder(16#d3#)) OR
 					(reg_q2552 AND symb_decoder(16#20#)) OR
 					(reg_q2552 AND symb_decoder(16#b1#)) OR
 					(reg_q2552 AND symb_decoder(16#51#)) OR
 					(reg_q2552 AND symb_decoder(16#95#)) OR
 					(reg_q2552 AND symb_decoder(16#b0#)) OR
 					(reg_q2552 AND symb_decoder(16#35#)) OR
 					(reg_q2552 AND symb_decoder(16#1a#)) OR
 					(reg_q2552 AND symb_decoder(16#06#)) OR
 					(reg_q2552 AND symb_decoder(16#54#)) OR
 					(reg_q2552 AND symb_decoder(16#ae#)) OR
 					(reg_q2552 AND symb_decoder(16#c4#)) OR
 					(reg_q2552 AND symb_decoder(16#3e#)) OR
 					(reg_q2552 AND symb_decoder(16#0a#)) OR
 					(reg_q2552 AND symb_decoder(16#a9#)) OR
 					(reg_q2552 AND symb_decoder(16#da#)) OR
 					(reg_q2552 AND symb_decoder(16#a3#)) OR
 					(reg_q2552 AND symb_decoder(16#86#)) OR
 					(reg_q2552 AND symb_decoder(16#07#)) OR
 					(reg_q2552 AND symb_decoder(16#a7#)) OR
 					(reg_q2552 AND symb_decoder(16#7e#)) OR
 					(reg_q2552 AND symb_decoder(16#15#)) OR
 					(reg_q2552 AND symb_decoder(16#b4#)) OR
 					(reg_q2552 AND symb_decoder(16#5b#)) OR
 					(reg_q2552 AND symb_decoder(16#55#)) OR
 					(reg_q2552 AND symb_decoder(16#02#)) OR
 					(reg_q2552 AND symb_decoder(16#3d#)) OR
 					(reg_q2552 AND symb_decoder(16#fd#)) OR
 					(reg_q2552 AND symb_decoder(16#c2#)) OR
 					(reg_q2552 AND symb_decoder(16#74#)) OR
 					(reg_q2552 AND symb_decoder(16#ce#)) OR
 					(reg_q2552 AND symb_decoder(16#fa#)) OR
 					(reg_q2552 AND symb_decoder(16#91#)) OR
 					(reg_q2552 AND symb_decoder(16#a8#)) OR
 					(reg_q2552 AND symb_decoder(16#12#)) OR
 					(reg_q2552 AND symb_decoder(16#78#)) OR
 					(reg_q2552 AND symb_decoder(16#18#)) OR
 					(reg_q2552 AND symb_decoder(16#01#)) OR
 					(reg_q2552 AND symb_decoder(16#f1#)) OR
 					(reg_q2552 AND symb_decoder(16#e3#)) OR
 					(reg_q2552 AND symb_decoder(16#7b#)) OR
 					(reg_q2552 AND symb_decoder(16#eb#)) OR
 					(reg_q2552 AND symb_decoder(16#f3#)) OR
 					(reg_q2552 AND symb_decoder(16#11#)) OR
 					(reg_q2552 AND symb_decoder(16#19#)) OR
 					(reg_q2552 AND symb_decoder(16#25#)) OR
 					(reg_q2552 AND symb_decoder(16#b9#)) OR
 					(reg_q2552 AND symb_decoder(16#cc#)) OR
 					(reg_q2552 AND symb_decoder(16#8a#)) OR
 					(reg_q2552 AND symb_decoder(16#38#)) OR
 					(reg_q2552 AND symb_decoder(16#71#)) OR
 					(reg_q2552 AND symb_decoder(16#52#)) OR
 					(reg_q2552 AND symb_decoder(16#58#)) OR
 					(reg_q2552 AND symb_decoder(16#df#)) OR
 					(reg_q2552 AND symb_decoder(16#ad#)) OR
 					(reg_q2552 AND symb_decoder(16#fc#)) OR
 					(reg_q2552 AND symb_decoder(16#f0#)) OR
 					(reg_q2552 AND symb_decoder(16#dd#)) OR
 					(reg_q2552 AND symb_decoder(16#79#)) OR
 					(reg_q2552 AND symb_decoder(16#45#)) OR
 					(reg_q2552 AND symb_decoder(16#a2#)) OR
 					(reg_q2552 AND symb_decoder(16#4b#)) OR
 					(reg_q2552 AND symb_decoder(16#8f#)) OR
 					(reg_q2552 AND symb_decoder(16#cb#)) OR
 					(reg_q2552 AND symb_decoder(16#bd#)) OR
 					(reg_q2552 AND symb_decoder(16#1c#)) OR
 					(reg_q2552 AND symb_decoder(16#3a#)) OR
 					(reg_q2552 AND symb_decoder(16#99#)) OR
 					(reg_q2552 AND symb_decoder(16#2c#)) OR
 					(reg_q2552 AND symb_decoder(16#ed#)) OR
 					(reg_q2552 AND symb_decoder(16#13#)) OR
 					(reg_q2552 AND symb_decoder(16#b5#)) OR
 					(reg_q2552 AND symb_decoder(16#1d#)) OR
 					(reg_q2552 AND symb_decoder(16#b6#)) OR
 					(reg_q2552 AND symb_decoder(16#77#)) OR
 					(reg_q2552 AND symb_decoder(16#39#)) OR
 					(reg_q2552 AND symb_decoder(16#5a#)) OR
 					(reg_q2552 AND symb_decoder(16#37#)) OR
 					(reg_q2552 AND symb_decoder(16#9f#)) OR
 					(reg_q2552 AND symb_decoder(16#a4#)) OR
 					(reg_q2552 AND symb_decoder(16#6e#)) OR
 					(reg_q2552 AND symb_decoder(16#84#)) OR
 					(reg_q2552 AND symb_decoder(16#1b#)) OR
 					(reg_q2552 AND symb_decoder(16#17#)) OR
 					(reg_q2552 AND symb_decoder(16#a5#)) OR
 					(reg_q2552 AND symb_decoder(16#4d#)) OR
 					(reg_q2552 AND symb_decoder(16#23#)) OR
 					(reg_q2552 AND symb_decoder(16#e6#)) OR
 					(reg_q2552 AND symb_decoder(16#b8#)) OR
 					(reg_q2552 AND symb_decoder(16#ea#)) OR
 					(reg_q2552 AND symb_decoder(16#2f#)) OR
 					(reg_q2552 AND symb_decoder(16#c1#)) OR
 					(reg_q2552 AND symb_decoder(16#0c#)) OR
 					(reg_q2552 AND symb_decoder(16#05#)) OR
 					(reg_q2552 AND symb_decoder(16#81#)) OR
 					(reg_q2552 AND symb_decoder(16#0b#)) OR
 					(reg_q2552 AND symb_decoder(16#fb#)) OR
 					(reg_q2552 AND symb_decoder(16#03#)) OR
 					(reg_q2552 AND symb_decoder(16#61#)) OR
 					(reg_q2552 AND symb_decoder(16#34#)) OR
 					(reg_q2552 AND symb_decoder(16#6f#)) OR
 					(reg_q2552 AND symb_decoder(16#04#)) OR
 					(reg_q2552 AND symb_decoder(16#44#)) OR
 					(reg_q2552 AND symb_decoder(16#3f#)) OR
 					(reg_q2552 AND symb_decoder(16#5d#)) OR
 					(reg_q2552 AND symb_decoder(16#f5#)) OR
 					(reg_q2552 AND symb_decoder(16#b3#)) OR
 					(reg_q2552 AND symb_decoder(16#d7#)) OR
 					(reg_q2552 AND symb_decoder(16#f8#)) OR
 					(reg_q2552 AND symb_decoder(16#60#)) OR
 					(reg_q2552 AND symb_decoder(16#3c#)) OR
 					(reg_q2552 AND symb_decoder(16#29#)) OR
 					(reg_q2552 AND symb_decoder(16#2a#)) OR
 					(reg_q2552 AND symb_decoder(16#09#)) OR
 					(reg_q2552 AND symb_decoder(16#e5#)) OR
 					(reg_q2552 AND symb_decoder(16#e8#)) OR
 					(reg_q2552 AND symb_decoder(16#27#)) OR
 					(reg_q2552 AND symb_decoder(16#c6#)) OR
 					(reg_q2552 AND symb_decoder(16#ba#)) OR
 					(reg_q2552 AND symb_decoder(16#53#)) OR
 					(reg_q2552 AND symb_decoder(16#59#)) OR
 					(reg_q2552 AND symb_decoder(16#9c#)) OR
 					(reg_q2552 AND symb_decoder(16#82#)) OR
 					(reg_q2552 AND symb_decoder(16#36#)) OR
 					(reg_q2552 AND symb_decoder(16#8c#)) OR
 					(reg_q2552 AND symb_decoder(16#de#)) OR
 					(reg_q2552 AND symb_decoder(16#21#)) OR
 					(reg_q2552 AND symb_decoder(16#8b#)) OR
 					(reg_q2552 AND symb_decoder(16#e7#)) OR
 					(reg_q2552 AND symb_decoder(16#31#));
reg_q2552_init <= '0' ;
	p_reg_q2552: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2552 <= reg_q2552_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2552 <= reg_q2552_init;
        else
          reg_q2552 <= reg_q2552_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1482_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1482 AND symb_decoder(16#2c#)) OR
 					(reg_q1482 AND symb_decoder(16#cf#)) OR
 					(reg_q1482 AND symb_decoder(16#92#)) OR
 					(reg_q1482 AND symb_decoder(16#d2#)) OR
 					(reg_q1482 AND symb_decoder(16#f7#)) OR
 					(reg_q1482 AND symb_decoder(16#fc#)) OR
 					(reg_q1482 AND symb_decoder(16#53#)) OR
 					(reg_q1482 AND symb_decoder(16#16#)) OR
 					(reg_q1482 AND symb_decoder(16#e2#)) OR
 					(reg_q1482 AND symb_decoder(16#cc#)) OR
 					(reg_q1482 AND symb_decoder(16#ed#)) OR
 					(reg_q1482 AND symb_decoder(16#20#)) OR
 					(reg_q1482 AND symb_decoder(16#f4#)) OR
 					(reg_q1482 AND symb_decoder(16#11#)) OR
 					(reg_q1482 AND symb_decoder(16#bc#)) OR
 					(reg_q1482 AND symb_decoder(16#31#)) OR
 					(reg_q1482 AND symb_decoder(16#97#)) OR
 					(reg_q1482 AND symb_decoder(16#28#)) OR
 					(reg_q1482 AND symb_decoder(16#e1#)) OR
 					(reg_q1482 AND symb_decoder(16#ae#)) OR
 					(reg_q1482 AND symb_decoder(16#76#)) OR
 					(reg_q1482 AND symb_decoder(16#bd#)) OR
 					(reg_q1482 AND symb_decoder(16#e6#)) OR
 					(reg_q1482 AND symb_decoder(16#e4#)) OR
 					(reg_q1482 AND symb_decoder(16#f8#)) OR
 					(reg_q1482 AND symb_decoder(16#a0#)) OR
 					(reg_q1482 AND symb_decoder(16#47#)) OR
 					(reg_q1482 AND symb_decoder(16#0d#)) OR
 					(reg_q1482 AND symb_decoder(16#a9#)) OR
 					(reg_q1482 AND symb_decoder(16#6b#)) OR
 					(reg_q1482 AND symb_decoder(16#59#)) OR
 					(reg_q1482 AND symb_decoder(16#af#)) OR
 					(reg_q1482 AND symb_decoder(16#23#)) OR
 					(reg_q1482 AND symb_decoder(16#4e#)) OR
 					(reg_q1482 AND symb_decoder(16#70#)) OR
 					(reg_q1482 AND symb_decoder(16#36#)) OR
 					(reg_q1482 AND symb_decoder(16#75#)) OR
 					(reg_q1482 AND symb_decoder(16#08#)) OR
 					(reg_q1482 AND symb_decoder(16#a8#)) OR
 					(reg_q1482 AND symb_decoder(16#f5#)) OR
 					(reg_q1482 AND symb_decoder(16#3f#)) OR
 					(reg_q1482 AND symb_decoder(16#be#)) OR
 					(reg_q1482 AND symb_decoder(16#04#)) OR
 					(reg_q1482 AND symb_decoder(16#91#)) OR
 					(reg_q1482 AND symb_decoder(16#1f#)) OR
 					(reg_q1482 AND symb_decoder(16#1c#)) OR
 					(reg_q1482 AND symb_decoder(16#7e#)) OR
 					(reg_q1482 AND symb_decoder(16#b7#)) OR
 					(reg_q1482 AND symb_decoder(16#b9#)) OR
 					(reg_q1482 AND symb_decoder(16#b5#)) OR
 					(reg_q1482 AND symb_decoder(16#4c#)) OR
 					(reg_q1482 AND symb_decoder(16#0f#)) OR
 					(reg_q1482 AND symb_decoder(16#12#)) OR
 					(reg_q1482 AND symb_decoder(16#b4#)) OR
 					(reg_q1482 AND symb_decoder(16#40#)) OR
 					(reg_q1482 AND symb_decoder(16#8d#)) OR
 					(reg_q1482 AND symb_decoder(16#c6#)) OR
 					(reg_q1482 AND symb_decoder(16#7c#)) OR
 					(reg_q1482 AND symb_decoder(16#9f#)) OR
 					(reg_q1482 AND symb_decoder(16#6d#)) OR
 					(reg_q1482 AND symb_decoder(16#4b#)) OR
 					(reg_q1482 AND symb_decoder(16#0c#)) OR
 					(reg_q1482 AND symb_decoder(16#9a#)) OR
 					(reg_q1482 AND symb_decoder(16#c3#)) OR
 					(reg_q1482 AND symb_decoder(16#63#)) OR
 					(reg_q1482 AND symb_decoder(16#ca#)) OR
 					(reg_q1482 AND symb_decoder(16#ff#)) OR
 					(reg_q1482 AND symb_decoder(16#02#)) OR
 					(reg_q1482 AND symb_decoder(16#6c#)) OR
 					(reg_q1482 AND symb_decoder(16#9c#)) OR
 					(reg_q1482 AND symb_decoder(16#ba#)) OR
 					(reg_q1482 AND symb_decoder(16#66#)) OR
 					(reg_q1482 AND symb_decoder(16#fd#)) OR
 					(reg_q1482 AND symb_decoder(16#65#)) OR
 					(reg_q1482 AND symb_decoder(16#45#)) OR
 					(reg_q1482 AND symb_decoder(16#d4#)) OR
 					(reg_q1482 AND symb_decoder(16#8f#)) OR
 					(reg_q1482 AND symb_decoder(16#a1#)) OR
 					(reg_q1482 AND symb_decoder(16#29#)) OR
 					(reg_q1482 AND symb_decoder(16#8e#)) OR
 					(reg_q1482 AND symb_decoder(16#83#)) OR
 					(reg_q1482 AND symb_decoder(16#2f#)) OR
 					(reg_q1482 AND symb_decoder(16#d1#)) OR
 					(reg_q1482 AND symb_decoder(16#c9#)) OR
 					(reg_q1482 AND symb_decoder(16#fb#)) OR
 					(reg_q1482 AND symb_decoder(16#69#)) OR
 					(reg_q1482 AND symb_decoder(16#ab#)) OR
 					(reg_q1482 AND symb_decoder(16#42#)) OR
 					(reg_q1482 AND symb_decoder(16#6e#)) OR
 					(reg_q1482 AND symb_decoder(16#2b#)) OR
 					(reg_q1482 AND symb_decoder(16#8c#)) OR
 					(reg_q1482 AND symb_decoder(16#54#)) OR
 					(reg_q1482 AND symb_decoder(16#3d#)) OR
 					(reg_q1482 AND symb_decoder(16#aa#)) OR
 					(reg_q1482 AND symb_decoder(16#44#)) OR
 					(reg_q1482 AND symb_decoder(16#62#)) OR
 					(reg_q1482 AND symb_decoder(16#c7#)) OR
 					(reg_q1482 AND symb_decoder(16#dd#)) OR
 					(reg_q1482 AND symb_decoder(16#50#)) OR
 					(reg_q1482 AND symb_decoder(16#4d#)) OR
 					(reg_q1482 AND symb_decoder(16#eb#)) OR
 					(reg_q1482 AND symb_decoder(16#0e#)) OR
 					(reg_q1482 AND symb_decoder(16#3a#)) OR
 					(reg_q1482 AND symb_decoder(16#3c#)) OR
 					(reg_q1482 AND symb_decoder(16#2d#)) OR
 					(reg_q1482 AND symb_decoder(16#b0#)) OR
 					(reg_q1482 AND symb_decoder(16#db#)) OR
 					(reg_q1482 AND symb_decoder(16#b3#)) OR
 					(reg_q1482 AND symb_decoder(16#55#)) OR
 					(reg_q1482 AND symb_decoder(16#5a#)) OR
 					(reg_q1482 AND symb_decoder(16#3e#)) OR
 					(reg_q1482 AND symb_decoder(16#05#)) OR
 					(reg_q1482 AND symb_decoder(16#d8#)) OR
 					(reg_q1482 AND symb_decoder(16#56#)) OR
 					(reg_q1482 AND symb_decoder(16#19#)) OR
 					(reg_q1482 AND symb_decoder(16#e7#)) OR
 					(reg_q1482 AND symb_decoder(16#d0#)) OR
 					(reg_q1482 AND symb_decoder(16#c0#)) OR
 					(reg_q1482 AND symb_decoder(16#a5#)) OR
 					(reg_q1482 AND symb_decoder(16#f6#)) OR
 					(reg_q1482 AND symb_decoder(16#48#)) OR
 					(reg_q1482 AND symb_decoder(16#ad#)) OR
 					(reg_q1482 AND symb_decoder(16#43#)) OR
 					(reg_q1482 AND symb_decoder(16#c5#)) OR
 					(reg_q1482 AND symb_decoder(16#cd#)) OR
 					(reg_q1482 AND symb_decoder(16#9e#)) OR
 					(reg_q1482 AND symb_decoder(16#c8#)) OR
 					(reg_q1482 AND symb_decoder(16#37#)) OR
 					(reg_q1482 AND symb_decoder(16#87#)) OR
 					(reg_q1482 AND symb_decoder(16#27#)) OR
 					(reg_q1482 AND symb_decoder(16#32#)) OR
 					(reg_q1482 AND symb_decoder(16#bb#)) OR
 					(reg_q1482 AND symb_decoder(16#b8#)) OR
 					(reg_q1482 AND symb_decoder(16#5e#)) OR
 					(reg_q1482 AND symb_decoder(16#93#)) OR
 					(reg_q1482 AND symb_decoder(16#67#)) OR
 					(reg_q1482 AND symb_decoder(16#ac#)) OR
 					(reg_q1482 AND symb_decoder(16#1b#)) OR
 					(reg_q1482 AND symb_decoder(16#60#)) OR
 					(reg_q1482 AND symb_decoder(16#78#)) OR
 					(reg_q1482 AND symb_decoder(16#98#)) OR
 					(reg_q1482 AND symb_decoder(16#15#)) OR
 					(reg_q1482 AND symb_decoder(16#e0#)) OR
 					(reg_q1482 AND symb_decoder(16#3b#)) OR
 					(reg_q1482 AND symb_decoder(16#0a#)) OR
 					(reg_q1482 AND symb_decoder(16#72#)) OR
 					(reg_q1482 AND symb_decoder(16#39#)) OR
 					(reg_q1482 AND symb_decoder(16#71#)) OR
 					(reg_q1482 AND symb_decoder(16#1a#)) OR
 					(reg_q1482 AND symb_decoder(16#5b#)) OR
 					(reg_q1482 AND symb_decoder(16#35#)) OR
 					(reg_q1482 AND symb_decoder(16#8b#)) OR
 					(reg_q1482 AND symb_decoder(16#fa#)) OR
 					(reg_q1482 AND symb_decoder(16#77#)) OR
 					(reg_q1482 AND symb_decoder(16#0b#)) OR
 					(reg_q1482 AND symb_decoder(16#96#)) OR
 					(reg_q1482 AND symb_decoder(16#ce#)) OR
 					(reg_q1482 AND symb_decoder(16#d6#)) OR
 					(reg_q1482 AND symb_decoder(16#f0#)) OR
 					(reg_q1482 AND symb_decoder(16#01#)) OR
 					(reg_q1482 AND symb_decoder(16#b1#)) OR
 					(reg_q1482 AND symb_decoder(16#d5#)) OR
 					(reg_q1482 AND symb_decoder(16#6a#)) OR
 					(reg_q1482 AND symb_decoder(16#09#)) OR
 					(reg_q1482 AND symb_decoder(16#c2#)) OR
 					(reg_q1482 AND symb_decoder(16#84#)) OR
 					(reg_q1482 AND symb_decoder(16#7b#)) OR
 					(reg_q1482 AND symb_decoder(16#c1#)) OR
 					(reg_q1482 AND symb_decoder(16#5c#)) OR
 					(reg_q1482 AND symb_decoder(16#f1#)) OR
 					(reg_q1482 AND symb_decoder(16#2e#)) OR
 					(reg_q1482 AND symb_decoder(16#86#)) OR
 					(reg_q1482 AND symb_decoder(16#2a#)) OR
 					(reg_q1482 AND symb_decoder(16#a4#)) OR
 					(reg_q1482 AND symb_decoder(16#57#)) OR
 					(reg_q1482 AND symb_decoder(16#52#)) OR
 					(reg_q1482 AND symb_decoder(16#a3#)) OR
 					(reg_q1482 AND symb_decoder(16#cb#)) OR
 					(reg_q1482 AND symb_decoder(16#9b#)) OR
 					(reg_q1482 AND symb_decoder(16#bf#)) OR
 					(reg_q1482 AND symb_decoder(16#79#)) OR
 					(reg_q1482 AND symb_decoder(16#d3#)) OR
 					(reg_q1482 AND symb_decoder(16#99#)) OR
 					(reg_q1482 AND symb_decoder(16#85#)) OR
 					(reg_q1482 AND symb_decoder(16#7f#)) OR
 					(reg_q1482 AND symb_decoder(16#a7#)) OR
 					(reg_q1482 AND symb_decoder(16#34#)) OR
 					(reg_q1482 AND symb_decoder(16#5d#)) OR
 					(reg_q1482 AND symb_decoder(16#fe#)) OR
 					(reg_q1482 AND symb_decoder(16#17#)) OR
 					(reg_q1482 AND symb_decoder(16#95#)) OR
 					(reg_q1482 AND symb_decoder(16#7a#)) OR
 					(reg_q1482 AND symb_decoder(16#90#)) OR
 					(reg_q1482 AND symb_decoder(16#68#)) OR
 					(reg_q1482 AND symb_decoder(16#dc#)) OR
 					(reg_q1482 AND symb_decoder(16#81#)) OR
 					(reg_q1482 AND symb_decoder(16#9d#)) OR
 					(reg_q1482 AND symb_decoder(16#00#)) OR
 					(reg_q1482 AND symb_decoder(16#41#)) OR
 					(reg_q1482 AND symb_decoder(16#e5#)) OR
 					(reg_q1482 AND symb_decoder(16#58#)) OR
 					(reg_q1482 AND symb_decoder(16#14#)) OR
 					(reg_q1482 AND symb_decoder(16#ee#)) OR
 					(reg_q1482 AND symb_decoder(16#26#)) OR
 					(reg_q1482 AND symb_decoder(16#30#)) OR
 					(reg_q1482 AND symb_decoder(16#ec#)) OR
 					(reg_q1482 AND symb_decoder(16#ea#)) OR
 					(reg_q1482 AND symb_decoder(16#f3#)) OR
 					(reg_q1482 AND symb_decoder(16#07#)) OR
 					(reg_q1482 AND symb_decoder(16#94#)) OR
 					(reg_q1482 AND symb_decoder(16#4f#)) OR
 					(reg_q1482 AND symb_decoder(16#a2#)) OR
 					(reg_q1482 AND symb_decoder(16#f2#)) OR
 					(reg_q1482 AND symb_decoder(16#e3#)) OR
 					(reg_q1482 AND symb_decoder(16#24#)) OR
 					(reg_q1482 AND symb_decoder(16#18#)) OR
 					(reg_q1482 AND symb_decoder(16#06#)) OR
 					(reg_q1482 AND symb_decoder(16#da#)) OR
 					(reg_q1482 AND symb_decoder(16#73#)) OR
 					(reg_q1482 AND symb_decoder(16#49#)) OR
 					(reg_q1482 AND symb_decoder(16#f9#)) OR
 					(reg_q1482 AND symb_decoder(16#38#)) OR
 					(reg_q1482 AND symb_decoder(16#de#)) OR
 					(reg_q1482 AND symb_decoder(16#c4#)) OR
 					(reg_q1482 AND symb_decoder(16#10#)) OR
 					(reg_q1482 AND symb_decoder(16#89#)) OR
 					(reg_q1482 AND symb_decoder(16#1e#)) OR
 					(reg_q1482 AND symb_decoder(16#1d#)) OR
 					(reg_q1482 AND symb_decoder(16#e9#)) OR
 					(reg_q1482 AND symb_decoder(16#d7#)) OR
 					(reg_q1482 AND symb_decoder(16#d9#)) OR
 					(reg_q1482 AND symb_decoder(16#03#)) OR
 					(reg_q1482 AND symb_decoder(16#64#)) OR
 					(reg_q1482 AND symb_decoder(16#ef#)) OR
 					(reg_q1482 AND symb_decoder(16#22#)) OR
 					(reg_q1482 AND symb_decoder(16#8a#)) OR
 					(reg_q1482 AND symb_decoder(16#88#)) OR
 					(reg_q1482 AND symb_decoder(16#82#)) OR
 					(reg_q1482 AND symb_decoder(16#e8#)) OR
 					(reg_q1482 AND symb_decoder(16#b2#)) OR
 					(reg_q1482 AND symb_decoder(16#61#)) OR
 					(reg_q1482 AND symb_decoder(16#5f#)) OR
 					(reg_q1482 AND symb_decoder(16#25#)) OR
 					(reg_q1482 AND symb_decoder(16#46#)) OR
 					(reg_q1482 AND symb_decoder(16#33#)) OR
 					(reg_q1482 AND symb_decoder(16#a6#)) OR
 					(reg_q1482 AND symb_decoder(16#74#)) OR
 					(reg_q1482 AND symb_decoder(16#7d#)) OR
 					(reg_q1482 AND symb_decoder(16#4a#)) OR
 					(reg_q1482 AND symb_decoder(16#df#)) OR
 					(reg_q1482 AND symb_decoder(16#80#)) OR
 					(reg_q1482 AND symb_decoder(16#13#)) OR
 					(reg_q1482 AND symb_decoder(16#6f#)) OR
 					(reg_q1482 AND symb_decoder(16#21#)) OR
 					(reg_q1482 AND symb_decoder(16#51#)) OR
 					(reg_q1482 AND symb_decoder(16#b6#));
reg_q1482_init <= '0' ;
	p_reg_q1482: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1482 <= reg_q1482_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1482 <= reg_q1482_init;
        else
          reg_q1482 <= reg_q1482_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph55

reg_q2080_in <= (reg_q2078 AND symb_decoder(16#2f#));
reg_q606_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q604 AND symb_decoder(16#73#)) OR
 					(reg_q604 AND symb_decoder(16#53#));
reg_q342_in <= (reg_q342 AND symb_decoder(16#33#)) OR
 					(reg_q342 AND symb_decoder(16#30#)) OR
 					(reg_q342 AND symb_decoder(16#37#)) OR
 					(reg_q342 AND symb_decoder(16#34#)) OR
 					(reg_q342 AND symb_decoder(16#39#)) OR
 					(reg_q342 AND symb_decoder(16#35#)) OR
 					(reg_q342 AND symb_decoder(16#36#)) OR
 					(reg_q342 AND symb_decoder(16#38#)) OR
 					(reg_q342 AND symb_decoder(16#31#)) OR
 					(reg_q342 AND symb_decoder(16#32#)) OR
 					(reg_q340 AND symb_decoder(16#34#)) OR
 					(reg_q340 AND symb_decoder(16#36#)) OR
 					(reg_q340 AND symb_decoder(16#38#)) OR
 					(reg_q340 AND symb_decoder(16#37#)) OR
 					(reg_q340 AND symb_decoder(16#31#)) OR
 					(reg_q340 AND symb_decoder(16#35#)) OR
 					(reg_q340 AND symb_decoder(16#39#)) OR
 					(reg_q340 AND symb_decoder(16#30#)) OR
 					(reg_q340 AND symb_decoder(16#32#)) OR
 					(reg_q340 AND symb_decoder(16#33#));
reg_q2435_in <= (reg_q2433 AND symb_decoder(16#2f#));
reg_q2641_in <= (reg_q2641 AND symb_decoder(16#31#)) OR
 					(reg_q2641 AND symb_decoder(16#33#)) OR
 					(reg_q2641 AND symb_decoder(16#37#)) OR
 					(reg_q2641 AND symb_decoder(16#36#)) OR
 					(reg_q2641 AND symb_decoder(16#35#)) OR
 					(reg_q2641 AND symb_decoder(16#30#)) OR
 					(reg_q2641 AND symb_decoder(16#32#)) OR
 					(reg_q2641 AND symb_decoder(16#39#)) OR
 					(reg_q2641 AND symb_decoder(16#38#)) OR
 					(reg_q2641 AND symb_decoder(16#34#)) OR
 					(reg_q2639 AND symb_decoder(16#39#)) OR
 					(reg_q2639 AND symb_decoder(16#34#)) OR
 					(reg_q2639 AND symb_decoder(16#38#)) OR
 					(reg_q2639 AND symb_decoder(16#36#)) OR
 					(reg_q2639 AND symb_decoder(16#32#)) OR
 					(reg_q2639 AND symb_decoder(16#31#)) OR
 					(reg_q2639 AND symb_decoder(16#37#)) OR
 					(reg_q2639 AND symb_decoder(16#33#)) OR
 					(reg_q2639 AND symb_decoder(16#30#)) OR
 					(reg_q2639 AND symb_decoder(16#35#));
reg_q435_in <= (reg_q433 AND symb_decoder(16#57#)) OR
 					(reg_q433 AND symb_decoder(16#77#));
reg_q2116_in <= (reg_q2218 AND symb_decoder(16#6e#)) OR
 					(reg_q2218 AND symb_decoder(16#4e#)) OR
 					(reg_q2112 AND symb_decoder(16#6e#)) OR
 					(reg_q2112 AND symb_decoder(16#4e#));
reg_q1465_in <= (reg_q1465 AND symb_decoder(16#0c#)) OR
 					(reg_q1465 AND symb_decoder(16#20#)) OR
 					(reg_q1465 AND symb_decoder(16#09#)) OR
 					(reg_q1465 AND symb_decoder(16#0a#)) OR
 					(reg_q1465 AND symb_decoder(16#0d#)) OR
 					(reg_q1463 AND symb_decoder(16#20#)) OR
 					(reg_q1463 AND symb_decoder(16#09#)) OR
 					(reg_q1463 AND symb_decoder(16#0a#)) OR
 					(reg_q1463 AND symb_decoder(16#0c#)) OR
 					(reg_q1463 AND symb_decoder(16#0d#));
reg_q2643_in <= (reg_q2641 AND symb_decoder(16#2e#));
reg_q296_in <= (reg_q294 AND symb_decoder(16#49#)) OR
 					(reg_q294 AND symb_decoder(16#69#));
reg_q2241_in <= (reg_q2241 AND symb_decoder(16#37#)) OR
 					(reg_q2241 AND symb_decoder(16#32#)) OR
 					(reg_q2241 AND symb_decoder(16#35#)) OR
 					(reg_q2241 AND symb_decoder(16#33#)) OR
 					(reg_q2241 AND symb_decoder(16#34#)) OR
 					(reg_q2241 AND symb_decoder(16#31#)) OR
 					(reg_q2241 AND symb_decoder(16#38#)) OR
 					(reg_q2241 AND symb_decoder(16#39#)) OR
 					(reg_q2241 AND symb_decoder(16#36#)) OR
 					(reg_q2241 AND symb_decoder(16#30#)) OR
 					(reg_q2239 AND symb_decoder(16#37#)) OR
 					(reg_q2239 AND symb_decoder(16#31#)) OR
 					(reg_q2239 AND symb_decoder(16#36#)) OR
 					(reg_q2239 AND symb_decoder(16#34#)) OR
 					(reg_q2239 AND symb_decoder(16#32#)) OR
 					(reg_q2239 AND symb_decoder(16#39#)) OR
 					(reg_q2239 AND symb_decoder(16#33#)) OR
 					(reg_q2239 AND symb_decoder(16#35#)) OR
 					(reg_q2239 AND symb_decoder(16#38#)) OR
 					(reg_q2239 AND symb_decoder(16#30#));
reg_q2237_in <= (reg_q2235 AND symb_decoder(16#38#)) OR
 					(reg_q2235 AND symb_decoder(16#39#)) OR
 					(reg_q2235 AND symb_decoder(16#37#)) OR
 					(reg_q2235 AND symb_decoder(16#31#)) OR
 					(reg_q2235 AND symb_decoder(16#34#)) OR
 					(reg_q2235 AND symb_decoder(16#36#)) OR
 					(reg_q2235 AND symb_decoder(16#35#)) OR
 					(reg_q2235 AND symb_decoder(16#33#)) OR
 					(reg_q2235 AND symb_decoder(16#30#)) OR
 					(reg_q2235 AND symb_decoder(16#32#)) OR
 					(reg_q2237 AND symb_decoder(16#35#)) OR
 					(reg_q2237 AND symb_decoder(16#34#)) OR
 					(reg_q2237 AND symb_decoder(16#39#)) OR
 					(reg_q2237 AND symb_decoder(16#36#)) OR
 					(reg_q2237 AND symb_decoder(16#33#)) OR
 					(reg_q2237 AND symb_decoder(16#38#)) OR
 					(reg_q2237 AND symb_decoder(16#32#)) OR
 					(reg_q2237 AND symb_decoder(16#37#)) OR
 					(reg_q2237 AND symb_decoder(16#30#)) OR
 					(reg_q2237 AND symb_decoder(16#31#));
reg_q2647_in <= (reg_q2645 AND symb_decoder(16#2e#));
reg_q2649_in <= (reg_q2647 AND symb_decoder(16#32#)) OR
 					(reg_q2647 AND symb_decoder(16#37#)) OR
 					(reg_q2647 AND symb_decoder(16#39#)) OR
 					(reg_q2647 AND symb_decoder(16#33#)) OR
 					(reg_q2647 AND symb_decoder(16#36#)) OR
 					(reg_q2647 AND symb_decoder(16#35#)) OR
 					(reg_q2647 AND symb_decoder(16#30#)) OR
 					(reg_q2647 AND symb_decoder(16#34#)) OR
 					(reg_q2647 AND symb_decoder(16#31#)) OR
 					(reg_q2647 AND symb_decoder(16#38#)) OR
 					(reg_q2649 AND symb_decoder(16#35#)) OR
 					(reg_q2649 AND symb_decoder(16#30#)) OR
 					(reg_q2649 AND symb_decoder(16#39#)) OR
 					(reg_q2649 AND symb_decoder(16#36#)) OR
 					(reg_q2649 AND symb_decoder(16#38#)) OR
 					(reg_q2649 AND symb_decoder(16#33#)) OR
 					(reg_q2649 AND symb_decoder(16#34#)) OR
 					(reg_q2649 AND symb_decoder(16#37#)) OR
 					(reg_q2649 AND symb_decoder(16#32#)) OR
 					(reg_q2649 AND symb_decoder(16#31#));
reg_q1457_in <= (reg_q1455 AND symb_decoder(16#4f#)) OR
 					(reg_q1455 AND symb_decoder(16#6f#));
reg_q1411_in <= (reg_q1409 AND symb_decoder(16#54#)) OR
 					(reg_q1409 AND symb_decoder(16#74#));
reg_q2064_in <= (reg_q2062 AND symb_decoder(16#49#)) OR
 					(reg_q2062 AND symb_decoder(16#69#));
reg_q1820_in <= (reg_q1818 AND symb_decoder(16#31#));
reg_q1463_in <= (reg_q1461 AND symb_decoder(16#6c#)) OR
 					(reg_q1461 AND symb_decoder(16#4c#));
reg_q2118_in <= (reg_q2116 AND symb_decoder(16#69#)) OR
 					(reg_q2116 AND symb_decoder(16#49#));
reg_q294_in <= (reg_q292 AND symb_decoder(16#77#)) OR
 					(reg_q292 AND symb_decoder(16#57#));
reg_q1034_in <= (reg_q1032 AND symb_decoder(16#32#));
reg_q2673_in <= (reg_q2671 AND symb_decoder(16#39#)) OR
 					(reg_q2671 AND symb_decoder(16#35#)) OR
 					(reg_q2671 AND symb_decoder(16#38#)) OR
 					(reg_q2671 AND symb_decoder(16#30#)) OR
 					(reg_q2671 AND symb_decoder(16#32#)) OR
 					(reg_q2671 AND symb_decoder(16#31#)) OR
 					(reg_q2671 AND symb_decoder(16#37#)) OR
 					(reg_q2671 AND symb_decoder(16#33#)) OR
 					(reg_q2671 AND symb_decoder(16#36#)) OR
 					(reg_q2671 AND symb_decoder(16#34#)) OR
 					(reg_q2673 AND symb_decoder(16#39#)) OR
 					(reg_q2673 AND symb_decoder(16#34#)) OR
 					(reg_q2673 AND symb_decoder(16#32#)) OR
 					(reg_q2673 AND symb_decoder(16#35#)) OR
 					(reg_q2673 AND symb_decoder(16#31#)) OR
 					(reg_q2673 AND symb_decoder(16#30#)) OR
 					(reg_q2673 AND symb_decoder(16#38#)) OR
 					(reg_q2673 AND symb_decoder(16#33#)) OR
 					(reg_q2673 AND symb_decoder(16#37#)) OR
 					(reg_q2673 AND symb_decoder(16#36#));
reg_q2635_in <= (reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2633 AND symb_decoder(16#7c#));
reg_q2637_in <= (reg_q2635 AND symb_decoder(16#39#)) OR
 					(reg_q2635 AND symb_decoder(16#36#)) OR
 					(reg_q2635 AND symb_decoder(16#32#)) OR
 					(reg_q2635 AND symb_decoder(16#38#)) OR
 					(reg_q2635 AND symb_decoder(16#37#)) OR
 					(reg_q2635 AND symb_decoder(16#34#)) OR
 					(reg_q2635 AND symb_decoder(16#33#)) OR
 					(reg_q2635 AND symb_decoder(16#31#)) OR
 					(reg_q2635 AND symb_decoder(16#30#)) OR
 					(reg_q2635 AND symb_decoder(16#35#)) OR
 					(reg_q2637 AND symb_decoder(16#34#)) OR
 					(reg_q2637 AND symb_decoder(16#31#)) OR
 					(reg_q2637 AND symb_decoder(16#38#)) OR
 					(reg_q2637 AND symb_decoder(16#33#)) OR
 					(reg_q2637 AND symb_decoder(16#30#)) OR
 					(reg_q2637 AND symb_decoder(16#35#)) OR
 					(reg_q2637 AND symb_decoder(16#39#)) OR
 					(reg_q2637 AND symb_decoder(16#37#)) OR
 					(reg_q2637 AND symb_decoder(16#36#)) OR
 					(reg_q2637 AND symb_decoder(16#32#));
reg_q2060_in <= (reg_q2058 AND symb_decoder(16#46#)) OR
 					(reg_q2058 AND symb_decoder(16#66#));
reg_q2062_in <= (reg_q2060 AND symb_decoder(16#72#)) OR
 					(reg_q2060 AND symb_decoder(16#52#));
reg_q1369_in <= (reg_q1367 AND symb_decoder(16#49#)) OR
 					(reg_q1367 AND symb_decoder(16#69#));
reg_q1636_in <= (reg_q1634 AND symb_decoder(16#49#)) OR
 					(reg_q1634 AND symb_decoder(16#69#));
reg_q2645_in <= (reg_q2643 AND symb_decoder(16#30#)) OR
 					(reg_q2643 AND symb_decoder(16#35#)) OR
 					(reg_q2643 AND symb_decoder(16#39#)) OR
 					(reg_q2643 AND symb_decoder(16#38#)) OR
 					(reg_q2643 AND symb_decoder(16#37#)) OR
 					(reg_q2643 AND symb_decoder(16#32#)) OR
 					(reg_q2643 AND symb_decoder(16#31#)) OR
 					(reg_q2643 AND symb_decoder(16#34#)) OR
 					(reg_q2643 AND symb_decoder(16#33#)) OR
 					(reg_q2643 AND symb_decoder(16#36#)) OR
 					(reg_q2645 AND symb_decoder(16#34#)) OR
 					(reg_q2645 AND symb_decoder(16#33#)) OR
 					(reg_q2645 AND symb_decoder(16#38#)) OR
 					(reg_q2645 AND symb_decoder(16#35#)) OR
 					(reg_q2645 AND symb_decoder(16#37#)) OR
 					(reg_q2645 AND symb_decoder(16#36#)) OR
 					(reg_q2645 AND symb_decoder(16#31#)) OR
 					(reg_q2645 AND symb_decoder(16#32#)) OR
 					(reg_q2645 AND symb_decoder(16#30#)) OR
 					(reg_q2645 AND symb_decoder(16#39#));
reg_q2433_in <= (reg_q2429 AND symb_decoder(16#3c#)) OR
 					(reg_q2447 AND symb_decoder(16#3c#));
reg_q1399_in <= (reg_q1397 AND symb_decoder(16#65#)) OR
 					(reg_q1397 AND symb_decoder(16#45#));
reg_q2239_in <= (reg_q2237 AND symb_decoder(16#3b#));
reg_q2122_in <= (reg_q2120 AND symb_decoder(16#4b#)) OR
 					(reg_q2120 AND symb_decoder(16#6b#));
reg_q1578_in <= (reg_q1576 AND symb_decoder(16#70#)) OR
 					(reg_q1576 AND symb_decoder(16#50#));
reg_q1848_in <= (reg_q1846 AND symb_decoder(16#49#)) OR
 					(reg_q1846 AND symb_decoder(16#69#));
reg_q1389_in <= (reg_q1387 AND symb_decoder(16#6f#)) OR
 					(reg_q1387 AND symb_decoder(16#4f#));
reg_q1385_in <= (reg_q1383 AND symb_decoder(16#65#)) OR
 					(reg_q1383 AND symb_decoder(16#45#));
reg_q1387_in <= (reg_q1385 AND symb_decoder(16#4d#)) OR
 					(reg_q1385 AND symb_decoder(16#6d#));
reg_q1644_in <= (reg_q1642 AND symb_decoder(16#75#)) OR
 					(reg_q1642 AND symb_decoder(16#55#));
reg_q1530_in <= (reg_q1528 AND symb_decoder(16#44#)) OR
 					(reg_q1528 AND symb_decoder(16#64#));
reg_q1592_in <= (reg_q1590 AND symb_decoder(16#64#)) OR
 					(reg_q1590 AND symb_decoder(16#44#));
reg_q1884_in <= (reg_q1882 AND symb_decoder(16#32#));
reg_q1026_in <= (reg_q1024 AND symb_decoder(16#68#));
reg_q2639_in <= (reg_q2637 AND symb_decoder(16#2e#));
reg_q2074_in <= (reg_q2072 AND symb_decoder(16#68#)) OR
 					(reg_q2072 AND symb_decoder(16#48#));
reg_q1818_in <= (reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q1816 AND symb_decoder(16#23#));
reg_q1461_in <= (reg_q1459 AND symb_decoder(16#41#)) OR
 					(reg_q1459 AND symb_decoder(16#61#));
reg_q1634_in <= (reg_q1632 AND symb_decoder(16#2d#));
reg_q1467_in <= (reg_q1465 AND symb_decoder(16#64#)) OR
 					(reg_q1465 AND symb_decoder(16#44#));
reg_q2172_in <= (reg_q2170 AND symb_decoder(16#43#)) OR
 					(reg_q2170 AND symb_decoder(16#63#));
reg_q1640_in <= (reg_q1638 AND symb_decoder(16#63#)) OR
 					(reg_q1638 AND symb_decoder(16#43#));
reg_q1642_in <= (reg_q1640 AND symb_decoder(16#4c#)) OR
 					(reg_q1640 AND symb_decoder(16#6c#));
reg_q1594_in <= (reg_q1592 AND symb_decoder(16#45#)) OR
 					(reg_q1592 AND symb_decoder(16#65#));
reg_q1365_in <= (reg_q1363 AND symb_decoder(16#63#)) OR
 					(reg_q1363 AND symb_decoder(16#43#));
reg_q2538_in <= (reg_q2534 AND symb_decoder(16#5c#)) OR
 					(reg_q2552 AND symb_decoder(16#5c#));
reg_q1598_in <= (reg_q1596 AND symb_decoder(16#2f#));
reg_q1270_in <= (reg_q1268 AND symb_decoder(16#49#)) OR
 					(reg_q1268 AND symb_decoder(16#69#));
reg_q411_in <= (reg_q409 AND symb_decoder(16#77#)) OR
 					(reg_q409 AND symb_decoder(16#57#));
reg_q1453_in <= (reg_q1451 AND symb_decoder(16#54#)) OR
 					(reg_q1451 AND symb_decoder(16#74#));
reg_q1469_in <= (reg_q1467 AND symb_decoder(16#61#)) OR
 					(reg_q1467 AND symb_decoder(16#41#));
reg_q1534_in <= (reg_q1532 AND symb_decoder(16#57#)) OR
 					(reg_q1532 AND symb_decoder(16#77#));
reg_q461_in <= (reg_q459 AND symb_decoder(16#77#)) OR
 					(reg_q459 AND symb_decoder(16#57#));
reg_q492_in <= (reg_q490 AND symb_decoder(16#3a#));
reg_q1973_in <= (reg_q1971 AND symb_decoder(16#2b#));
reg_q2160_in <= (reg_q2158 AND symb_decoder(16#65#)) OR
 					(reg_q2158 AND symb_decoder(16#45#));
reg_q1028_in <= (reg_q1026 AND symb_decoder(16#65#));
reg_q2164_in <= (reg_q2162 AND symb_decoder(16#44#)) OR
 					(reg_q2162 AND symb_decoder(16#64#));
reg_fullgraph55_init <= "0000000";

reg_fullgraph55_sel <= "000000000000000000000000000000000000000000000000000000000000" & reg_q2164_in & reg_q1028_in & reg_q2160_in & reg_q1973_in & reg_q492_in & reg_q461_in & reg_q1534_in & reg_q1469_in & reg_q1453_in & reg_q411_in & reg_q1270_in & reg_q1598_in & reg_q2538_in & reg_q1365_in & reg_q1594_in & reg_q1642_in & reg_q1640_in & reg_q2172_in & reg_q1467_in & reg_q1634_in & reg_q1461_in & reg_q1818_in & reg_q2074_in & reg_q2639_in & reg_q1026_in & reg_q1884_in & reg_q1592_in & reg_q1530_in & reg_q1644_in & reg_q1387_in & reg_q1385_in & reg_q1389_in & reg_q1848_in & reg_q1578_in & reg_q2122_in & reg_q2239_in & reg_q1399_in & reg_q2433_in & reg_q2645_in & reg_q1636_in & reg_q1369_in & reg_q2062_in & reg_q2060_in & reg_q2637_in & reg_q2635_in & reg_q2673_in & reg_q1034_in & reg_q294_in & reg_q2118_in & reg_q1463_in & reg_q1820_in & reg_q2064_in & reg_q1411_in & reg_q1457_in & reg_q2649_in & reg_q2647_in & reg_q2237_in & reg_q2241_in & reg_q296_in & reg_q2643_in & reg_q1465_in & reg_q2116_in & reg_q435_in & reg_q2641_in & reg_q2435_in & reg_q342_in & reg_q606_in & reg_q2080_in;

	--coder fullgraph55
with reg_fullgraph55_sel select
reg_fullgraph55_in <=
	"0000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001",
	"0000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010",
	"0000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100",
	"0000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000",
	"0000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000",
	"0000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000",
	"0000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000",
	"0001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000",
	"0001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
	"0001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000",
	"0001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000",
	"0001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000",
	"0001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000",
	"0001110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000",
	"0001111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000",
	"0010000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000",
	"0010001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000",
	"0010010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000",
	"0010011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000",
	"0010100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000",
	"0010101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000",
	"0010110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000",
	"0010111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000",
	"0011000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000",
	"0011001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000",
	"0011010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000",
	"0011011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000",
	"0011100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000",
	"0011101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000",
	"0011110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000",
	"0011111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000",
	"0100000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000",
	"0100001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000",
	"0100010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000",
	"0100011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000",
	"0100100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000",
	"0100101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000",
	"0100110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000",
	"0100111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000",
	"0101000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000",
	"0101001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000",
	"0101010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000",
	"0101011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000",
	"0101100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000",
	"0101101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"0101110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000",
	"0101111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000",
	"0110000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000",
	"0110001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000",
	"0110010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000",
	"0110011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000",
	"0110100" when "00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000",
	"0110101" when "00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000",
	"0110110" when "00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000",
	"0110111" when "00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000",
	"0111000" when "00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000",
	"0111001" when "00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000",
	"0111010" when "00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000",
	"0111011" when "00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000",
	"0111100" when "00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000",
	"0111101" when "00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000",
	"0111110" when "00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000",
	"0111111" when "00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000",
	"1000000" when "00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000",
	"1000001" when "00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000",
	"1000010" when "00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000",
	"1000011" when "00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000",
	"1000100" when "00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000",
	"0000000" when others;
 --end coder

	p_reg_fullgraph55: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph55 <= reg_fullgraph55_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph55 <= reg_fullgraph55_init;
        else
          reg_fullgraph55 <= reg_fullgraph55_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph55

		reg_q2080 <= '1' when reg_fullgraph55 = "0000001" else '0'; 
		reg_q606 <= '1' when reg_fullgraph55 = "0000010" else '0'; 
		reg_q342 <= '1' when reg_fullgraph55 = "0000011" else '0'; 
		reg_q2435 <= '1' when reg_fullgraph55 = "0000100" else '0'; 
		reg_q2641 <= '1' when reg_fullgraph55 = "0000101" else '0'; 
		reg_q435 <= '1' when reg_fullgraph55 = "0000110" else '0'; 
		reg_q2116 <= '1' when reg_fullgraph55 = "0000111" else '0'; 
		reg_q1465 <= '1' when reg_fullgraph55 = "0001000" else '0'; 
		reg_q2643 <= '1' when reg_fullgraph55 = "0001001" else '0'; 
		reg_q296 <= '1' when reg_fullgraph55 = "0001010" else '0'; 
		reg_q2241 <= '1' when reg_fullgraph55 = "0001011" else '0'; 
		reg_q2237 <= '1' when reg_fullgraph55 = "0001100" else '0'; 
		reg_q2647 <= '1' when reg_fullgraph55 = "0001101" else '0'; 
		reg_q2649 <= '1' when reg_fullgraph55 = "0001110" else '0'; 
		reg_q1457 <= '1' when reg_fullgraph55 = "0001111" else '0'; 
		reg_q1411 <= '1' when reg_fullgraph55 = "0010000" else '0'; 
		reg_q2064 <= '1' when reg_fullgraph55 = "0010001" else '0'; 
		reg_q1820 <= '1' when reg_fullgraph55 = "0010010" else '0'; 
		reg_q1463 <= '1' when reg_fullgraph55 = "0010011" else '0'; 
		reg_q2118 <= '1' when reg_fullgraph55 = "0010100" else '0'; 
		reg_q294 <= '1' when reg_fullgraph55 = "0010101" else '0'; 
		reg_q1034 <= '1' when reg_fullgraph55 = "0010110" else '0'; 
		reg_q2673 <= '1' when reg_fullgraph55 = "0010111" else '0'; 
		reg_q2635 <= '1' when reg_fullgraph55 = "0011000" else '0'; 
		reg_q2637 <= '1' when reg_fullgraph55 = "0011001" else '0'; 
		reg_q2060 <= '1' when reg_fullgraph55 = "0011010" else '0'; 
		reg_q2062 <= '1' when reg_fullgraph55 = "0011011" else '0'; 
		reg_q1369 <= '1' when reg_fullgraph55 = "0011100" else '0'; 
		reg_q1636 <= '1' when reg_fullgraph55 = "0011101" else '0'; 
		reg_q2645 <= '1' when reg_fullgraph55 = "0011110" else '0'; 
		reg_q2433 <= '1' when reg_fullgraph55 = "0011111" else '0'; 
		reg_q1399 <= '1' when reg_fullgraph55 = "0100000" else '0'; 
		reg_q2239 <= '1' when reg_fullgraph55 = "0100001" else '0'; 
		reg_q2122 <= '1' when reg_fullgraph55 = "0100010" else '0'; 
		reg_q1578 <= '1' when reg_fullgraph55 = "0100011" else '0'; 
		reg_q1848 <= '1' when reg_fullgraph55 = "0100100" else '0'; 
		reg_q1389 <= '1' when reg_fullgraph55 = "0100101" else '0'; 
		reg_q1385 <= '1' when reg_fullgraph55 = "0100110" else '0'; 
		reg_q1387 <= '1' when reg_fullgraph55 = "0100111" else '0'; 
		reg_q1644 <= '1' when reg_fullgraph55 = "0101000" else '0'; 
		reg_q1530 <= '1' when reg_fullgraph55 = "0101001" else '0'; 
		reg_q1592 <= '1' when reg_fullgraph55 = "0101010" else '0'; 
		reg_q1884 <= '1' when reg_fullgraph55 = "0101011" else '0'; 
		reg_q1026 <= '1' when reg_fullgraph55 = "0101100" else '0'; 
		reg_q2639 <= '1' when reg_fullgraph55 = "0101101" else '0'; 
		reg_q2074 <= '1' when reg_fullgraph55 = "0101110" else '0'; 
		reg_q1818 <= '1' when reg_fullgraph55 = "0101111" else '0'; 
		reg_q1461 <= '1' when reg_fullgraph55 = "0110000" else '0'; 
		reg_q1634 <= '1' when reg_fullgraph55 = "0110001" else '0'; 
		reg_q1467 <= '1' when reg_fullgraph55 = "0110010" else '0'; 
		reg_q2172 <= '1' when reg_fullgraph55 = "0110011" else '0'; 
		reg_q1640 <= '1' when reg_fullgraph55 = "0110100" else '0'; 
		reg_q1642 <= '1' when reg_fullgraph55 = "0110101" else '0'; 
		reg_q1594 <= '1' when reg_fullgraph55 = "0110110" else '0'; 
		reg_q1365 <= '1' when reg_fullgraph55 = "0110111" else '0'; 
		reg_q2538 <= '1' when reg_fullgraph55 = "0111000" else '0'; 
		reg_q1598 <= '1' when reg_fullgraph55 = "0111001" else '0'; 
		reg_q1270 <= '1' when reg_fullgraph55 = "0111010" else '0'; 
		reg_q411 <= '1' when reg_fullgraph55 = "0111011" else '0'; 
		reg_q1453 <= '1' when reg_fullgraph55 = "0111100" else '0'; 
		reg_q1469 <= '1' when reg_fullgraph55 = "0111101" else '0'; 
		reg_q1534 <= '1' when reg_fullgraph55 = "0111110" else '0'; 
		reg_q461 <= '1' when reg_fullgraph55 = "0111111" else '0'; 
		reg_q492 <= '1' when reg_fullgraph55 = "1000000" else '0'; 
		reg_q1973 <= '1' when reg_fullgraph55 = "1000001" else '0'; 
		reg_q2160 <= '1' when reg_fullgraph55 = "1000010" else '0'; 
		reg_q1028 <= '1' when reg_fullgraph55 = "1000011" else '0'; 
		reg_q2164 <= '1' when reg_fullgraph55 = "1000100" else '0'; 
--end decoder 

reg_q1522_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1522 AND symb_decoder(16#a0#)) OR
 					(reg_q1522 AND symb_decoder(16#c1#)) OR
 					(reg_q1522 AND symb_decoder(16#b1#)) OR
 					(reg_q1522 AND symb_decoder(16#e9#)) OR
 					(reg_q1522 AND symb_decoder(16#16#)) OR
 					(reg_q1522 AND symb_decoder(16#0e#)) OR
 					(reg_q1522 AND symb_decoder(16#b0#)) OR
 					(reg_q1522 AND symb_decoder(16#73#)) OR
 					(reg_q1522 AND symb_decoder(16#f3#)) OR
 					(reg_q1522 AND symb_decoder(16#15#)) OR
 					(reg_q1522 AND symb_decoder(16#ad#)) OR
 					(reg_q1522 AND symb_decoder(16#0c#)) OR
 					(reg_q1522 AND symb_decoder(16#4f#)) OR
 					(reg_q1522 AND symb_decoder(16#7f#)) OR
 					(reg_q1522 AND symb_decoder(16#88#)) OR
 					(reg_q1522 AND symb_decoder(16#30#)) OR
 					(reg_q1522 AND symb_decoder(16#b7#)) OR
 					(reg_q1522 AND symb_decoder(16#a2#)) OR
 					(reg_q1522 AND symb_decoder(16#63#)) OR
 					(reg_q1522 AND symb_decoder(16#8e#)) OR
 					(reg_q1522 AND symb_decoder(16#94#)) OR
 					(reg_q1522 AND symb_decoder(16#f4#)) OR
 					(reg_q1522 AND symb_decoder(16#7c#)) OR
 					(reg_q1522 AND symb_decoder(16#2e#)) OR
 					(reg_q1522 AND symb_decoder(16#6e#)) OR
 					(reg_q1522 AND symb_decoder(16#07#)) OR
 					(reg_q1522 AND symb_decoder(16#2c#)) OR
 					(reg_q1522 AND symb_decoder(16#c0#)) OR
 					(reg_q1522 AND symb_decoder(16#5a#)) OR
 					(reg_q1522 AND symb_decoder(16#86#)) OR
 					(reg_q1522 AND symb_decoder(16#6a#)) OR
 					(reg_q1522 AND symb_decoder(16#66#)) OR
 					(reg_q1522 AND symb_decoder(16#0a#)) OR
 					(reg_q1522 AND symb_decoder(16#62#)) OR
 					(reg_q1522 AND symb_decoder(16#7e#)) OR
 					(reg_q1522 AND symb_decoder(16#e4#)) OR
 					(reg_q1522 AND symb_decoder(16#5c#)) OR
 					(reg_q1522 AND symb_decoder(16#82#)) OR
 					(reg_q1522 AND symb_decoder(16#ce#)) OR
 					(reg_q1522 AND symb_decoder(16#fe#)) OR
 					(reg_q1522 AND symb_decoder(16#08#)) OR
 					(reg_q1522 AND symb_decoder(16#85#)) OR
 					(reg_q1522 AND symb_decoder(16#9a#)) OR
 					(reg_q1522 AND symb_decoder(16#db#)) OR
 					(reg_q1522 AND symb_decoder(16#b4#)) OR
 					(reg_q1522 AND symb_decoder(16#92#)) OR
 					(reg_q1522 AND symb_decoder(16#6d#)) OR
 					(reg_q1522 AND symb_decoder(16#41#)) OR
 					(reg_q1522 AND symb_decoder(16#3f#)) OR
 					(reg_q1522 AND symb_decoder(16#39#)) OR
 					(reg_q1522 AND symb_decoder(16#72#)) OR
 					(reg_q1522 AND symb_decoder(16#97#)) OR
 					(reg_q1522 AND symb_decoder(16#cc#)) OR
 					(reg_q1522 AND symb_decoder(16#71#)) OR
 					(reg_q1522 AND symb_decoder(16#bc#)) OR
 					(reg_q1522 AND symb_decoder(16#60#)) OR
 					(reg_q1522 AND symb_decoder(16#04#)) OR
 					(reg_q1522 AND symb_decoder(16#c4#)) OR
 					(reg_q1522 AND symb_decoder(16#0d#)) OR
 					(reg_q1522 AND symb_decoder(16#23#)) OR
 					(reg_q1522 AND symb_decoder(16#02#)) OR
 					(reg_q1522 AND symb_decoder(16#c9#)) OR
 					(reg_q1522 AND symb_decoder(16#74#)) OR
 					(reg_q1522 AND symb_decoder(16#83#)) OR
 					(reg_q1522 AND symb_decoder(16#43#)) OR
 					(reg_q1522 AND symb_decoder(16#ba#)) OR
 					(reg_q1522 AND symb_decoder(16#67#)) OR
 					(reg_q1522 AND symb_decoder(16#26#)) OR
 					(reg_q1522 AND symb_decoder(16#b3#)) OR
 					(reg_q1522 AND symb_decoder(16#5f#)) OR
 					(reg_q1522 AND symb_decoder(16#d2#)) OR
 					(reg_q1522 AND symb_decoder(16#4a#)) OR
 					(reg_q1522 AND symb_decoder(16#a8#)) OR
 					(reg_q1522 AND symb_decoder(16#6f#)) OR
 					(reg_q1522 AND symb_decoder(16#2b#)) OR
 					(reg_q1522 AND symb_decoder(16#28#)) OR
 					(reg_q1522 AND symb_decoder(16#64#)) OR
 					(reg_q1522 AND symb_decoder(16#ca#)) OR
 					(reg_q1522 AND symb_decoder(16#b8#)) OR
 					(reg_q1522 AND symb_decoder(16#ea#)) OR
 					(reg_q1522 AND symb_decoder(16#bd#)) OR
 					(reg_q1522 AND symb_decoder(16#af#)) OR
 					(reg_q1522 AND symb_decoder(16#fd#)) OR
 					(reg_q1522 AND symb_decoder(16#77#)) OR
 					(reg_q1522 AND symb_decoder(16#42#)) OR
 					(reg_q1522 AND symb_decoder(16#d7#)) OR
 					(reg_q1522 AND symb_decoder(16#0f#)) OR
 					(reg_q1522 AND symb_decoder(16#44#)) OR
 					(reg_q1522 AND symb_decoder(16#57#)) OR
 					(reg_q1522 AND symb_decoder(16#0b#)) OR
 					(reg_q1522 AND symb_decoder(16#e2#)) OR
 					(reg_q1522 AND symb_decoder(16#55#)) OR
 					(reg_q1522 AND symb_decoder(16#c6#)) OR
 					(reg_q1522 AND symb_decoder(16#70#)) OR
 					(reg_q1522 AND symb_decoder(16#9c#)) OR
 					(reg_q1522 AND symb_decoder(16#cf#)) OR
 					(reg_q1522 AND symb_decoder(16#10#)) OR
 					(reg_q1522 AND symb_decoder(16#31#)) OR
 					(reg_q1522 AND symb_decoder(16#52#)) OR
 					(reg_q1522 AND symb_decoder(16#90#)) OR
 					(reg_q1522 AND symb_decoder(16#59#)) OR
 					(reg_q1522 AND symb_decoder(16#dd#)) OR
 					(reg_q1522 AND symb_decoder(16#ae#)) OR
 					(reg_q1522 AND symb_decoder(16#1a#)) OR
 					(reg_q1522 AND symb_decoder(16#1f#)) OR
 					(reg_q1522 AND symb_decoder(16#34#)) OR
 					(reg_q1522 AND symb_decoder(16#68#)) OR
 					(reg_q1522 AND symb_decoder(16#38#)) OR
 					(reg_q1522 AND symb_decoder(16#8d#)) OR
 					(reg_q1522 AND symb_decoder(16#17#)) OR
 					(reg_q1522 AND symb_decoder(16#78#)) OR
 					(reg_q1522 AND symb_decoder(16#2a#)) OR
 					(reg_q1522 AND symb_decoder(16#fa#)) OR
 					(reg_q1522 AND symb_decoder(16#98#)) OR
 					(reg_q1522 AND symb_decoder(16#c2#)) OR
 					(reg_q1522 AND symb_decoder(16#4d#)) OR
 					(reg_q1522 AND symb_decoder(16#29#)) OR
 					(reg_q1522 AND symb_decoder(16#bb#)) OR
 					(reg_q1522 AND symb_decoder(16#fb#)) OR
 					(reg_q1522 AND symb_decoder(16#ab#)) OR
 					(reg_q1522 AND symb_decoder(16#3c#)) OR
 					(reg_q1522 AND symb_decoder(16#51#)) OR
 					(reg_q1522 AND symb_decoder(16#cd#)) OR
 					(reg_q1522 AND symb_decoder(16#56#)) OR
 					(reg_q1522 AND symb_decoder(16#8b#)) OR
 					(reg_q1522 AND symb_decoder(16#65#)) OR
 					(reg_q1522 AND symb_decoder(16#05#)) OR
 					(reg_q1522 AND symb_decoder(16#69#)) OR
 					(reg_q1522 AND symb_decoder(16#32#)) OR
 					(reg_q1522 AND symb_decoder(16#4b#)) OR
 					(reg_q1522 AND symb_decoder(16#1b#)) OR
 					(reg_q1522 AND symb_decoder(16#5d#)) OR
 					(reg_q1522 AND symb_decoder(16#4e#)) OR
 					(reg_q1522 AND symb_decoder(16#a1#)) OR
 					(reg_q1522 AND symb_decoder(16#21#)) OR
 					(reg_q1522 AND symb_decoder(16#00#)) OR
 					(reg_q1522 AND symb_decoder(16#8a#)) OR
 					(reg_q1522 AND symb_decoder(16#f5#)) OR
 					(reg_q1522 AND symb_decoder(16#f1#)) OR
 					(reg_q1522 AND symb_decoder(16#61#)) OR
 					(reg_q1522 AND symb_decoder(16#2d#)) OR
 					(reg_q1522 AND symb_decoder(16#09#)) OR
 					(reg_q1522 AND symb_decoder(16#75#)) OR
 					(reg_q1522 AND symb_decoder(16#aa#)) OR
 					(reg_q1522 AND symb_decoder(16#3d#)) OR
 					(reg_q1522 AND symb_decoder(16#7d#)) OR
 					(reg_q1522 AND symb_decoder(16#d6#)) OR
 					(reg_q1522 AND symb_decoder(16#a3#)) OR
 					(reg_q1522 AND symb_decoder(16#fc#)) OR
 					(reg_q1522 AND symb_decoder(16#50#)) OR
 					(reg_q1522 AND symb_decoder(16#9b#)) OR
 					(reg_q1522 AND symb_decoder(16#22#)) OR
 					(reg_q1522 AND symb_decoder(16#18#)) OR
 					(reg_q1522 AND symb_decoder(16#2f#)) OR
 					(reg_q1522 AND symb_decoder(16#3b#)) OR
 					(reg_q1522 AND symb_decoder(16#f2#)) OR
 					(reg_q1522 AND symb_decoder(16#96#)) OR
 					(reg_q1522 AND symb_decoder(16#91#)) OR
 					(reg_q1522 AND symb_decoder(16#24#)) OR
 					(reg_q1522 AND symb_decoder(16#eb#)) OR
 					(reg_q1522 AND symb_decoder(16#b9#)) OR
 					(reg_q1522 AND symb_decoder(16#1d#)) OR
 					(reg_q1522 AND symb_decoder(16#35#)) OR
 					(reg_q1522 AND symb_decoder(16#ed#)) OR
 					(reg_q1522 AND symb_decoder(16#45#)) OR
 					(reg_q1522 AND symb_decoder(16#36#)) OR
 					(reg_q1522 AND symb_decoder(16#f9#)) OR
 					(reg_q1522 AND symb_decoder(16#54#)) OR
 					(reg_q1522 AND symb_decoder(16#d1#)) OR
 					(reg_q1522 AND symb_decoder(16#8f#)) OR
 					(reg_q1522 AND symb_decoder(16#da#)) OR
 					(reg_q1522 AND symb_decoder(16#3e#)) OR
 					(reg_q1522 AND symb_decoder(16#93#)) OR
 					(reg_q1522 AND symb_decoder(16#25#)) OR
 					(reg_q1522 AND symb_decoder(16#6c#)) OR
 					(reg_q1522 AND symb_decoder(16#12#)) OR
 					(reg_q1522 AND symb_decoder(16#14#)) OR
 					(reg_q1522 AND symb_decoder(16#4c#)) OR
 					(reg_q1522 AND symb_decoder(16#a4#)) OR
 					(reg_q1522 AND symb_decoder(16#5b#)) OR
 					(reg_q1522 AND symb_decoder(16#ac#)) OR
 					(reg_q1522 AND symb_decoder(16#87#)) OR
 					(reg_q1522 AND symb_decoder(16#c7#)) OR
 					(reg_q1522 AND symb_decoder(16#7b#)) OR
 					(reg_q1522 AND symb_decoder(16#1c#)) OR
 					(reg_q1522 AND symb_decoder(16#19#)) OR
 					(reg_q1522 AND symb_decoder(16#f6#)) OR
 					(reg_q1522 AND symb_decoder(16#3a#)) OR
 					(reg_q1522 AND symb_decoder(16#9e#)) OR
 					(reg_q1522 AND symb_decoder(16#27#)) OR
 					(reg_q1522 AND symb_decoder(16#d9#)) OR
 					(reg_q1522 AND symb_decoder(16#ff#)) OR
 					(reg_q1522 AND symb_decoder(16#df#)) OR
 					(reg_q1522 AND symb_decoder(16#f7#)) OR
 					(reg_q1522 AND symb_decoder(16#ef#)) OR
 					(reg_q1522 AND symb_decoder(16#01#)) OR
 					(reg_q1522 AND symb_decoder(16#37#)) OR
 					(reg_q1522 AND symb_decoder(16#cb#)) OR
 					(reg_q1522 AND symb_decoder(16#d0#)) OR
 					(reg_q1522 AND symb_decoder(16#48#)) OR
 					(reg_q1522 AND symb_decoder(16#a5#)) OR
 					(reg_q1522 AND symb_decoder(16#80#)) OR
 					(reg_q1522 AND symb_decoder(16#11#)) OR
 					(reg_q1522 AND symb_decoder(16#20#)) OR
 					(reg_q1522 AND symb_decoder(16#89#)) OR
 					(reg_q1522 AND symb_decoder(16#d4#)) OR
 					(reg_q1522 AND symb_decoder(16#49#)) OR
 					(reg_q1522 AND symb_decoder(16#b2#)) OR
 					(reg_q1522 AND symb_decoder(16#58#)) OR
 					(reg_q1522 AND symb_decoder(16#81#)) OR
 					(reg_q1522 AND symb_decoder(16#79#)) OR
 					(reg_q1522 AND symb_decoder(16#8c#)) OR
 					(reg_q1522 AND symb_decoder(16#84#)) OR
 					(reg_q1522 AND symb_decoder(16#76#)) OR
 					(reg_q1522 AND symb_decoder(16#c3#)) OR
 					(reg_q1522 AND symb_decoder(16#e5#)) OR
 					(reg_q1522 AND symb_decoder(16#ec#)) OR
 					(reg_q1522 AND symb_decoder(16#ee#)) OR
 					(reg_q1522 AND symb_decoder(16#c5#)) OR
 					(reg_q1522 AND symb_decoder(16#13#)) OR
 					(reg_q1522 AND symb_decoder(16#be#)) OR
 					(reg_q1522 AND symb_decoder(16#b6#)) OR
 					(reg_q1522 AND symb_decoder(16#06#)) OR
 					(reg_q1522 AND symb_decoder(16#dc#)) OR
 					(reg_q1522 AND symb_decoder(16#b5#)) OR
 					(reg_q1522 AND symb_decoder(16#e3#)) OR
 					(reg_q1522 AND symb_decoder(16#5e#)) OR
 					(reg_q1522 AND symb_decoder(16#46#)) OR
 					(reg_q1522 AND symb_decoder(16#e0#)) OR
 					(reg_q1522 AND symb_decoder(16#53#)) OR
 					(reg_q1522 AND symb_decoder(16#d8#)) OR
 					(reg_q1522 AND symb_decoder(16#95#)) OR
 					(reg_q1522 AND symb_decoder(16#d3#)) OR
 					(reg_q1522 AND symb_decoder(16#a9#)) OR
 					(reg_q1522 AND symb_decoder(16#f8#)) OR
 					(reg_q1522 AND symb_decoder(16#a7#)) OR
 					(reg_q1522 AND symb_decoder(16#7a#)) OR
 					(reg_q1522 AND symb_decoder(16#bf#)) OR
 					(reg_q1522 AND symb_decoder(16#6b#)) OR
 					(reg_q1522 AND symb_decoder(16#9d#)) OR
 					(reg_q1522 AND symb_decoder(16#c8#)) OR
 					(reg_q1522 AND symb_decoder(16#99#)) OR
 					(reg_q1522 AND symb_decoder(16#33#)) OR
 					(reg_q1522 AND symb_decoder(16#e1#)) OR
 					(reg_q1522 AND symb_decoder(16#e7#)) OR
 					(reg_q1522 AND symb_decoder(16#d5#)) OR
 					(reg_q1522 AND symb_decoder(16#e8#)) OR
 					(reg_q1522 AND symb_decoder(16#9f#)) OR
 					(reg_q1522 AND symb_decoder(16#1e#)) OR
 					(reg_q1522 AND symb_decoder(16#e6#)) OR
 					(reg_q1522 AND symb_decoder(16#40#)) OR
 					(reg_q1522 AND symb_decoder(16#de#)) OR
 					(reg_q1522 AND symb_decoder(16#47#)) OR
 					(reg_q1522 AND symb_decoder(16#03#)) OR
 					(reg_q1522 AND symb_decoder(16#f0#)) OR
 					(reg_q1522 AND symb_decoder(16#a6#));
reg_q1522_init <= '0' ;
	p_reg_q1522: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1522 <= reg_q1522_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1522 <= reg_q1522_init;
        else
          reg_q1522 <= reg_q1522_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q661_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q661 AND symb_decoder(16#d1#)) OR
 					(reg_q661 AND symb_decoder(16#18#)) OR
 					(reg_q661 AND symb_decoder(16#fd#)) OR
 					(reg_q661 AND symb_decoder(16#cc#)) OR
 					(reg_q661 AND symb_decoder(16#7c#)) OR
 					(reg_q661 AND symb_decoder(16#3c#)) OR
 					(reg_q661 AND symb_decoder(16#75#)) OR
 					(reg_q661 AND symb_decoder(16#e3#)) OR
 					(reg_q661 AND symb_decoder(16#67#)) OR
 					(reg_q661 AND symb_decoder(16#d5#)) OR
 					(reg_q661 AND symb_decoder(16#26#)) OR
 					(reg_q661 AND symb_decoder(16#ff#)) OR
 					(reg_q661 AND symb_decoder(16#09#)) OR
 					(reg_q661 AND symb_decoder(16#1a#)) OR
 					(reg_q661 AND symb_decoder(16#c7#)) OR
 					(reg_q661 AND symb_decoder(16#7d#)) OR
 					(reg_q661 AND symb_decoder(16#49#)) OR
 					(reg_q661 AND symb_decoder(16#38#)) OR
 					(reg_q661 AND symb_decoder(16#5b#)) OR
 					(reg_q661 AND symb_decoder(16#ea#)) OR
 					(reg_q661 AND symb_decoder(16#f1#)) OR
 					(reg_q661 AND symb_decoder(16#b1#)) OR
 					(reg_q661 AND symb_decoder(16#79#)) OR
 					(reg_q661 AND symb_decoder(16#20#)) OR
 					(reg_q661 AND symb_decoder(16#ef#)) OR
 					(reg_q661 AND symb_decoder(16#1f#)) OR
 					(reg_q661 AND symb_decoder(16#93#)) OR
 					(reg_q661 AND symb_decoder(16#ae#)) OR
 					(reg_q661 AND symb_decoder(16#35#)) OR
 					(reg_q661 AND symb_decoder(16#3b#)) OR
 					(reg_q661 AND symb_decoder(16#fb#)) OR
 					(reg_q661 AND symb_decoder(16#ed#)) OR
 					(reg_q661 AND symb_decoder(16#c6#)) OR
 					(reg_q661 AND symb_decoder(16#14#)) OR
 					(reg_q661 AND symb_decoder(16#7f#)) OR
 					(reg_q661 AND symb_decoder(16#0d#)) OR
 					(reg_q661 AND symb_decoder(16#6e#)) OR
 					(reg_q661 AND symb_decoder(16#dd#)) OR
 					(reg_q661 AND symb_decoder(16#df#)) OR
 					(reg_q661 AND symb_decoder(16#23#)) OR
 					(reg_q661 AND symb_decoder(16#a3#)) OR
 					(reg_q661 AND symb_decoder(16#4f#)) OR
 					(reg_q661 AND symb_decoder(16#ce#)) OR
 					(reg_q661 AND symb_decoder(16#5d#)) OR
 					(reg_q661 AND symb_decoder(16#10#)) OR
 					(reg_q661 AND symb_decoder(16#88#)) OR
 					(reg_q661 AND symb_decoder(16#d4#)) OR
 					(reg_q661 AND symb_decoder(16#2f#)) OR
 					(reg_q661 AND symb_decoder(16#32#)) OR
 					(reg_q661 AND symb_decoder(16#74#)) OR
 					(reg_q661 AND symb_decoder(16#e1#)) OR
 					(reg_q661 AND symb_decoder(16#4e#)) OR
 					(reg_q661 AND symb_decoder(16#90#)) OR
 					(reg_q661 AND symb_decoder(16#55#)) OR
 					(reg_q661 AND symb_decoder(16#89#)) OR
 					(reg_q661 AND symb_decoder(16#a0#)) OR
 					(reg_q661 AND symb_decoder(16#4a#)) OR
 					(reg_q661 AND symb_decoder(16#f8#)) OR
 					(reg_q661 AND symb_decoder(16#b3#)) OR
 					(reg_q661 AND symb_decoder(16#a2#)) OR
 					(reg_q661 AND symb_decoder(16#95#)) OR
 					(reg_q661 AND symb_decoder(16#17#)) OR
 					(reg_q661 AND symb_decoder(16#b4#)) OR
 					(reg_q661 AND symb_decoder(16#e8#)) OR
 					(reg_q661 AND symb_decoder(16#4b#)) OR
 					(reg_q661 AND symb_decoder(16#61#)) OR
 					(reg_q661 AND symb_decoder(16#1c#)) OR
 					(reg_q661 AND symb_decoder(16#e6#)) OR
 					(reg_q661 AND symb_decoder(16#bb#)) OR
 					(reg_q661 AND symb_decoder(16#99#)) OR
 					(reg_q661 AND symb_decoder(16#12#)) OR
 					(reg_q661 AND symb_decoder(16#72#)) OR
 					(reg_q661 AND symb_decoder(16#84#)) OR
 					(reg_q661 AND symb_decoder(16#c5#)) OR
 					(reg_q661 AND symb_decoder(16#68#)) OR
 					(reg_q661 AND symb_decoder(16#8a#)) OR
 					(reg_q661 AND symb_decoder(16#dc#)) OR
 					(reg_q661 AND symb_decoder(16#8e#)) OR
 					(reg_q661 AND symb_decoder(16#a8#)) OR
 					(reg_q661 AND symb_decoder(16#25#)) OR
 					(reg_q661 AND symb_decoder(16#2c#)) OR
 					(reg_q661 AND symb_decoder(16#5e#)) OR
 					(reg_q661 AND symb_decoder(16#d9#)) OR
 					(reg_q661 AND symb_decoder(16#4d#)) OR
 					(reg_q661 AND symb_decoder(16#ab#)) OR
 					(reg_q661 AND symb_decoder(16#2d#)) OR
 					(reg_q661 AND symb_decoder(16#c4#)) OR
 					(reg_q661 AND symb_decoder(16#e4#)) OR
 					(reg_q661 AND symb_decoder(16#37#)) OR
 					(reg_q661 AND symb_decoder(16#2e#)) OR
 					(reg_q661 AND symb_decoder(16#21#)) OR
 					(reg_q661 AND symb_decoder(16#01#)) OR
 					(reg_q661 AND symb_decoder(16#16#)) OR
 					(reg_q661 AND symb_decoder(16#1e#)) OR
 					(reg_q661 AND symb_decoder(16#fa#)) OR
 					(reg_q661 AND symb_decoder(16#07#)) OR
 					(reg_q661 AND symb_decoder(16#c9#)) OR
 					(reg_q661 AND symb_decoder(16#1b#)) OR
 					(reg_q661 AND symb_decoder(16#58#)) OR
 					(reg_q661 AND symb_decoder(16#9f#)) OR
 					(reg_q661 AND symb_decoder(16#34#)) OR
 					(reg_q661 AND symb_decoder(16#f0#)) OR
 					(reg_q661 AND symb_decoder(16#c0#)) OR
 					(reg_q661 AND symb_decoder(16#b5#)) OR
 					(reg_q661 AND symb_decoder(16#77#)) OR
 					(reg_q661 AND symb_decoder(16#11#)) OR
 					(reg_q661 AND symb_decoder(16#1d#)) OR
 					(reg_q661 AND symb_decoder(16#59#)) OR
 					(reg_q661 AND symb_decoder(16#cb#)) OR
 					(reg_q661 AND symb_decoder(16#7b#)) OR
 					(reg_q661 AND symb_decoder(16#3a#)) OR
 					(reg_q661 AND symb_decoder(16#d2#)) OR
 					(reg_q661 AND symb_decoder(16#91#)) OR
 					(reg_q661 AND symb_decoder(16#eb#)) OR
 					(reg_q661 AND symb_decoder(16#57#)) OR
 					(reg_q661 AND symb_decoder(16#9b#)) OR
 					(reg_q661 AND symb_decoder(16#ac#)) OR
 					(reg_q661 AND symb_decoder(16#3d#)) OR
 					(reg_q661 AND symb_decoder(16#2b#)) OR
 					(reg_q661 AND symb_decoder(16#24#)) OR
 					(reg_q661 AND symb_decoder(16#80#)) OR
 					(reg_q661 AND symb_decoder(16#45#)) OR
 					(reg_q661 AND symb_decoder(16#82#)) OR
 					(reg_q661 AND symb_decoder(16#bf#)) OR
 					(reg_q661 AND symb_decoder(16#4c#)) OR
 					(reg_q661 AND symb_decoder(16#f6#)) OR
 					(reg_q661 AND symb_decoder(16#6d#)) OR
 					(reg_q661 AND symb_decoder(16#9e#)) OR
 					(reg_q661 AND symb_decoder(16#6f#)) OR
 					(reg_q661 AND symb_decoder(16#78#)) OR
 					(reg_q661 AND symb_decoder(16#a7#)) OR
 					(reg_q661 AND symb_decoder(16#33#)) OR
 					(reg_q661 AND symb_decoder(16#d3#)) OR
 					(reg_q661 AND symb_decoder(16#30#)) OR
 					(reg_q661 AND symb_decoder(16#d0#)) OR
 					(reg_q661 AND symb_decoder(16#50#)) OR
 					(reg_q661 AND symb_decoder(16#94#)) OR
 					(reg_q661 AND symb_decoder(16#f3#)) OR
 					(reg_q661 AND symb_decoder(16#9c#)) OR
 					(reg_q661 AND symb_decoder(16#0e#)) OR
 					(reg_q661 AND symb_decoder(16#63#)) OR
 					(reg_q661 AND symb_decoder(16#44#)) OR
 					(reg_q661 AND symb_decoder(16#8c#)) OR
 					(reg_q661 AND symb_decoder(16#0b#)) OR
 					(reg_q661 AND symb_decoder(16#f5#)) OR
 					(reg_q661 AND symb_decoder(16#19#)) OR
 					(reg_q661 AND symb_decoder(16#5a#)) OR
 					(reg_q661 AND symb_decoder(16#0f#)) OR
 					(reg_q661 AND symb_decoder(16#0a#)) OR
 					(reg_q661 AND symb_decoder(16#60#)) OR
 					(reg_q661 AND symb_decoder(16#af#)) OR
 					(reg_q661 AND symb_decoder(16#71#)) OR
 					(reg_q661 AND symb_decoder(16#e2#)) OR
 					(reg_q661 AND symb_decoder(16#bc#)) OR
 					(reg_q661 AND symb_decoder(16#b6#)) OR
 					(reg_q661 AND symb_decoder(16#c8#)) OR
 					(reg_q661 AND symb_decoder(16#2a#)) OR
 					(reg_q661 AND symb_decoder(16#42#)) OR
 					(reg_q661 AND symb_decoder(16#28#)) OR
 					(reg_q661 AND symb_decoder(16#02#)) OR
 					(reg_q661 AND symb_decoder(16#39#)) OR
 					(reg_q661 AND symb_decoder(16#be#)) OR
 					(reg_q661 AND symb_decoder(16#c2#)) OR
 					(reg_q661 AND symb_decoder(16#ad#)) OR
 					(reg_q661 AND symb_decoder(16#e9#)) OR
 					(reg_q661 AND symb_decoder(16#53#)) OR
 					(reg_q661 AND symb_decoder(16#cd#)) OR
 					(reg_q661 AND symb_decoder(16#f4#)) OR
 					(reg_q661 AND symb_decoder(16#47#)) OR
 					(reg_q661 AND symb_decoder(16#b0#)) OR
 					(reg_q661 AND symb_decoder(16#48#)) OR
 					(reg_q661 AND symb_decoder(16#5c#)) OR
 					(reg_q661 AND symb_decoder(16#08#)) OR
 					(reg_q661 AND symb_decoder(16#bd#)) OR
 					(reg_q661 AND symb_decoder(16#5f#)) OR
 					(reg_q661 AND symb_decoder(16#ca#)) OR
 					(reg_q661 AND symb_decoder(16#e5#)) OR
 					(reg_q661 AND symb_decoder(16#62#)) OR
 					(reg_q661 AND symb_decoder(16#73#)) OR
 					(reg_q661 AND symb_decoder(16#27#)) OR
 					(reg_q661 AND symb_decoder(16#b7#)) OR
 					(reg_q661 AND symb_decoder(16#13#)) OR
 					(reg_q661 AND symb_decoder(16#56#)) OR
 					(reg_q661 AND symb_decoder(16#a9#)) OR
 					(reg_q661 AND symb_decoder(16#a4#)) OR
 					(reg_q661 AND symb_decoder(16#65#)) OR
 					(reg_q661 AND symb_decoder(16#c1#)) OR
 					(reg_q661 AND symb_decoder(16#69#)) OR
 					(reg_q661 AND symb_decoder(16#0c#)) OR
 					(reg_q661 AND symb_decoder(16#00#)) OR
 					(reg_q661 AND symb_decoder(16#aa#)) OR
 					(reg_q661 AND symb_decoder(16#6a#)) OR
 					(reg_q661 AND symb_decoder(16#76#)) OR
 					(reg_q661 AND symb_decoder(16#40#)) OR
 					(reg_q661 AND symb_decoder(16#fe#)) OR
 					(reg_q661 AND symb_decoder(16#41#)) OR
 					(reg_q661 AND symb_decoder(16#22#)) OR
 					(reg_q661 AND symb_decoder(16#f2#)) OR
 					(reg_q661 AND symb_decoder(16#83#)) OR
 					(reg_q661 AND symb_decoder(16#b2#)) OR
 					(reg_q661 AND symb_decoder(16#7a#)) OR
 					(reg_q661 AND symb_decoder(16#ec#)) OR
 					(reg_q661 AND symb_decoder(16#e0#)) OR
 					(reg_q661 AND symb_decoder(16#a6#)) OR
 					(reg_q661 AND symb_decoder(16#cf#)) OR
 					(reg_q661 AND symb_decoder(16#96#)) OR
 					(reg_q661 AND symb_decoder(16#15#)) OR
 					(reg_q661 AND symb_decoder(16#46#)) OR
 					(reg_q661 AND symb_decoder(16#43#)) OR
 					(reg_q661 AND symb_decoder(16#86#)) OR
 					(reg_q661 AND symb_decoder(16#d8#)) OR
 					(reg_q661 AND symb_decoder(16#ba#)) OR
 					(reg_q661 AND symb_decoder(16#64#)) OR
 					(reg_q661 AND symb_decoder(16#db#)) OR
 					(reg_q661 AND symb_decoder(16#85#)) OR
 					(reg_q661 AND symb_decoder(16#b8#)) OR
 					(reg_q661 AND symb_decoder(16#7e#)) OR
 					(reg_q661 AND symb_decoder(16#31#)) OR
 					(reg_q661 AND symb_decoder(16#9d#)) OR
 					(reg_q661 AND symb_decoder(16#6c#)) OR
 					(reg_q661 AND symb_decoder(16#98#)) OR
 					(reg_q661 AND symb_decoder(16#3f#)) OR
 					(reg_q661 AND symb_decoder(16#da#)) OR
 					(reg_q661 AND symb_decoder(16#fc#)) OR
 					(reg_q661 AND symb_decoder(16#8b#)) OR
 					(reg_q661 AND symb_decoder(16#b9#)) OR
 					(reg_q661 AND symb_decoder(16#52#)) OR
 					(reg_q661 AND symb_decoder(16#de#)) OR
 					(reg_q661 AND symb_decoder(16#06#)) OR
 					(reg_q661 AND symb_decoder(16#3e#)) OR
 					(reg_q661 AND symb_decoder(16#6b#)) OR
 					(reg_q661 AND symb_decoder(16#d7#)) OR
 					(reg_q661 AND symb_decoder(16#81#)) OR
 					(reg_q661 AND symb_decoder(16#05#)) OR
 					(reg_q661 AND symb_decoder(16#8d#)) OR
 					(reg_q661 AND symb_decoder(16#9a#)) OR
 					(reg_q661 AND symb_decoder(16#a1#)) OR
 					(reg_q661 AND symb_decoder(16#54#)) OR
 					(reg_q661 AND symb_decoder(16#66#)) OR
 					(reg_q661 AND symb_decoder(16#8f#)) OR
 					(reg_q661 AND symb_decoder(16#f7#)) OR
 					(reg_q661 AND symb_decoder(16#92#)) OR
 					(reg_q661 AND symb_decoder(16#29#)) OR
 					(reg_q661 AND symb_decoder(16#70#)) OR
 					(reg_q661 AND symb_decoder(16#51#)) OR
 					(reg_q661 AND symb_decoder(16#87#)) OR
 					(reg_q661 AND symb_decoder(16#04#)) OR
 					(reg_q661 AND symb_decoder(16#a5#)) OR
 					(reg_q661 AND symb_decoder(16#c3#)) OR
 					(reg_q661 AND symb_decoder(16#03#)) OR
 					(reg_q661 AND symb_decoder(16#36#)) OR
 					(reg_q661 AND symb_decoder(16#f9#)) OR
 					(reg_q661 AND symb_decoder(16#97#)) OR
 					(reg_q661 AND symb_decoder(16#e7#)) OR
 					(reg_q661 AND symb_decoder(16#ee#)) OR
 					(reg_q661 AND symb_decoder(16#d6#));
reg_q661_init <= '0' ;
	p_reg_q661: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q661 <= reg_q661_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q661 <= reg_q661_init;
        else
          reg_q661 <= reg_q661_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2329_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q2329 AND symb_decoder(16#26#)) OR
 					(reg_q2329 AND symb_decoder(16#de#)) OR
 					(reg_q2329 AND symb_decoder(16#2f#)) OR
 					(reg_q2329 AND symb_decoder(16#95#)) OR
 					(reg_q2329 AND symb_decoder(16#66#)) OR
 					(reg_q2329 AND symb_decoder(16#93#)) OR
 					(reg_q2329 AND symb_decoder(16#97#)) OR
 					(reg_q2329 AND symb_decoder(16#d9#)) OR
 					(reg_q2329 AND symb_decoder(16#f3#)) OR
 					(reg_q2329 AND symb_decoder(16#02#)) OR
 					(reg_q2329 AND symb_decoder(16#1d#)) OR
 					(reg_q2329 AND symb_decoder(16#99#)) OR
 					(reg_q2329 AND symb_decoder(16#48#)) OR
 					(reg_q2329 AND symb_decoder(16#8e#)) OR
 					(reg_q2329 AND symb_decoder(16#61#)) OR
 					(reg_q2329 AND symb_decoder(16#ef#)) OR
 					(reg_q2329 AND symb_decoder(16#12#)) OR
 					(reg_q2329 AND symb_decoder(16#5d#)) OR
 					(reg_q2329 AND symb_decoder(16#4d#)) OR
 					(reg_q2329 AND symb_decoder(16#35#)) OR
 					(reg_q2329 AND symb_decoder(16#da#)) OR
 					(reg_q2329 AND symb_decoder(16#1c#)) OR
 					(reg_q2329 AND symb_decoder(16#b7#)) OR
 					(reg_q2329 AND symb_decoder(16#81#)) OR
 					(reg_q2329 AND symb_decoder(16#cc#)) OR
 					(reg_q2329 AND symb_decoder(16#86#)) OR
 					(reg_q2329 AND symb_decoder(16#c3#)) OR
 					(reg_q2329 AND symb_decoder(16#44#)) OR
 					(reg_q2329 AND symb_decoder(16#b5#)) OR
 					(reg_q2329 AND symb_decoder(16#cb#)) OR
 					(reg_q2329 AND symb_decoder(16#34#)) OR
 					(reg_q2329 AND symb_decoder(16#31#)) OR
 					(reg_q2329 AND symb_decoder(16#0a#)) OR
 					(reg_q2329 AND symb_decoder(16#6b#)) OR
 					(reg_q2329 AND symb_decoder(16#32#)) OR
 					(reg_q2329 AND symb_decoder(16#74#)) OR
 					(reg_q2329 AND symb_decoder(16#5c#)) OR
 					(reg_q2329 AND symb_decoder(16#3b#)) OR
 					(reg_q2329 AND symb_decoder(16#dd#)) OR
 					(reg_q2329 AND symb_decoder(16#bd#)) OR
 					(reg_q2329 AND symb_decoder(16#8b#)) OR
 					(reg_q2329 AND symb_decoder(16#c6#)) OR
 					(reg_q2329 AND symb_decoder(16#eb#)) OR
 					(reg_q2329 AND symb_decoder(16#0e#)) OR
 					(reg_q2329 AND symb_decoder(16#aa#)) OR
 					(reg_q2329 AND symb_decoder(16#3d#)) OR
 					(reg_q2329 AND symb_decoder(16#4e#)) OR
 					(reg_q2329 AND symb_decoder(16#d7#)) OR
 					(reg_q2329 AND symb_decoder(16#fb#)) OR
 					(reg_q2329 AND symb_decoder(16#15#)) OR
 					(reg_q2329 AND symb_decoder(16#8f#)) OR
 					(reg_q2329 AND symb_decoder(16#c1#)) OR
 					(reg_q2329 AND symb_decoder(16#6d#)) OR
 					(reg_q2329 AND symb_decoder(16#d5#)) OR
 					(reg_q2329 AND symb_decoder(16#d2#)) OR
 					(reg_q2329 AND symb_decoder(16#00#)) OR
 					(reg_q2329 AND symb_decoder(16#21#)) OR
 					(reg_q2329 AND symb_decoder(16#d0#)) OR
 					(reg_q2329 AND symb_decoder(16#05#)) OR
 					(reg_q2329 AND symb_decoder(16#7a#)) OR
 					(reg_q2329 AND symb_decoder(16#04#)) OR
 					(reg_q2329 AND symb_decoder(16#ae#)) OR
 					(reg_q2329 AND symb_decoder(16#fe#)) OR
 					(reg_q2329 AND symb_decoder(16#01#)) OR
 					(reg_q2329 AND symb_decoder(16#e3#)) OR
 					(reg_q2329 AND symb_decoder(16#58#)) OR
 					(reg_q2329 AND symb_decoder(16#50#)) OR
 					(reg_q2329 AND symb_decoder(16#9d#)) OR
 					(reg_q2329 AND symb_decoder(16#78#)) OR
 					(reg_q2329 AND symb_decoder(16#3a#)) OR
 					(reg_q2329 AND symb_decoder(16#88#)) OR
 					(reg_q2329 AND symb_decoder(16#fd#)) OR
 					(reg_q2329 AND symb_decoder(16#68#)) OR
 					(reg_q2329 AND symb_decoder(16#69#)) OR
 					(reg_q2329 AND symb_decoder(16#0d#)) OR
 					(reg_q2329 AND symb_decoder(16#39#)) OR
 					(reg_q2329 AND symb_decoder(16#30#)) OR
 					(reg_q2329 AND symb_decoder(16#37#)) OR
 					(reg_q2329 AND symb_decoder(16#e6#)) OR
 					(reg_q2329 AND symb_decoder(16#2b#)) OR
 					(reg_q2329 AND symb_decoder(16#27#)) OR
 					(reg_q2329 AND symb_decoder(16#ca#)) OR
 					(reg_q2329 AND symb_decoder(16#07#)) OR
 					(reg_q2329 AND symb_decoder(16#e8#)) OR
 					(reg_q2329 AND symb_decoder(16#b8#)) OR
 					(reg_q2329 AND symb_decoder(16#51#)) OR
 					(reg_q2329 AND symb_decoder(16#73#)) OR
 					(reg_q2329 AND symb_decoder(16#a1#)) OR
 					(reg_q2329 AND symb_decoder(16#d1#)) OR
 					(reg_q2329 AND symb_decoder(16#fc#)) OR
 					(reg_q2329 AND symb_decoder(16#d4#)) OR
 					(reg_q2329 AND symb_decoder(16#38#)) OR
 					(reg_q2329 AND symb_decoder(16#03#)) OR
 					(reg_q2329 AND symb_decoder(16#ea#)) OR
 					(reg_q2329 AND symb_decoder(16#f0#)) OR
 					(reg_q2329 AND symb_decoder(16#c0#)) OR
 					(reg_q2329 AND symb_decoder(16#c9#)) OR
 					(reg_q2329 AND symb_decoder(16#b3#)) OR
 					(reg_q2329 AND symb_decoder(16#d8#)) OR
 					(reg_q2329 AND symb_decoder(16#bc#)) OR
 					(reg_q2329 AND symb_decoder(16#fa#)) OR
 					(reg_q2329 AND symb_decoder(16#70#)) OR
 					(reg_q2329 AND symb_decoder(16#b2#)) OR
 					(reg_q2329 AND symb_decoder(16#90#)) OR
 					(reg_q2329 AND symb_decoder(16#7c#)) OR
 					(reg_q2329 AND symb_decoder(16#e5#)) OR
 					(reg_q2329 AND symb_decoder(16#6e#)) OR
 					(reg_q2329 AND symb_decoder(16#cf#)) OR
 					(reg_q2329 AND symb_decoder(16#0c#)) OR
 					(reg_q2329 AND symb_decoder(16#45#)) OR
 					(reg_q2329 AND symb_decoder(16#57#)) OR
 					(reg_q2329 AND symb_decoder(16#ce#)) OR
 					(reg_q2329 AND symb_decoder(16#29#)) OR
 					(reg_q2329 AND symb_decoder(16#a2#)) OR
 					(reg_q2329 AND symb_decoder(16#f9#)) OR
 					(reg_q2329 AND symb_decoder(16#4b#)) OR
 					(reg_q2329 AND symb_decoder(16#65#)) OR
 					(reg_q2329 AND symb_decoder(16#bf#)) OR
 					(reg_q2329 AND symb_decoder(16#14#)) OR
 					(reg_q2329 AND symb_decoder(16#77#)) OR
 					(reg_q2329 AND symb_decoder(16#83#)) OR
 					(reg_q2329 AND symb_decoder(16#17#)) OR
 					(reg_q2329 AND symb_decoder(16#4f#)) OR
 					(reg_q2329 AND symb_decoder(16#84#)) OR
 					(reg_q2329 AND symb_decoder(16#f2#)) OR
 					(reg_q2329 AND symb_decoder(16#56#)) OR
 					(reg_q2329 AND symb_decoder(16#94#)) OR
 					(reg_q2329 AND symb_decoder(16#6a#)) OR
 					(reg_q2329 AND symb_decoder(16#7b#)) OR
 					(reg_q2329 AND symb_decoder(16#d6#)) OR
 					(reg_q2329 AND symb_decoder(16#c2#)) OR
 					(reg_q2329 AND symb_decoder(16#60#)) OR
 					(reg_q2329 AND symb_decoder(16#20#)) OR
 					(reg_q2329 AND symb_decoder(16#0b#)) OR
 					(reg_q2329 AND symb_decoder(16#b0#)) OR
 					(reg_q2329 AND symb_decoder(16#91#)) OR
 					(reg_q2329 AND symb_decoder(16#f5#)) OR
 					(reg_q2329 AND symb_decoder(16#5f#)) OR
 					(reg_q2329 AND symb_decoder(16#b4#)) OR
 					(reg_q2329 AND symb_decoder(16#62#)) OR
 					(reg_q2329 AND symb_decoder(16#5a#)) OR
 					(reg_q2329 AND symb_decoder(16#c4#)) OR
 					(reg_q2329 AND symb_decoder(16#75#)) OR
 					(reg_q2329 AND symb_decoder(16#4a#)) OR
 					(reg_q2329 AND symb_decoder(16#af#)) OR
 					(reg_q2329 AND symb_decoder(16#72#)) OR
 					(reg_q2329 AND symb_decoder(16#98#)) OR
 					(reg_q2329 AND symb_decoder(16#b1#)) OR
 					(reg_q2329 AND symb_decoder(16#ad#)) OR
 					(reg_q2329 AND symb_decoder(16#23#)) OR
 					(reg_q2329 AND symb_decoder(16#1a#)) OR
 					(reg_q2329 AND symb_decoder(16#dc#)) OR
 					(reg_q2329 AND symb_decoder(16#a7#)) OR
 					(reg_q2329 AND symb_decoder(16#ed#)) OR
 					(reg_q2329 AND symb_decoder(16#be#)) OR
 					(reg_q2329 AND symb_decoder(16#85#)) OR
 					(reg_q2329 AND symb_decoder(16#9b#)) OR
 					(reg_q2329 AND symb_decoder(16#ee#)) OR
 					(reg_q2329 AND symb_decoder(16#a9#)) OR
 					(reg_q2329 AND symb_decoder(16#40#)) OR
 					(reg_q2329 AND symb_decoder(16#7e#)) OR
 					(reg_q2329 AND symb_decoder(16#87#)) OR
 					(reg_q2329 AND symb_decoder(16#e7#)) OR
 					(reg_q2329 AND symb_decoder(16#10#)) OR
 					(reg_q2329 AND symb_decoder(16#e0#)) OR
 					(reg_q2329 AND symb_decoder(16#ac#)) OR
 					(reg_q2329 AND symb_decoder(16#1e#)) OR
 					(reg_q2329 AND symb_decoder(16#6f#)) OR
 					(reg_q2329 AND symb_decoder(16#52#)) OR
 					(reg_q2329 AND symb_decoder(16#ba#)) OR
 					(reg_q2329 AND symb_decoder(16#1f#)) OR
 					(reg_q2329 AND symb_decoder(16#a6#)) OR
 					(reg_q2329 AND symb_decoder(16#55#)) OR
 					(reg_q2329 AND symb_decoder(16#3e#)) OR
 					(reg_q2329 AND symb_decoder(16#79#)) OR
 					(reg_q2329 AND symb_decoder(16#53#)) OR
 					(reg_q2329 AND symb_decoder(16#3f#)) OR
 					(reg_q2329 AND symb_decoder(16#92#)) OR
 					(reg_q2329 AND symb_decoder(16#59#)) OR
 					(reg_q2329 AND symb_decoder(16#4c#)) OR
 					(reg_q2329 AND symb_decoder(16#71#)) OR
 					(reg_q2329 AND symb_decoder(16#f7#)) OR
 					(reg_q2329 AND symb_decoder(16#6c#)) OR
 					(reg_q2329 AND symb_decoder(16#54#)) OR
 					(reg_q2329 AND symb_decoder(16#43#)) OR
 					(reg_q2329 AND symb_decoder(16#ff#)) OR
 					(reg_q2329 AND symb_decoder(16#a3#)) OR
 					(reg_q2329 AND symb_decoder(16#e4#)) OR
 					(reg_q2329 AND symb_decoder(16#22#)) OR
 					(reg_q2329 AND symb_decoder(16#1b#)) OR
 					(reg_q2329 AND symb_decoder(16#ec#)) OR
 					(reg_q2329 AND symb_decoder(16#09#)) OR
 					(reg_q2329 AND symb_decoder(16#80#)) OR
 					(reg_q2329 AND symb_decoder(16#c8#)) OR
 					(reg_q2329 AND symb_decoder(16#47#)) OR
 					(reg_q2329 AND symb_decoder(16#46#)) OR
 					(reg_q2329 AND symb_decoder(16#9a#)) OR
 					(reg_q2329 AND symb_decoder(16#24#)) OR
 					(reg_q2329 AND symb_decoder(16#a8#)) OR
 					(reg_q2329 AND symb_decoder(16#b9#)) OR
 					(reg_q2329 AND symb_decoder(16#19#)) OR
 					(reg_q2329 AND symb_decoder(16#7f#)) OR
 					(reg_q2329 AND symb_decoder(16#9e#)) OR
 					(reg_q2329 AND symb_decoder(16#8c#)) OR
 					(reg_q2329 AND symb_decoder(16#2e#)) OR
 					(reg_q2329 AND symb_decoder(16#f4#)) OR
 					(reg_q2329 AND symb_decoder(16#67#)) OR
 					(reg_q2329 AND symb_decoder(16#33#)) OR
 					(reg_q2329 AND symb_decoder(16#d3#)) OR
 					(reg_q2329 AND symb_decoder(16#16#)) OR
 					(reg_q2329 AND symb_decoder(16#64#)) OR
 					(reg_q2329 AND symb_decoder(16#b6#)) OR
 					(reg_q2329 AND symb_decoder(16#c7#)) OR
 					(reg_q2329 AND symb_decoder(16#e9#)) OR
 					(reg_q2329 AND symb_decoder(16#bb#)) OR
 					(reg_q2329 AND symb_decoder(16#cd#)) OR
 					(reg_q2329 AND symb_decoder(16#25#)) OR
 					(reg_q2329 AND symb_decoder(16#df#)) OR
 					(reg_q2329 AND symb_decoder(16#a0#)) OR
 					(reg_q2329 AND symb_decoder(16#96#)) OR
 					(reg_q2329 AND symb_decoder(16#49#)) OR
 					(reg_q2329 AND symb_decoder(16#28#)) OR
 					(reg_q2329 AND symb_decoder(16#18#)) OR
 					(reg_q2329 AND symb_decoder(16#63#)) OR
 					(reg_q2329 AND symb_decoder(16#a4#)) OR
 					(reg_q2329 AND symb_decoder(16#db#)) OR
 					(reg_q2329 AND symb_decoder(16#42#)) OR
 					(reg_q2329 AND symb_decoder(16#9f#)) OR
 					(reg_q2329 AND symb_decoder(16#5b#)) OR
 					(reg_q2329 AND symb_decoder(16#a5#)) OR
 					(reg_q2329 AND symb_decoder(16#2d#)) OR
 					(reg_q2329 AND symb_decoder(16#2a#)) OR
 					(reg_q2329 AND symb_decoder(16#89#)) OR
 					(reg_q2329 AND symb_decoder(16#7d#)) OR
 					(reg_q2329 AND symb_decoder(16#c5#)) OR
 					(reg_q2329 AND symb_decoder(16#f8#)) OR
 					(reg_q2329 AND symb_decoder(16#41#)) OR
 					(reg_q2329 AND symb_decoder(16#11#)) OR
 					(reg_q2329 AND symb_decoder(16#82#)) OR
 					(reg_q2329 AND symb_decoder(16#36#)) OR
 					(reg_q2329 AND symb_decoder(16#f6#)) OR
 					(reg_q2329 AND symb_decoder(16#ab#)) OR
 					(reg_q2329 AND symb_decoder(16#08#)) OR
 					(reg_q2329 AND symb_decoder(16#e2#)) OR
 					(reg_q2329 AND symb_decoder(16#9c#)) OR
 					(reg_q2329 AND symb_decoder(16#06#)) OR
 					(reg_q2329 AND symb_decoder(16#e1#)) OR
 					(reg_q2329 AND symb_decoder(16#2c#)) OR
 					(reg_q2329 AND symb_decoder(16#0f#)) OR
 					(reg_q2329 AND symb_decoder(16#13#)) OR
 					(reg_q2329 AND symb_decoder(16#3c#)) OR
 					(reg_q2329 AND symb_decoder(16#f1#)) OR
 					(reg_q2329 AND symb_decoder(16#76#)) OR
 					(reg_q2329 AND symb_decoder(16#5e#)) OR
 					(reg_q2329 AND symb_decoder(16#8d#)) OR
 					(reg_q2329 AND symb_decoder(16#8a#));
reg_q2329_init <= '0' ;
	p_reg_q2329: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2329 <= reg_q2329_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2329 <= reg_q2329_init;
        else
          reg_q2329 <= reg_q2329_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q803_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q803 AND symb_decoder(16#2b#)) OR
 					(reg_q803 AND symb_decoder(16#52#)) OR
 					(reg_q803 AND symb_decoder(16#12#)) OR
 					(reg_q803 AND symb_decoder(16#0f#)) OR
 					(reg_q803 AND symb_decoder(16#64#)) OR
 					(reg_q803 AND symb_decoder(16#6a#)) OR
 					(reg_q803 AND symb_decoder(16#c9#)) OR
 					(reg_q803 AND symb_decoder(16#51#)) OR
 					(reg_q803 AND symb_decoder(16#5a#)) OR
 					(reg_q803 AND symb_decoder(16#a9#)) OR
 					(reg_q803 AND symb_decoder(16#83#)) OR
 					(reg_q803 AND symb_decoder(16#2a#)) OR
 					(reg_q803 AND symb_decoder(16#de#)) OR
 					(reg_q803 AND symb_decoder(16#fe#)) OR
 					(reg_q803 AND symb_decoder(16#af#)) OR
 					(reg_q803 AND symb_decoder(16#d3#)) OR
 					(reg_q803 AND symb_decoder(16#3a#)) OR
 					(reg_q803 AND symb_decoder(16#97#)) OR
 					(reg_q803 AND symb_decoder(16#10#)) OR
 					(reg_q803 AND symb_decoder(16#9f#)) OR
 					(reg_q803 AND symb_decoder(16#c8#)) OR
 					(reg_q803 AND symb_decoder(16#b1#)) OR
 					(reg_q803 AND symb_decoder(16#e3#)) OR
 					(reg_q803 AND symb_decoder(16#24#)) OR
 					(reg_q803 AND symb_decoder(16#75#)) OR
 					(reg_q803 AND symb_decoder(16#8f#)) OR
 					(reg_q803 AND symb_decoder(16#50#)) OR
 					(reg_q803 AND symb_decoder(16#fc#)) OR
 					(reg_q803 AND symb_decoder(16#dc#)) OR
 					(reg_q803 AND symb_decoder(16#b4#)) OR
 					(reg_q803 AND symb_decoder(16#57#)) OR
 					(reg_q803 AND symb_decoder(16#77#)) OR
 					(reg_q803 AND symb_decoder(16#6e#)) OR
 					(reg_q803 AND symb_decoder(16#4c#)) OR
 					(reg_q803 AND symb_decoder(16#cc#)) OR
 					(reg_q803 AND symb_decoder(16#cd#)) OR
 					(reg_q803 AND symb_decoder(16#15#)) OR
 					(reg_q803 AND symb_decoder(16#46#)) OR
 					(reg_q803 AND symb_decoder(16#5f#)) OR
 					(reg_q803 AND symb_decoder(16#5b#)) OR
 					(reg_q803 AND symb_decoder(16#45#)) OR
 					(reg_q803 AND symb_decoder(16#d2#)) OR
 					(reg_q803 AND symb_decoder(16#05#)) OR
 					(reg_q803 AND symb_decoder(16#bf#)) OR
 					(reg_q803 AND symb_decoder(16#d5#)) OR
 					(reg_q803 AND symb_decoder(16#ba#)) OR
 					(reg_q803 AND symb_decoder(16#b7#)) OR
 					(reg_q803 AND symb_decoder(16#ce#)) OR
 					(reg_q803 AND symb_decoder(16#f4#)) OR
 					(reg_q803 AND symb_decoder(16#e5#)) OR
 					(reg_q803 AND symb_decoder(16#7f#)) OR
 					(reg_q803 AND symb_decoder(16#42#)) OR
 					(reg_q803 AND symb_decoder(16#95#)) OR
 					(reg_q803 AND symb_decoder(16#78#)) OR
 					(reg_q803 AND symb_decoder(16#4f#)) OR
 					(reg_q803 AND symb_decoder(16#06#)) OR
 					(reg_q803 AND symb_decoder(16#58#)) OR
 					(reg_q803 AND symb_decoder(16#da#)) OR
 					(reg_q803 AND symb_decoder(16#cb#)) OR
 					(reg_q803 AND symb_decoder(16#be#)) OR
 					(reg_q803 AND symb_decoder(16#0e#)) OR
 					(reg_q803 AND symb_decoder(16#9e#)) OR
 					(reg_q803 AND symb_decoder(16#61#)) OR
 					(reg_q803 AND symb_decoder(16#6b#)) OR
 					(reg_q803 AND symb_decoder(16#37#)) OR
 					(reg_q803 AND symb_decoder(16#ea#)) OR
 					(reg_q803 AND symb_decoder(16#84#)) OR
 					(reg_q803 AND symb_decoder(16#16#)) OR
 					(reg_q803 AND symb_decoder(16#65#)) OR
 					(reg_q803 AND symb_decoder(16#19#)) OR
 					(reg_q803 AND symb_decoder(16#c6#)) OR
 					(reg_q803 AND symb_decoder(16#99#)) OR
 					(reg_q803 AND symb_decoder(16#67#)) OR
 					(reg_q803 AND symb_decoder(16#f7#)) OR
 					(reg_q803 AND symb_decoder(16#30#)) OR
 					(reg_q803 AND symb_decoder(16#c2#)) OR
 					(reg_q803 AND symb_decoder(16#76#)) OR
 					(reg_q803 AND symb_decoder(16#6c#)) OR
 					(reg_q803 AND symb_decoder(16#f0#)) OR
 					(reg_q803 AND symb_decoder(16#d9#)) OR
 					(reg_q803 AND symb_decoder(16#55#)) OR
 					(reg_q803 AND symb_decoder(16#f8#)) OR
 					(reg_q803 AND symb_decoder(16#8e#)) OR
 					(reg_q803 AND symb_decoder(16#d8#)) OR
 					(reg_q803 AND symb_decoder(16#13#)) OR
 					(reg_q803 AND symb_decoder(16#27#)) OR
 					(reg_q803 AND symb_decoder(16#41#)) OR
 					(reg_q803 AND symb_decoder(16#5e#)) OR
 					(reg_q803 AND symb_decoder(16#0c#)) OR
 					(reg_q803 AND symb_decoder(16#3c#)) OR
 					(reg_q803 AND symb_decoder(16#90#)) OR
 					(reg_q803 AND symb_decoder(16#e2#)) OR
 					(reg_q803 AND symb_decoder(16#40#)) OR
 					(reg_q803 AND symb_decoder(16#54#)) OR
 					(reg_q803 AND symb_decoder(16#89#)) OR
 					(reg_q803 AND symb_decoder(16#7c#)) OR
 					(reg_q803 AND symb_decoder(16#ae#)) OR
 					(reg_q803 AND symb_decoder(16#38#)) OR
 					(reg_q803 AND symb_decoder(16#d4#)) OR
 					(reg_q803 AND symb_decoder(16#a5#)) OR
 					(reg_q803 AND symb_decoder(16#fd#)) OR
 					(reg_q803 AND symb_decoder(16#8c#)) OR
 					(reg_q803 AND symb_decoder(16#ca#)) OR
 					(reg_q803 AND symb_decoder(16#b5#)) OR
 					(reg_q803 AND symb_decoder(16#e0#)) OR
 					(reg_q803 AND symb_decoder(16#0a#)) OR
 					(reg_q803 AND symb_decoder(16#a3#)) OR
 					(reg_q803 AND symb_decoder(16#2c#)) OR
 					(reg_q803 AND symb_decoder(16#21#)) OR
 					(reg_q803 AND symb_decoder(16#88#)) OR
 					(reg_q803 AND symb_decoder(16#bd#)) OR
 					(reg_q803 AND symb_decoder(16#9b#)) OR
 					(reg_q803 AND symb_decoder(16#81#)) OR
 					(reg_q803 AND symb_decoder(16#d0#)) OR
 					(reg_q803 AND symb_decoder(16#18#)) OR
 					(reg_q803 AND symb_decoder(16#aa#)) OR
 					(reg_q803 AND symb_decoder(16#b3#)) OR
 					(reg_q803 AND symb_decoder(16#b2#)) OR
 					(reg_q803 AND symb_decoder(16#4b#)) OR
 					(reg_q803 AND symb_decoder(16#e8#)) OR
 					(reg_q803 AND symb_decoder(16#4e#)) OR
 					(reg_q803 AND symb_decoder(16#07#)) OR
 					(reg_q803 AND symb_decoder(16#dd#)) OR
 					(reg_q803 AND symb_decoder(16#f9#)) OR
 					(reg_q803 AND symb_decoder(16#3e#)) OR
 					(reg_q803 AND symb_decoder(16#a7#)) OR
 					(reg_q803 AND symb_decoder(16#11#)) OR
 					(reg_q803 AND symb_decoder(16#8d#)) OR
 					(reg_q803 AND symb_decoder(16#7a#)) OR
 					(reg_q803 AND symb_decoder(16#b6#)) OR
 					(reg_q803 AND symb_decoder(16#49#)) OR
 					(reg_q803 AND symb_decoder(16#33#)) OR
 					(reg_q803 AND symb_decoder(16#00#)) OR
 					(reg_q803 AND symb_decoder(16#92#)) OR
 					(reg_q803 AND symb_decoder(16#bc#)) OR
 					(reg_q803 AND symb_decoder(16#1f#)) OR
 					(reg_q803 AND symb_decoder(16#0b#)) OR
 					(reg_q803 AND symb_decoder(16#29#)) OR
 					(reg_q803 AND symb_decoder(16#14#)) OR
 					(reg_q803 AND symb_decoder(16#db#)) OR
 					(reg_q803 AND symb_decoder(16#70#)) OR
 					(reg_q803 AND symb_decoder(16#f2#)) OR
 					(reg_q803 AND symb_decoder(16#62#)) OR
 					(reg_q803 AND symb_decoder(16#0d#)) OR
 					(reg_q803 AND symb_decoder(16#36#)) OR
 					(reg_q803 AND symb_decoder(16#c4#)) OR
 					(reg_q803 AND symb_decoder(16#35#)) OR
 					(reg_q803 AND symb_decoder(16#31#)) OR
 					(reg_q803 AND symb_decoder(16#a1#)) OR
 					(reg_q803 AND symb_decoder(16#2f#)) OR
 					(reg_q803 AND symb_decoder(16#f6#)) OR
 					(reg_q803 AND symb_decoder(16#b8#)) OR
 					(reg_q803 AND symb_decoder(16#e1#)) OR
 					(reg_q803 AND symb_decoder(16#e7#)) OR
 					(reg_q803 AND symb_decoder(16#ad#)) OR
 					(reg_q803 AND symb_decoder(16#c5#)) OR
 					(reg_q803 AND symb_decoder(16#b9#)) OR
 					(reg_q803 AND symb_decoder(16#8b#)) OR
 					(reg_q803 AND symb_decoder(16#1a#)) OR
 					(reg_q803 AND symb_decoder(16#48#)) OR
 					(reg_q803 AND symb_decoder(16#28#)) OR
 					(reg_q803 AND symb_decoder(16#96#)) OR
 					(reg_q803 AND symb_decoder(16#c0#)) OR
 					(reg_q803 AND symb_decoder(16#a2#)) OR
 					(reg_q803 AND symb_decoder(16#1c#)) OR
 					(reg_q803 AND symb_decoder(16#9d#)) OR
 					(reg_q803 AND symb_decoder(16#d1#)) OR
 					(reg_q803 AND symb_decoder(16#c3#)) OR
 					(reg_q803 AND symb_decoder(16#a0#)) OR
 					(reg_q803 AND symb_decoder(16#68#)) OR
 					(reg_q803 AND symb_decoder(16#df#)) OR
 					(reg_q803 AND symb_decoder(16#1d#)) OR
 					(reg_q803 AND symb_decoder(16#53#)) OR
 					(reg_q803 AND symb_decoder(16#26#)) OR
 					(reg_q803 AND symb_decoder(16#93#)) OR
 					(reg_q803 AND symb_decoder(16#94#)) OR
 					(reg_q803 AND symb_decoder(16#e9#)) OR
 					(reg_q803 AND symb_decoder(16#c1#)) OR
 					(reg_q803 AND symb_decoder(16#ef#)) OR
 					(reg_q803 AND symb_decoder(16#32#)) OR
 					(reg_q803 AND symb_decoder(16#22#)) OR
 					(reg_q803 AND symb_decoder(16#1e#)) OR
 					(reg_q803 AND symb_decoder(16#e4#)) OR
 					(reg_q803 AND symb_decoder(16#7b#)) OR
 					(reg_q803 AND symb_decoder(16#9a#)) OR
 					(reg_q803 AND symb_decoder(16#cf#)) OR
 					(reg_q803 AND symb_decoder(16#d6#)) OR
 					(reg_q803 AND symb_decoder(16#91#)) OR
 					(reg_q803 AND symb_decoder(16#01#)) OR
 					(reg_q803 AND symb_decoder(16#eb#)) OR
 					(reg_q803 AND symb_decoder(16#63#)) OR
 					(reg_q803 AND symb_decoder(16#6f#)) OR
 					(reg_q803 AND symb_decoder(16#6d#)) OR
 					(reg_q803 AND symb_decoder(16#66#)) OR
 					(reg_q803 AND symb_decoder(16#7d#)) OR
 					(reg_q803 AND symb_decoder(16#d7#)) OR
 					(reg_q803 AND symb_decoder(16#4d#)) OR
 					(reg_q803 AND symb_decoder(16#86#)) OR
 					(reg_q803 AND symb_decoder(16#bb#)) OR
 					(reg_q803 AND symb_decoder(16#ec#)) OR
 					(reg_q803 AND symb_decoder(16#5d#)) OR
 					(reg_q803 AND symb_decoder(16#1b#)) OR
 					(reg_q803 AND symb_decoder(16#72#)) OR
 					(reg_q803 AND symb_decoder(16#ee#)) OR
 					(reg_q803 AND symb_decoder(16#74#)) OR
 					(reg_q803 AND symb_decoder(16#56#)) OR
 					(reg_q803 AND symb_decoder(16#87#)) OR
 					(reg_q803 AND symb_decoder(16#39#)) OR
 					(reg_q803 AND symb_decoder(16#47#)) OR
 					(reg_q803 AND symb_decoder(16#4a#)) OR
 					(reg_q803 AND symb_decoder(16#3b#)) OR
 					(reg_q803 AND symb_decoder(16#08#)) OR
 					(reg_q803 AND symb_decoder(16#9c#)) OR
 					(reg_q803 AND symb_decoder(16#02#)) OR
 					(reg_q803 AND symb_decoder(16#ac#)) OR
 					(reg_q803 AND symb_decoder(16#98#)) OR
 					(reg_q803 AND symb_decoder(16#43#)) OR
 					(reg_q803 AND symb_decoder(16#2e#)) OR
 					(reg_q803 AND symb_decoder(16#b0#)) OR
 					(reg_q803 AND symb_decoder(16#5c#)) OR
 					(reg_q803 AND symb_decoder(16#04#)) OR
 					(reg_q803 AND symb_decoder(16#73#)) OR
 					(reg_q803 AND symb_decoder(16#59#)) OR
 					(reg_q803 AND symb_decoder(16#25#)) OR
 					(reg_q803 AND symb_decoder(16#2d#)) OR
 					(reg_q803 AND symb_decoder(16#34#)) OR
 					(reg_q803 AND symb_decoder(16#e6#)) OR
 					(reg_q803 AND symb_decoder(16#80#)) OR
 					(reg_q803 AND symb_decoder(16#ff#)) OR
 					(reg_q803 AND symb_decoder(16#fb#)) OR
 					(reg_q803 AND symb_decoder(16#f1#)) OR
 					(reg_q803 AND symb_decoder(16#f5#)) OR
 					(reg_q803 AND symb_decoder(16#79#)) OR
 					(reg_q803 AND symb_decoder(16#3f#)) OR
 					(reg_q803 AND symb_decoder(16#03#)) OR
 					(reg_q803 AND symb_decoder(16#a6#)) OR
 					(reg_q803 AND symb_decoder(16#f3#)) OR
 					(reg_q803 AND symb_decoder(16#20#)) OR
 					(reg_q803 AND symb_decoder(16#17#)) OR
 					(reg_q803 AND symb_decoder(16#69#)) OR
 					(reg_q803 AND symb_decoder(16#a4#)) OR
 					(reg_q803 AND symb_decoder(16#fa#)) OR
 					(reg_q803 AND symb_decoder(16#ed#)) OR
 					(reg_q803 AND symb_decoder(16#7e#)) OR
 					(reg_q803 AND symb_decoder(16#3d#)) OR
 					(reg_q803 AND symb_decoder(16#85#)) OR
 					(reg_q803 AND symb_decoder(16#ab#)) OR
 					(reg_q803 AND symb_decoder(16#44#)) OR
 					(reg_q803 AND symb_decoder(16#c7#)) OR
 					(reg_q803 AND symb_decoder(16#8a#)) OR
 					(reg_q803 AND symb_decoder(16#23#)) OR
 					(reg_q803 AND symb_decoder(16#09#)) OR
 					(reg_q803 AND symb_decoder(16#a8#)) OR
 					(reg_q803 AND symb_decoder(16#82#)) OR
 					(reg_q803 AND symb_decoder(16#60#)) OR
 					(reg_q803 AND symb_decoder(16#71#));
reg_q803_init <= '0' ;
	p_reg_q803: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q803 <= reg_q803_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q803 <= reg_q803_init;
        else
          reg_q803 <= reg_q803_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q604_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q604 AND symb_decoder(16#09#)) OR
 					(reg_q604 AND symb_decoder(16#d1#)) OR
 					(reg_q604 AND symb_decoder(16#2d#)) OR
 					(reg_q604 AND symb_decoder(16#d6#)) OR
 					(reg_q604 AND symb_decoder(16#b6#)) OR
 					(reg_q604 AND symb_decoder(16#9f#)) OR
 					(reg_q604 AND symb_decoder(16#1a#)) OR
 					(reg_q604 AND symb_decoder(16#d7#)) OR
 					(reg_q604 AND symb_decoder(16#c8#)) OR
 					(reg_q604 AND symb_decoder(16#ba#)) OR
 					(reg_q604 AND symb_decoder(16#34#)) OR
 					(reg_q604 AND symb_decoder(16#f9#)) OR
 					(reg_q604 AND symb_decoder(16#22#)) OR
 					(reg_q604 AND symb_decoder(16#f3#)) OR
 					(reg_q604 AND symb_decoder(16#6e#)) OR
 					(reg_q604 AND symb_decoder(16#4c#)) OR
 					(reg_q604 AND symb_decoder(16#d9#)) OR
 					(reg_q604 AND symb_decoder(16#df#)) OR
 					(reg_q604 AND symb_decoder(16#0a#)) OR
 					(reg_q604 AND symb_decoder(16#04#)) OR
 					(reg_q604 AND symb_decoder(16#00#)) OR
 					(reg_q604 AND symb_decoder(16#bf#)) OR
 					(reg_q604 AND symb_decoder(16#6b#)) OR
 					(reg_q604 AND symb_decoder(16#ef#)) OR
 					(reg_q604 AND symb_decoder(16#d4#)) OR
 					(reg_q604 AND symb_decoder(16#bc#)) OR
 					(reg_q604 AND symb_decoder(16#37#)) OR
 					(reg_q604 AND symb_decoder(16#7a#)) OR
 					(reg_q604 AND symb_decoder(16#3f#)) OR
 					(reg_q604 AND symb_decoder(16#69#)) OR
 					(reg_q604 AND symb_decoder(16#f0#)) OR
 					(reg_q604 AND symb_decoder(16#bd#)) OR
 					(reg_q604 AND symb_decoder(16#a2#)) OR
 					(reg_q604 AND symb_decoder(16#91#)) OR
 					(reg_q604 AND symb_decoder(16#a0#)) OR
 					(reg_q604 AND symb_decoder(16#74#)) OR
 					(reg_q604 AND symb_decoder(16#c2#)) OR
 					(reg_q604 AND symb_decoder(16#3e#)) OR
 					(reg_q604 AND symb_decoder(16#da#)) OR
 					(reg_q604 AND symb_decoder(16#c6#)) OR
 					(reg_q604 AND symb_decoder(16#25#)) OR
 					(reg_q604 AND symb_decoder(16#7e#)) OR
 					(reg_q604 AND symb_decoder(16#11#)) OR
 					(reg_q604 AND symb_decoder(16#1c#)) OR
 					(reg_q604 AND symb_decoder(16#56#)) OR
 					(reg_q604 AND symb_decoder(16#39#)) OR
 					(reg_q604 AND symb_decoder(16#b7#)) OR
 					(reg_q604 AND symb_decoder(16#13#)) OR
 					(reg_q604 AND symb_decoder(16#28#)) OR
 					(reg_q604 AND symb_decoder(16#ec#)) OR
 					(reg_q604 AND symb_decoder(16#0e#)) OR
 					(reg_q604 AND symb_decoder(16#1b#)) OR
 					(reg_q604 AND symb_decoder(16#e8#)) OR
 					(reg_q604 AND symb_decoder(16#87#)) OR
 					(reg_q604 AND symb_decoder(16#8c#)) OR
 					(reg_q604 AND symb_decoder(16#e4#)) OR
 					(reg_q604 AND symb_decoder(16#40#)) OR
 					(reg_q604 AND symb_decoder(16#a9#)) OR
 					(reg_q604 AND symb_decoder(16#21#)) OR
 					(reg_q604 AND symb_decoder(16#a5#)) OR
 					(reg_q604 AND symb_decoder(16#71#)) OR
 					(reg_q604 AND symb_decoder(16#b4#)) OR
 					(reg_q604 AND symb_decoder(16#65#)) OR
 					(reg_q604 AND symb_decoder(16#3d#)) OR
 					(reg_q604 AND symb_decoder(16#14#)) OR
 					(reg_q604 AND symb_decoder(16#31#)) OR
 					(reg_q604 AND symb_decoder(16#2c#)) OR
 					(reg_q604 AND symb_decoder(16#26#)) OR
 					(reg_q604 AND symb_decoder(16#b1#)) OR
 					(reg_q604 AND symb_decoder(16#73#)) OR
 					(reg_q604 AND symb_decoder(16#ac#)) OR
 					(reg_q604 AND symb_decoder(16#67#)) OR
 					(reg_q604 AND symb_decoder(16#17#)) OR
 					(reg_q604 AND symb_decoder(16#0b#)) OR
 					(reg_q604 AND symb_decoder(16#0c#)) OR
 					(reg_q604 AND symb_decoder(16#98#)) OR
 					(reg_q604 AND symb_decoder(16#a6#)) OR
 					(reg_q604 AND symb_decoder(16#96#)) OR
 					(reg_q604 AND symb_decoder(16#f4#)) OR
 					(reg_q604 AND symb_decoder(16#77#)) OR
 					(reg_q604 AND symb_decoder(16#05#)) OR
 					(reg_q604 AND symb_decoder(16#4e#)) OR
 					(reg_q604 AND symb_decoder(16#9b#)) OR
 					(reg_q604 AND symb_decoder(16#19#)) OR
 					(reg_q604 AND symb_decoder(16#a4#)) OR
 					(reg_q604 AND symb_decoder(16#53#)) OR
 					(reg_q604 AND symb_decoder(16#e6#)) OR
 					(reg_q604 AND symb_decoder(16#de#)) OR
 					(reg_q604 AND symb_decoder(16#be#)) OR
 					(reg_q604 AND symb_decoder(16#ed#)) OR
 					(reg_q604 AND symb_decoder(16#5d#)) OR
 					(reg_q604 AND symb_decoder(16#aa#)) OR
 					(reg_q604 AND symb_decoder(16#e9#)) OR
 					(reg_q604 AND symb_decoder(16#a1#)) OR
 					(reg_q604 AND symb_decoder(16#8d#)) OR
 					(reg_q604 AND symb_decoder(16#6f#)) OR
 					(reg_q604 AND symb_decoder(16#e1#)) OR
 					(reg_q604 AND symb_decoder(16#7b#)) OR
 					(reg_q604 AND symb_decoder(16#4b#)) OR
 					(reg_q604 AND symb_decoder(16#15#)) OR
 					(reg_q604 AND symb_decoder(16#82#)) OR
 					(reg_q604 AND symb_decoder(16#cf#)) OR
 					(reg_q604 AND symb_decoder(16#ff#)) OR
 					(reg_q604 AND symb_decoder(16#eb#)) OR
 					(reg_q604 AND symb_decoder(16#fa#)) OR
 					(reg_q604 AND symb_decoder(16#78#)) OR
 					(reg_q604 AND symb_decoder(16#42#)) OR
 					(reg_q604 AND symb_decoder(16#4f#)) OR
 					(reg_q604 AND symb_decoder(16#db#)) OR
 					(reg_q604 AND symb_decoder(16#9e#)) OR
 					(reg_q604 AND symb_decoder(16#24#)) OR
 					(reg_q604 AND symb_decoder(16#97#)) OR
 					(reg_q604 AND symb_decoder(16#35#)) OR
 					(reg_q604 AND symb_decoder(16#51#)) OR
 					(reg_q604 AND symb_decoder(16#d0#)) OR
 					(reg_q604 AND symb_decoder(16#2e#)) OR
 					(reg_q604 AND symb_decoder(16#7c#)) OR
 					(reg_q604 AND symb_decoder(16#2f#)) OR
 					(reg_q604 AND symb_decoder(16#12#)) OR
 					(reg_q604 AND symb_decoder(16#ea#)) OR
 					(reg_q604 AND symb_decoder(16#75#)) OR
 					(reg_q604 AND symb_decoder(16#76#)) OR
 					(reg_q604 AND symb_decoder(16#83#)) OR
 					(reg_q604 AND symb_decoder(16#cc#)) OR
 					(reg_q604 AND symb_decoder(16#02#)) OR
 					(reg_q604 AND symb_decoder(16#a3#)) OR
 					(reg_q604 AND symb_decoder(16#59#)) OR
 					(reg_q604 AND symb_decoder(16#cd#)) OR
 					(reg_q604 AND symb_decoder(16#a8#)) OR
 					(reg_q604 AND symb_decoder(16#30#)) OR
 					(reg_q604 AND symb_decoder(16#e2#)) OR
 					(reg_q604 AND symb_decoder(16#38#)) OR
 					(reg_q604 AND symb_decoder(16#47#)) OR
 					(reg_q604 AND symb_decoder(16#52#)) OR
 					(reg_q604 AND symb_decoder(16#f8#)) OR
 					(reg_q604 AND symb_decoder(16#48#)) OR
 					(reg_q604 AND symb_decoder(16#49#)) OR
 					(reg_q604 AND symb_decoder(16#63#)) OR
 					(reg_q604 AND symb_decoder(16#b8#)) OR
 					(reg_q604 AND symb_decoder(16#2a#)) OR
 					(reg_q604 AND symb_decoder(16#10#)) OR
 					(reg_q604 AND symb_decoder(16#ae#)) OR
 					(reg_q604 AND symb_decoder(16#79#)) OR
 					(reg_q604 AND symb_decoder(16#41#)) OR
 					(reg_q604 AND symb_decoder(16#fb#)) OR
 					(reg_q604 AND symb_decoder(16#0d#)) OR
 					(reg_q604 AND symb_decoder(16#c0#)) OR
 					(reg_q604 AND symb_decoder(16#36#)) OR
 					(reg_q604 AND symb_decoder(16#ca#)) OR
 					(reg_q604 AND symb_decoder(16#5f#)) OR
 					(reg_q604 AND symb_decoder(16#f5#)) OR
 					(reg_q604 AND symb_decoder(16#f1#)) OR
 					(reg_q604 AND symb_decoder(16#b0#)) OR
 					(reg_q604 AND symb_decoder(16#45#)) OR
 					(reg_q604 AND symb_decoder(16#ce#)) OR
 					(reg_q604 AND symb_decoder(16#5c#)) OR
 					(reg_q604 AND symb_decoder(16#c1#)) OR
 					(reg_q604 AND symb_decoder(16#dc#)) OR
 					(reg_q604 AND symb_decoder(16#8e#)) OR
 					(reg_q604 AND symb_decoder(16#18#)) OR
 					(reg_q604 AND symb_decoder(16#bb#)) OR
 					(reg_q604 AND symb_decoder(16#86#)) OR
 					(reg_q604 AND symb_decoder(16#ad#)) OR
 					(reg_q604 AND symb_decoder(16#c4#)) OR
 					(reg_q604 AND symb_decoder(16#1e#)) OR
 					(reg_q604 AND symb_decoder(16#fc#)) OR
 					(reg_q604 AND symb_decoder(16#61#)) OR
 					(reg_q604 AND symb_decoder(16#4d#)) OR
 					(reg_q604 AND symb_decoder(16#92#)) OR
 					(reg_q604 AND symb_decoder(16#c3#)) OR
 					(reg_q604 AND symb_decoder(16#55#)) OR
 					(reg_q604 AND symb_decoder(16#43#)) OR
 					(reg_q604 AND symb_decoder(16#08#)) OR
 					(reg_q604 AND symb_decoder(16#8b#)) OR
 					(reg_q604 AND symb_decoder(16#ab#)) OR
 					(reg_q604 AND symb_decoder(16#3a#)) OR
 					(reg_q604 AND symb_decoder(16#e0#)) OR
 					(reg_q604 AND symb_decoder(16#94#)) OR
 					(reg_q604 AND symb_decoder(16#c5#)) OR
 					(reg_q604 AND symb_decoder(16#54#)) OR
 					(reg_q604 AND symb_decoder(16#fd#)) OR
 					(reg_q604 AND symb_decoder(16#60#)) OR
 					(reg_q604 AND symb_decoder(16#9a#)) OR
 					(reg_q604 AND symb_decoder(16#32#)) OR
 					(reg_q604 AND symb_decoder(16#64#)) OR
 					(reg_q604 AND symb_decoder(16#6d#)) OR
 					(reg_q604 AND symb_decoder(16#9d#)) OR
 					(reg_q604 AND symb_decoder(16#b2#)) OR
 					(reg_q604 AND symb_decoder(16#72#)) OR
 					(reg_q604 AND symb_decoder(16#16#)) OR
 					(reg_q604 AND symb_decoder(16#70#)) OR
 					(reg_q604 AND symb_decoder(16#4a#)) OR
 					(reg_q604 AND symb_decoder(16#d8#)) OR
 					(reg_q604 AND symb_decoder(16#01#)) OR
 					(reg_q604 AND symb_decoder(16#5b#)) OR
 					(reg_q604 AND symb_decoder(16#e5#)) OR
 					(reg_q604 AND symb_decoder(16#b5#)) OR
 					(reg_q604 AND symb_decoder(16#af#)) OR
 					(reg_q604 AND symb_decoder(16#f7#)) OR
 					(reg_q604 AND symb_decoder(16#c7#)) OR
 					(reg_q604 AND symb_decoder(16#58#)) OR
 					(reg_q604 AND symb_decoder(16#33#)) OR
 					(reg_q604 AND symb_decoder(16#d2#)) OR
 					(reg_q604 AND symb_decoder(16#d3#)) OR
 					(reg_q604 AND symb_decoder(16#6c#)) OR
 					(reg_q604 AND symb_decoder(16#06#)) OR
 					(reg_q604 AND symb_decoder(16#1d#)) OR
 					(reg_q604 AND symb_decoder(16#66#)) OR
 					(reg_q604 AND symb_decoder(16#c9#)) OR
 					(reg_q604 AND symb_decoder(16#03#)) OR
 					(reg_q604 AND symb_decoder(16#07#)) OR
 					(reg_q604 AND symb_decoder(16#85#)) OR
 					(reg_q604 AND symb_decoder(16#5a#)) OR
 					(reg_q604 AND symb_decoder(16#50#)) OR
 					(reg_q604 AND symb_decoder(16#7d#)) OR
 					(reg_q604 AND symb_decoder(16#57#)) OR
 					(reg_q604 AND symb_decoder(16#99#)) OR
 					(reg_q604 AND symb_decoder(16#80#)) OR
 					(reg_q604 AND symb_decoder(16#cb#)) OR
 					(reg_q604 AND symb_decoder(16#44#)) OR
 					(reg_q604 AND symb_decoder(16#27#)) OR
 					(reg_q604 AND symb_decoder(16#f6#)) OR
 					(reg_q604 AND symb_decoder(16#84#)) OR
 					(reg_q604 AND symb_decoder(16#ee#)) OR
 					(reg_q604 AND symb_decoder(16#9c#)) OR
 					(reg_q604 AND symb_decoder(16#dd#)) OR
 					(reg_q604 AND symb_decoder(16#e7#)) OR
 					(reg_q604 AND symb_decoder(16#81#)) OR
 					(reg_q604 AND symb_decoder(16#b9#)) OR
 					(reg_q604 AND symb_decoder(16#6a#)) OR
 					(reg_q604 AND symb_decoder(16#88#)) OR
 					(reg_q604 AND symb_decoder(16#7f#)) OR
 					(reg_q604 AND symb_decoder(16#1f#)) OR
 					(reg_q604 AND symb_decoder(16#e3#)) OR
 					(reg_q604 AND symb_decoder(16#20#)) OR
 					(reg_q604 AND symb_decoder(16#f2#)) OR
 					(reg_q604 AND symb_decoder(16#5e#)) OR
 					(reg_q604 AND symb_decoder(16#fe#)) OR
 					(reg_q604 AND symb_decoder(16#62#)) OR
 					(reg_q604 AND symb_decoder(16#a7#)) OR
 					(reg_q604 AND symb_decoder(16#68#)) OR
 					(reg_q604 AND symb_decoder(16#89#)) OR
 					(reg_q604 AND symb_decoder(16#8a#)) OR
 					(reg_q604 AND symb_decoder(16#2b#)) OR
 					(reg_q604 AND symb_decoder(16#3c#)) OR
 					(reg_q604 AND symb_decoder(16#95#)) OR
 					(reg_q604 AND symb_decoder(16#0f#)) OR
 					(reg_q604 AND symb_decoder(16#46#)) OR
 					(reg_q604 AND symb_decoder(16#23#)) OR
 					(reg_q604 AND symb_decoder(16#93#)) OR
 					(reg_q604 AND symb_decoder(16#b3#)) OR
 					(reg_q604 AND symb_decoder(16#29#)) OR
 					(reg_q604 AND symb_decoder(16#90#)) OR
 					(reg_q604 AND symb_decoder(16#8f#)) OR
 					(reg_q604 AND symb_decoder(16#3b#)) OR
 					(reg_q604 AND symb_decoder(16#d5#));
reg_q604_init <= '0' ;
	p_reg_q604: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q604 <= reg_q604_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q604 <= reg_q604_init;
        else
          reg_q604 <= reg_q604_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1574_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1574 AND symb_decoder(16#11#)) OR
 					(reg_q1574 AND symb_decoder(16#88#)) OR
 					(reg_q1574 AND symb_decoder(16#f8#)) OR
 					(reg_q1574 AND symb_decoder(16#a2#)) OR
 					(reg_q1574 AND symb_decoder(16#39#)) OR
 					(reg_q1574 AND symb_decoder(16#24#)) OR
 					(reg_q1574 AND symb_decoder(16#1f#)) OR
 					(reg_q1574 AND symb_decoder(16#b7#)) OR
 					(reg_q1574 AND symb_decoder(16#84#)) OR
 					(reg_q1574 AND symb_decoder(16#b8#)) OR
 					(reg_q1574 AND symb_decoder(16#09#)) OR
 					(reg_q1574 AND symb_decoder(16#4d#)) OR
 					(reg_q1574 AND symb_decoder(16#3b#)) OR
 					(reg_q1574 AND symb_decoder(16#0c#)) OR
 					(reg_q1574 AND symb_decoder(16#ed#)) OR
 					(reg_q1574 AND symb_decoder(16#2e#)) OR
 					(reg_q1574 AND symb_decoder(16#19#)) OR
 					(reg_q1574 AND symb_decoder(16#db#)) OR
 					(reg_q1574 AND symb_decoder(16#ea#)) OR
 					(reg_q1574 AND symb_decoder(16#17#)) OR
 					(reg_q1574 AND symb_decoder(16#03#)) OR
 					(reg_q1574 AND symb_decoder(16#bf#)) OR
 					(reg_q1574 AND symb_decoder(16#72#)) OR
 					(reg_q1574 AND symb_decoder(16#32#)) OR
 					(reg_q1574 AND symb_decoder(16#a6#)) OR
 					(reg_q1574 AND symb_decoder(16#e1#)) OR
 					(reg_q1574 AND symb_decoder(16#95#)) OR
 					(reg_q1574 AND symb_decoder(16#dc#)) OR
 					(reg_q1574 AND symb_decoder(16#75#)) OR
 					(reg_q1574 AND symb_decoder(16#7a#)) OR
 					(reg_q1574 AND symb_decoder(16#53#)) OR
 					(reg_q1574 AND symb_decoder(16#b4#)) OR
 					(reg_q1574 AND symb_decoder(16#ce#)) OR
 					(reg_q1574 AND symb_decoder(16#2b#)) OR
 					(reg_q1574 AND symb_decoder(16#68#)) OR
 					(reg_q1574 AND symb_decoder(16#eb#)) OR
 					(reg_q1574 AND symb_decoder(16#6f#)) OR
 					(reg_q1574 AND symb_decoder(16#48#)) OR
 					(reg_q1574 AND symb_decoder(16#42#)) OR
 					(reg_q1574 AND symb_decoder(16#06#)) OR
 					(reg_q1574 AND symb_decoder(16#af#)) OR
 					(reg_q1574 AND symb_decoder(16#ef#)) OR
 					(reg_q1574 AND symb_decoder(16#ba#)) OR
 					(reg_q1574 AND symb_decoder(16#a3#)) OR
 					(reg_q1574 AND symb_decoder(16#8b#)) OR
 					(reg_q1574 AND symb_decoder(16#ca#)) OR
 					(reg_q1574 AND symb_decoder(16#c2#)) OR
 					(reg_q1574 AND symb_decoder(16#29#)) OR
 					(reg_q1574 AND symb_decoder(16#b3#)) OR
 					(reg_q1574 AND symb_decoder(16#d3#)) OR
 					(reg_q1574 AND symb_decoder(16#d6#)) OR
 					(reg_q1574 AND symb_decoder(16#89#)) OR
 					(reg_q1574 AND symb_decoder(16#73#)) OR
 					(reg_q1574 AND symb_decoder(16#fc#)) OR
 					(reg_q1574 AND symb_decoder(16#ee#)) OR
 					(reg_q1574 AND symb_decoder(16#ad#)) OR
 					(reg_q1574 AND symb_decoder(16#8f#)) OR
 					(reg_q1574 AND symb_decoder(16#a5#)) OR
 					(reg_q1574 AND symb_decoder(16#4e#)) OR
 					(reg_q1574 AND symb_decoder(16#85#)) OR
 					(reg_q1574 AND symb_decoder(16#79#)) OR
 					(reg_q1574 AND symb_decoder(16#64#)) OR
 					(reg_q1574 AND symb_decoder(16#fa#)) OR
 					(reg_q1574 AND symb_decoder(16#b5#)) OR
 					(reg_q1574 AND symb_decoder(16#e6#)) OR
 					(reg_q1574 AND symb_decoder(16#69#)) OR
 					(reg_q1574 AND symb_decoder(16#e0#)) OR
 					(reg_q1574 AND symb_decoder(16#be#)) OR
 					(reg_q1574 AND symb_decoder(16#d4#)) OR
 					(reg_q1574 AND symb_decoder(16#33#)) OR
 					(reg_q1574 AND symb_decoder(16#45#)) OR
 					(reg_q1574 AND symb_decoder(16#52#)) OR
 					(reg_q1574 AND symb_decoder(16#a7#)) OR
 					(reg_q1574 AND symb_decoder(16#67#)) OR
 					(reg_q1574 AND symb_decoder(16#f4#)) OR
 					(reg_q1574 AND symb_decoder(16#82#)) OR
 					(reg_q1574 AND symb_decoder(16#f3#)) OR
 					(reg_q1574 AND symb_decoder(16#fe#)) OR
 					(reg_q1574 AND symb_decoder(16#05#)) OR
 					(reg_q1574 AND symb_decoder(16#37#)) OR
 					(reg_q1574 AND symb_decoder(16#aa#)) OR
 					(reg_q1574 AND symb_decoder(16#83#)) OR
 					(reg_q1574 AND symb_decoder(16#10#)) OR
 					(reg_q1574 AND symb_decoder(16#d7#)) OR
 					(reg_q1574 AND symb_decoder(16#01#)) OR
 					(reg_q1574 AND symb_decoder(16#43#)) OR
 					(reg_q1574 AND symb_decoder(16#04#)) OR
 					(reg_q1574 AND symb_decoder(16#78#)) OR
 					(reg_q1574 AND symb_decoder(16#f7#)) OR
 					(reg_q1574 AND symb_decoder(16#b0#)) OR
 					(reg_q1574 AND symb_decoder(16#54#)) OR
 					(reg_q1574 AND symb_decoder(16#d5#)) OR
 					(reg_q1574 AND symb_decoder(16#3a#)) OR
 					(reg_q1574 AND symb_decoder(16#55#)) OR
 					(reg_q1574 AND symb_decoder(16#31#)) OR
 					(reg_q1574 AND symb_decoder(16#b1#)) OR
 					(reg_q1574 AND symb_decoder(16#49#)) OR
 					(reg_q1574 AND symb_decoder(16#30#)) OR
 					(reg_q1574 AND symb_decoder(16#fd#)) OR
 					(reg_q1574 AND symb_decoder(16#57#)) OR
 					(reg_q1574 AND symb_decoder(16#22#)) OR
 					(reg_q1574 AND symb_decoder(16#87#)) OR
 					(reg_q1574 AND symb_decoder(16#94#)) OR
 					(reg_q1574 AND symb_decoder(16#de#)) OR
 					(reg_q1574 AND symb_decoder(16#a4#)) OR
 					(reg_q1574 AND symb_decoder(16#c4#)) OR
 					(reg_q1574 AND symb_decoder(16#f1#)) OR
 					(reg_q1574 AND symb_decoder(16#9d#)) OR
 					(reg_q1574 AND symb_decoder(16#93#)) OR
 					(reg_q1574 AND symb_decoder(16#6a#)) OR
 					(reg_q1574 AND symb_decoder(16#1d#)) OR
 					(reg_q1574 AND symb_decoder(16#d9#)) OR
 					(reg_q1574 AND symb_decoder(16#02#)) OR
 					(reg_q1574 AND symb_decoder(16#9b#)) OR
 					(reg_q1574 AND symb_decoder(16#4b#)) OR
 					(reg_q1574 AND symb_decoder(16#26#)) OR
 					(reg_q1574 AND symb_decoder(16#00#)) OR
 					(reg_q1574 AND symb_decoder(16#9a#)) OR
 					(reg_q1574 AND symb_decoder(16#21#)) OR
 					(reg_q1574 AND symb_decoder(16#70#)) OR
 					(reg_q1574 AND symb_decoder(16#0d#)) OR
 					(reg_q1574 AND symb_decoder(16#15#)) OR
 					(reg_q1574 AND symb_decoder(16#9c#)) OR
 					(reg_q1574 AND symb_decoder(16#cf#)) OR
 					(reg_q1574 AND symb_decoder(16#da#)) OR
 					(reg_q1574 AND symb_decoder(16#4a#)) OR
 					(reg_q1574 AND symb_decoder(16#38#)) OR
 					(reg_q1574 AND symb_decoder(16#96#)) OR
 					(reg_q1574 AND symb_decoder(16#ec#)) OR
 					(reg_q1574 AND symb_decoder(16#81#)) OR
 					(reg_q1574 AND symb_decoder(16#cc#)) OR
 					(reg_q1574 AND symb_decoder(16#e3#)) OR
 					(reg_q1574 AND symb_decoder(16#20#)) OR
 					(reg_q1574 AND symb_decoder(16#d2#)) OR
 					(reg_q1574 AND symb_decoder(16#63#)) OR
 					(reg_q1574 AND symb_decoder(16#62#)) OR
 					(reg_q1574 AND symb_decoder(16#86#)) OR
 					(reg_q1574 AND symb_decoder(16#13#)) OR
 					(reg_q1574 AND symb_decoder(16#bd#)) OR
 					(reg_q1574 AND symb_decoder(16#f6#)) OR
 					(reg_q1574 AND symb_decoder(16#61#)) OR
 					(reg_q1574 AND symb_decoder(16#6c#)) OR
 					(reg_q1574 AND symb_decoder(16#2c#)) OR
 					(reg_q1574 AND symb_decoder(16#ac#)) OR
 					(reg_q1574 AND symb_decoder(16#91#)) OR
 					(reg_q1574 AND symb_decoder(16#9e#)) OR
 					(reg_q1574 AND symb_decoder(16#50#)) OR
 					(reg_q1574 AND symb_decoder(16#12#)) OR
 					(reg_q1574 AND symb_decoder(16#cb#)) OR
 					(reg_q1574 AND symb_decoder(16#07#)) OR
 					(reg_q1574 AND symb_decoder(16#6d#)) OR
 					(reg_q1574 AND symb_decoder(16#e2#)) OR
 					(reg_q1574 AND symb_decoder(16#a8#)) OR
 					(reg_q1574 AND symb_decoder(16#7c#)) OR
 					(reg_q1574 AND symb_decoder(16#ab#)) OR
 					(reg_q1574 AND symb_decoder(16#c9#)) OR
 					(reg_q1574 AND symb_decoder(16#8a#)) OR
 					(reg_q1574 AND symb_decoder(16#ae#)) OR
 					(reg_q1574 AND symb_decoder(16#76#)) OR
 					(reg_q1574 AND symb_decoder(16#3f#)) OR
 					(reg_q1574 AND symb_decoder(16#7f#)) OR
 					(reg_q1574 AND symb_decoder(16#77#)) OR
 					(reg_q1574 AND symb_decoder(16#2f#)) OR
 					(reg_q1574 AND symb_decoder(16#60#)) OR
 					(reg_q1574 AND symb_decoder(16#e7#)) OR
 					(reg_q1574 AND symb_decoder(16#b9#)) OR
 					(reg_q1574 AND symb_decoder(16#80#)) OR
 					(reg_q1574 AND symb_decoder(16#8e#)) OR
 					(reg_q1574 AND symb_decoder(16#5e#)) OR
 					(reg_q1574 AND symb_decoder(16#b2#)) OR
 					(reg_q1574 AND symb_decoder(16#a1#)) OR
 					(reg_q1574 AND symb_decoder(16#f5#)) OR
 					(reg_q1574 AND symb_decoder(16#16#)) OR
 					(reg_q1574 AND symb_decoder(16#71#)) OR
 					(reg_q1574 AND symb_decoder(16#0b#)) OR
 					(reg_q1574 AND symb_decoder(16#3d#)) OR
 					(reg_q1574 AND symb_decoder(16#e4#)) OR
 					(reg_q1574 AND symb_decoder(16#18#)) OR
 					(reg_q1574 AND symb_decoder(16#56#)) OR
 					(reg_q1574 AND symb_decoder(16#5a#)) OR
 					(reg_q1574 AND symb_decoder(16#9f#)) OR
 					(reg_q1574 AND symb_decoder(16#4c#)) OR
 					(reg_q1574 AND symb_decoder(16#c3#)) OR
 					(reg_q1574 AND symb_decoder(16#0a#)) OR
 					(reg_q1574 AND symb_decoder(16#35#)) OR
 					(reg_q1574 AND symb_decoder(16#90#)) OR
 					(reg_q1574 AND symb_decoder(16#8c#)) OR
 					(reg_q1574 AND symb_decoder(16#66#)) OR
 					(reg_q1574 AND symb_decoder(16#6b#)) OR
 					(reg_q1574 AND symb_decoder(16#0f#)) OR
 					(reg_q1574 AND symb_decoder(16#2a#)) OR
 					(reg_q1574 AND symb_decoder(16#74#)) OR
 					(reg_q1574 AND symb_decoder(16#36#)) OR
 					(reg_q1574 AND symb_decoder(16#7e#)) OR
 					(reg_q1574 AND symb_decoder(16#df#)) OR
 					(reg_q1574 AND symb_decoder(16#5b#)) OR
 					(reg_q1574 AND symb_decoder(16#2d#)) OR
 					(reg_q1574 AND symb_decoder(16#1e#)) OR
 					(reg_q1574 AND symb_decoder(16#7d#)) OR
 					(reg_q1574 AND symb_decoder(16#e5#)) OR
 					(reg_q1574 AND symb_decoder(16#d0#)) OR
 					(reg_q1574 AND symb_decoder(16#4f#)) OR
 					(reg_q1574 AND symb_decoder(16#1b#)) OR
 					(reg_q1574 AND symb_decoder(16#14#)) OR
 					(reg_q1574 AND symb_decoder(16#40#)) OR
 					(reg_q1574 AND symb_decoder(16#92#)) OR
 					(reg_q1574 AND symb_decoder(16#97#)) OR
 					(reg_q1574 AND symb_decoder(16#58#)) OR
 					(reg_q1574 AND symb_decoder(16#99#)) OR
 					(reg_q1574 AND symb_decoder(16#28#)) OR
 					(reg_q1574 AND symb_decoder(16#c1#)) OR
 					(reg_q1574 AND symb_decoder(16#8d#)) OR
 					(reg_q1574 AND symb_decoder(16#e9#)) OR
 					(reg_q1574 AND symb_decoder(16#b6#)) OR
 					(reg_q1574 AND symb_decoder(16#c5#)) OR
 					(reg_q1574 AND symb_decoder(16#0e#)) OR
 					(reg_q1574 AND symb_decoder(16#a9#)) OR
 					(reg_q1574 AND symb_decoder(16#fb#)) OR
 					(reg_q1574 AND symb_decoder(16#d8#)) OR
 					(reg_q1574 AND symb_decoder(16#ff#)) OR
 					(reg_q1574 AND symb_decoder(16#1a#)) OR
 					(reg_q1574 AND symb_decoder(16#27#)) OR
 					(reg_q1574 AND symb_decoder(16#6e#)) OR
 					(reg_q1574 AND symb_decoder(16#a0#)) OR
 					(reg_q1574 AND symb_decoder(16#3c#)) OR
 					(reg_q1574 AND symb_decoder(16#41#)) OR
 					(reg_q1574 AND symb_decoder(16#c0#)) OR
 					(reg_q1574 AND symb_decoder(16#23#)) OR
 					(reg_q1574 AND symb_decoder(16#f2#)) OR
 					(reg_q1574 AND symb_decoder(16#51#)) OR
 					(reg_q1574 AND symb_decoder(16#25#)) OR
 					(reg_q1574 AND symb_decoder(16#34#)) OR
 					(reg_q1574 AND symb_decoder(16#f9#)) OR
 					(reg_q1574 AND symb_decoder(16#98#)) OR
 					(reg_q1574 AND symb_decoder(16#bb#)) OR
 					(reg_q1574 AND symb_decoder(16#5f#)) OR
 					(reg_q1574 AND symb_decoder(16#e8#)) OR
 					(reg_q1574 AND symb_decoder(16#7b#)) OR
 					(reg_q1574 AND symb_decoder(16#c8#)) OR
 					(reg_q1574 AND symb_decoder(16#5d#)) OR
 					(reg_q1574 AND symb_decoder(16#47#)) OR
 					(reg_q1574 AND symb_decoder(16#c6#)) OR
 					(reg_q1574 AND symb_decoder(16#1c#)) OR
 					(reg_q1574 AND symb_decoder(16#59#)) OR
 					(reg_q1574 AND symb_decoder(16#c7#)) OR
 					(reg_q1574 AND symb_decoder(16#3e#)) OR
 					(reg_q1574 AND symb_decoder(16#bc#)) OR
 					(reg_q1574 AND symb_decoder(16#46#)) OR
 					(reg_q1574 AND symb_decoder(16#5c#)) OR
 					(reg_q1574 AND symb_decoder(16#08#)) OR
 					(reg_q1574 AND symb_decoder(16#f0#)) OR
 					(reg_q1574 AND symb_decoder(16#44#)) OR
 					(reg_q1574 AND symb_decoder(16#d1#)) OR
 					(reg_q1574 AND symb_decoder(16#65#)) OR
 					(reg_q1574 AND symb_decoder(16#dd#)) OR
 					(reg_q1574 AND symb_decoder(16#cd#));
reg_q1574_init <= '0' ;
	p_reg_q1574: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1574 <= reg_q1574_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1574 <= reg_q1574_init;
        else
          reg_q1574 <= reg_q1574_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph62

reg_q113_in <= (reg_q107 AND symb_decoder(16#03#)) OR
 					(reg_q107 AND symb_decoder(16#29#)) OR
 					(reg_q107 AND symb_decoder(16#f8#)) OR
 					(reg_q107 AND symb_decoder(16#72#)) OR
 					(reg_q107 AND symb_decoder(16#49#)) OR
 					(reg_q107 AND symb_decoder(16#3e#)) OR
 					(reg_q107 AND symb_decoder(16#e7#)) OR
 					(reg_q107 AND symb_decoder(16#f6#)) OR
 					(reg_q107 AND symb_decoder(16#22#)) OR
 					(reg_q107 AND symb_decoder(16#48#)) OR
 					(reg_q107 AND symb_decoder(16#23#)) OR
 					(reg_q107 AND symb_decoder(16#69#)) OR
 					(reg_q107 AND symb_decoder(16#13#)) OR
 					(reg_q107 AND symb_decoder(16#b2#)) OR
 					(reg_q107 AND symb_decoder(16#94#)) OR
 					(reg_q107 AND symb_decoder(16#4b#)) OR
 					(reg_q107 AND symb_decoder(16#a4#)) OR
 					(reg_q107 AND symb_decoder(16#32#)) OR
 					(reg_q107 AND symb_decoder(16#ee#)) OR
 					(reg_q107 AND symb_decoder(16#93#)) OR
 					(reg_q107 AND symb_decoder(16#26#)) OR
 					(reg_q107 AND symb_decoder(16#b0#)) OR
 					(reg_q107 AND symb_decoder(16#52#)) OR
 					(reg_q107 AND symb_decoder(16#80#)) OR
 					(reg_q107 AND symb_decoder(16#27#)) OR
 					(reg_q107 AND symb_decoder(16#b8#)) OR
 					(reg_q107 AND symb_decoder(16#7a#)) OR
 					(reg_q107 AND symb_decoder(16#39#)) OR
 					(reg_q107 AND symb_decoder(16#01#)) OR
 					(reg_q107 AND symb_decoder(16#96#)) OR
 					(reg_q107 AND symb_decoder(16#e9#)) OR
 					(reg_q107 AND symb_decoder(16#59#)) OR
 					(reg_q107 AND symb_decoder(16#71#)) OR
 					(reg_q107 AND symb_decoder(16#74#)) OR
 					(reg_q107 AND symb_decoder(16#3c#)) OR
 					(reg_q107 AND symb_decoder(16#99#)) OR
 					(reg_q107 AND symb_decoder(16#8d#)) OR
 					(reg_q107 AND symb_decoder(16#f7#)) OR
 					(reg_q107 AND symb_decoder(16#e1#)) OR
 					(reg_q107 AND symb_decoder(16#cb#)) OR
 					(reg_q107 AND symb_decoder(16#6a#)) OR
 					(reg_q107 AND symb_decoder(16#c9#)) OR
 					(reg_q107 AND symb_decoder(16#fa#)) OR
 					(reg_q107 AND symb_decoder(16#46#)) OR
 					(reg_q107 AND symb_decoder(16#07#)) OR
 					(reg_q107 AND symb_decoder(16#31#)) OR
 					(reg_q107 AND symb_decoder(16#2d#)) OR
 					(reg_q107 AND symb_decoder(16#65#)) OR
 					(reg_q107 AND symb_decoder(16#f1#)) OR
 					(reg_q107 AND symb_decoder(16#12#)) OR
 					(reg_q107 AND symb_decoder(16#c3#)) OR
 					(reg_q107 AND symb_decoder(16#5d#)) OR
 					(reg_q107 AND symb_decoder(16#90#)) OR
 					(reg_q107 AND symb_decoder(16#98#)) OR
 					(reg_q107 AND symb_decoder(16#c1#)) OR
 					(reg_q107 AND symb_decoder(16#02#)) OR
 					(reg_q107 AND symb_decoder(16#54#)) OR
 					(reg_q107 AND symb_decoder(16#3f#)) OR
 					(reg_q107 AND symb_decoder(16#d7#)) OR
 					(reg_q107 AND symb_decoder(16#aa#)) OR
 					(reg_q107 AND symb_decoder(16#db#)) OR
 					(reg_q107 AND symb_decoder(16#6d#)) OR
 					(reg_q107 AND symb_decoder(16#8c#)) OR
 					(reg_q107 AND symb_decoder(16#1b#)) OR
 					(reg_q107 AND symb_decoder(16#21#)) OR
 					(reg_q107 AND symb_decoder(16#61#)) OR
 					(reg_q107 AND symb_decoder(16#a5#)) OR
 					(reg_q107 AND symb_decoder(16#cc#)) OR
 					(reg_q107 AND symb_decoder(16#0c#)) OR
 					(reg_q107 AND symb_decoder(16#5a#)) OR
 					(reg_q107 AND symb_decoder(16#17#)) OR
 					(reg_q107 AND symb_decoder(16#6f#)) OR
 					(reg_q107 AND symb_decoder(16#36#)) OR
 					(reg_q107 AND symb_decoder(16#55#)) OR
 					(reg_q107 AND symb_decoder(16#b5#)) OR
 					(reg_q107 AND symb_decoder(16#24#)) OR
 					(reg_q107 AND symb_decoder(16#40#)) OR
 					(reg_q107 AND symb_decoder(16#97#)) OR
 					(reg_q107 AND symb_decoder(16#7b#)) OR
 					(reg_q107 AND symb_decoder(16#37#)) OR
 					(reg_q107 AND symb_decoder(16#cd#)) OR
 					(reg_q107 AND symb_decoder(16#53#)) OR
 					(reg_q107 AND symb_decoder(16#ea#)) OR
 					(reg_q107 AND symb_decoder(16#9f#)) OR
 					(reg_q107 AND symb_decoder(16#87#)) OR
 					(reg_q107 AND symb_decoder(16#11#)) OR
 					(reg_q107 AND symb_decoder(16#4f#)) OR
 					(reg_q107 AND symb_decoder(16#d2#)) OR
 					(reg_q107 AND symb_decoder(16#c4#)) OR
 					(reg_q107 AND symb_decoder(16#df#)) OR
 					(reg_q107 AND symb_decoder(16#7c#)) OR
 					(reg_q107 AND symb_decoder(16#83#)) OR
 					(reg_q107 AND symb_decoder(16#1c#)) OR
 					(reg_q107 AND symb_decoder(16#08#)) OR
 					(reg_q107 AND symb_decoder(16#4e#)) OR
 					(reg_q107 AND symb_decoder(16#66#)) OR
 					(reg_q107 AND symb_decoder(16#81#)) OR
 					(reg_q107 AND symb_decoder(16#77#)) OR
 					(reg_q107 AND symb_decoder(16#34#)) OR
 					(reg_q107 AND symb_decoder(16#9b#)) OR
 					(reg_q107 AND symb_decoder(16#c6#)) OR
 					(reg_q107 AND symb_decoder(16#fc#)) OR
 					(reg_q107 AND symb_decoder(16#1f#)) OR
 					(reg_q107 AND symb_decoder(16#d1#)) OR
 					(reg_q107 AND symb_decoder(16#a8#)) OR
 					(reg_q107 AND symb_decoder(16#2b#)) OR
 					(reg_q107 AND symb_decoder(16#43#)) OR
 					(reg_q107 AND symb_decoder(16#8e#)) OR
 					(reg_q107 AND symb_decoder(16#d8#)) OR
 					(reg_q107 AND symb_decoder(16#05#)) OR
 					(reg_q107 AND symb_decoder(16#c7#)) OR
 					(reg_q107 AND symb_decoder(16#d6#)) OR
 					(reg_q107 AND symb_decoder(16#47#)) OR
 					(reg_q107 AND symb_decoder(16#2e#)) OR
 					(reg_q107 AND symb_decoder(16#dd#)) OR
 					(reg_q107 AND symb_decoder(16#20#)) OR
 					(reg_q107 AND symb_decoder(16#63#)) OR
 					(reg_q107 AND symb_decoder(16#14#)) OR
 					(reg_q107 AND symb_decoder(16#19#)) OR
 					(reg_q107 AND symb_decoder(16#e4#)) OR
 					(reg_q107 AND symb_decoder(16#35#)) OR
 					(reg_q107 AND symb_decoder(16#f2#)) OR
 					(reg_q107 AND symb_decoder(16#09#)) OR
 					(reg_q107 AND symb_decoder(16#c8#)) OR
 					(reg_q107 AND symb_decoder(16#c5#)) OR
 					(reg_q107 AND symb_decoder(16#c0#)) OR
 					(reg_q107 AND symb_decoder(16#89#)) OR
 					(reg_q107 AND symb_decoder(16#4d#)) OR
 					(reg_q107 AND symb_decoder(16#85#)) OR
 					(reg_q107 AND symb_decoder(16#6e#)) OR
 					(reg_q107 AND symb_decoder(16#73#)) OR
 					(reg_q107 AND symb_decoder(16#ef#)) OR
 					(reg_q107 AND symb_decoder(16#eb#)) OR
 					(reg_q107 AND symb_decoder(16#04#)) OR
 					(reg_q107 AND symb_decoder(16#bc#)) OR
 					(reg_q107 AND symb_decoder(16#3a#)) OR
 					(reg_q107 AND symb_decoder(16#5f#)) OR
 					(reg_q107 AND symb_decoder(16#33#)) OR
 					(reg_q107 AND symb_decoder(16#ce#)) OR
 					(reg_q107 AND symb_decoder(16#ac#)) OR
 					(reg_q107 AND symb_decoder(16#56#)) OR
 					(reg_q107 AND symb_decoder(16#ec#)) OR
 					(reg_q107 AND symb_decoder(16#f3#)) OR
 					(reg_q107 AND symb_decoder(16#b6#)) OR
 					(reg_q107 AND symb_decoder(16#75#)) OR
 					(reg_q107 AND symb_decoder(16#3b#)) OR
 					(reg_q107 AND symb_decoder(16#25#)) OR
 					(reg_q107 AND symb_decoder(16#2c#)) OR
 					(reg_q107 AND symb_decoder(16#7d#)) OR
 					(reg_q107 AND symb_decoder(16#1e#)) OR
 					(reg_q107 AND symb_decoder(16#78#)) OR
 					(reg_q107 AND symb_decoder(16#0b#)) OR
 					(reg_q107 AND symb_decoder(16#60#)) OR
 					(reg_q107 AND symb_decoder(16#1d#)) OR
 					(reg_q107 AND symb_decoder(16#e6#)) OR
 					(reg_q107 AND symb_decoder(16#fb#)) OR
 					(reg_q107 AND symb_decoder(16#1a#)) OR
 					(reg_q107 AND symb_decoder(16#ed#)) OR
 					(reg_q107 AND symb_decoder(16#d3#)) OR
 					(reg_q107 AND symb_decoder(16#3d#)) OR
 					(reg_q107 AND symb_decoder(16#8b#)) OR
 					(reg_q107 AND symb_decoder(16#ad#)) OR
 					(reg_q107 AND symb_decoder(16#76#)) OR
 					(reg_q107 AND symb_decoder(16#41#)) OR
 					(reg_q107 AND symb_decoder(16#18#)) OR
 					(reg_q107 AND symb_decoder(16#b1#)) OR
 					(reg_q107 AND symb_decoder(16#ab#)) OR
 					(reg_q107 AND symb_decoder(16#2f#)) OR
 					(reg_q107 AND symb_decoder(16#30#)) OR
 					(reg_q107 AND symb_decoder(16#06#)) OR
 					(reg_q107 AND symb_decoder(16#10#)) OR
 					(reg_q107 AND symb_decoder(16#82#)) OR
 					(reg_q107 AND symb_decoder(16#f0#)) OR
 					(reg_q107 AND symb_decoder(16#b3#)) OR
 					(reg_q107 AND symb_decoder(16#ba#)) OR
 					(reg_q107 AND symb_decoder(16#af#)) OR
 					(reg_q107 AND symb_decoder(16#15#)) OR
 					(reg_q107 AND symb_decoder(16#7f#)) OR
 					(reg_q107 AND symb_decoder(16#79#)) OR
 					(reg_q107 AND symb_decoder(16#5e#)) OR
 					(reg_q107 AND symb_decoder(16#67#)) OR
 					(reg_q107 AND symb_decoder(16#5b#)) OR
 					(reg_q107 AND symb_decoder(16#e0#)) OR
 					(reg_q107 AND symb_decoder(16#9e#)) OR
 					(reg_q107 AND symb_decoder(16#16#)) OR
 					(reg_q107 AND symb_decoder(16#ca#)) OR
 					(reg_q107 AND symb_decoder(16#dc#)) OR
 					(reg_q107 AND symb_decoder(16#00#)) OR
 					(reg_q107 AND symb_decoder(16#68#)) OR
 					(reg_q107 AND symb_decoder(16#ff#)) OR
 					(reg_q107 AND symb_decoder(16#86#)) OR
 					(reg_q107 AND symb_decoder(16#91#)) OR
 					(reg_q107 AND symb_decoder(16#c2#)) OR
 					(reg_q107 AND symb_decoder(16#9a#)) OR
 					(reg_q107 AND symb_decoder(16#45#)) OR
 					(reg_q107 AND symb_decoder(16#50#)) OR
 					(reg_q107 AND symb_decoder(16#e2#)) OR
 					(reg_q107 AND symb_decoder(16#ae#)) OR
 					(reg_q107 AND symb_decoder(16#6c#)) OR
 					(reg_q107 AND symb_decoder(16#f4#)) OR
 					(reg_q107 AND symb_decoder(16#9d#)) OR
 					(reg_q107 AND symb_decoder(16#0f#)) OR
 					(reg_q107 AND symb_decoder(16#e8#)) OR
 					(reg_q107 AND symb_decoder(16#d0#)) OR
 					(reg_q107 AND symb_decoder(16#8a#)) OR
 					(reg_q107 AND symb_decoder(16#28#)) OR
 					(reg_q107 AND symb_decoder(16#be#)) OR
 					(reg_q107 AND symb_decoder(16#a7#)) OR
 					(reg_q107 AND symb_decoder(16#bf#)) OR
 					(reg_q107 AND symb_decoder(16#b7#)) OR
 					(reg_q107 AND symb_decoder(16#92#)) OR
 					(reg_q107 AND symb_decoder(16#4c#)) OR
 					(reg_q107 AND symb_decoder(16#a9#)) OR
 					(reg_q107 AND symb_decoder(16#fd#)) OR
 					(reg_q107 AND symb_decoder(16#0e#)) OR
 					(reg_q107 AND symb_decoder(16#7e#)) OR
 					(reg_q107 AND symb_decoder(16#38#)) OR
 					(reg_q107 AND symb_decoder(16#64#)) OR
 					(reg_q107 AND symb_decoder(16#a0#)) OR
 					(reg_q107 AND symb_decoder(16#62#)) OR
 					(reg_q107 AND symb_decoder(16#a6#)) OR
 					(reg_q107 AND symb_decoder(16#88#)) OR
 					(reg_q107 AND symb_decoder(16#57#)) OR
 					(reg_q107 AND symb_decoder(16#4a#)) OR
 					(reg_q107 AND symb_decoder(16#d9#)) OR
 					(reg_q107 AND symb_decoder(16#42#)) OR
 					(reg_q107 AND symb_decoder(16#8f#)) OR
 					(reg_q107 AND symb_decoder(16#44#)) OR
 					(reg_q107 AND symb_decoder(16#84#)) OR
 					(reg_q107 AND symb_decoder(16#5c#)) OR
 					(reg_q107 AND symb_decoder(16#fe#)) OR
 					(reg_q107 AND symb_decoder(16#a1#)) OR
 					(reg_q107 AND symb_decoder(16#de#)) OR
 					(reg_q107 AND symb_decoder(16#95#)) OR
 					(reg_q107 AND symb_decoder(16#a2#)) OR
 					(reg_q107 AND symb_decoder(16#e5#)) OR
 					(reg_q107 AND symb_decoder(16#58#)) OR
 					(reg_q107 AND symb_decoder(16#6b#)) OR
 					(reg_q107 AND symb_decoder(16#51#)) OR
 					(reg_q107 AND symb_decoder(16#d5#)) OR
 					(reg_q107 AND symb_decoder(16#b4#)) OR
 					(reg_q107 AND symb_decoder(16#e3#)) OR
 					(reg_q107 AND symb_decoder(16#f5#)) OR
 					(reg_q107 AND symb_decoder(16#b9#)) OR
 					(reg_q107 AND symb_decoder(16#cf#)) OR
 					(reg_q107 AND symb_decoder(16#9c#)) OR
 					(reg_q107 AND symb_decoder(16#70#)) OR
 					(reg_q107 AND symb_decoder(16#bb#)) OR
 					(reg_q107 AND symb_decoder(16#da#)) OR
 					(reg_q107 AND symb_decoder(16#bd#)) OR
 					(reg_q107 AND symb_decoder(16#d4#)) OR
 					(reg_q107 AND symb_decoder(16#f9#)) OR
 					(reg_q107 AND symb_decoder(16#a3#)) OR
 					(reg_q107 AND symb_decoder(16#2a#)) OR
 					(reg_q113 AND symb_decoder(16#69#)) OR
 					(reg_q113 AND symb_decoder(16#00#)) OR
 					(reg_q113 AND symb_decoder(16#da#)) OR
 					(reg_q113 AND symb_decoder(16#27#)) OR
 					(reg_q113 AND symb_decoder(16#5d#)) OR
 					(reg_q113 AND symb_decoder(16#33#)) OR
 					(reg_q113 AND symb_decoder(16#ed#)) OR
 					(reg_q113 AND symb_decoder(16#c2#)) OR
 					(reg_q113 AND symb_decoder(16#e5#)) OR
 					(reg_q113 AND symb_decoder(16#d2#)) OR
 					(reg_q113 AND symb_decoder(16#79#)) OR
 					(reg_q113 AND symb_decoder(16#18#)) OR
 					(reg_q113 AND symb_decoder(16#66#)) OR
 					(reg_q113 AND symb_decoder(16#15#)) OR
 					(reg_q113 AND symb_decoder(16#8f#)) OR
 					(reg_q113 AND symb_decoder(16#a5#)) OR
 					(reg_q113 AND symb_decoder(16#a7#)) OR
 					(reg_q113 AND symb_decoder(16#ea#)) OR
 					(reg_q113 AND symb_decoder(16#7e#)) OR
 					(reg_q113 AND symb_decoder(16#4e#)) OR
 					(reg_q113 AND symb_decoder(16#fc#)) OR
 					(reg_q113 AND symb_decoder(16#0f#)) OR
 					(reg_q113 AND symb_decoder(16#d5#)) OR
 					(reg_q113 AND symb_decoder(16#f5#)) OR
 					(reg_q113 AND symb_decoder(16#82#)) OR
 					(reg_q113 AND symb_decoder(16#d9#)) OR
 					(reg_q113 AND symb_decoder(16#45#)) OR
 					(reg_q113 AND symb_decoder(16#c5#)) OR
 					(reg_q113 AND symb_decoder(16#f6#)) OR
 					(reg_q113 AND symb_decoder(16#d1#)) OR
 					(reg_q113 AND symb_decoder(16#25#)) OR
 					(reg_q113 AND symb_decoder(16#14#)) OR
 					(reg_q113 AND symb_decoder(16#4a#)) OR
 					(reg_q113 AND symb_decoder(16#2d#)) OR
 					(reg_q113 AND symb_decoder(16#ca#)) OR
 					(reg_q113 AND symb_decoder(16#38#)) OR
 					(reg_q113 AND symb_decoder(16#7c#)) OR
 					(reg_q113 AND symb_decoder(16#13#)) OR
 					(reg_q113 AND symb_decoder(16#c3#)) OR
 					(reg_q113 AND symb_decoder(16#e6#)) OR
 					(reg_q113 AND symb_decoder(16#91#)) OR
 					(reg_q113 AND symb_decoder(16#6e#)) OR
 					(reg_q113 AND symb_decoder(16#f3#)) OR
 					(reg_q113 AND symb_decoder(16#d6#)) OR
 					(reg_q113 AND symb_decoder(16#e2#)) OR
 					(reg_q113 AND symb_decoder(16#a2#)) OR
 					(reg_q113 AND symb_decoder(16#aa#)) OR
 					(reg_q113 AND symb_decoder(16#db#)) OR
 					(reg_q113 AND symb_decoder(16#21#)) OR
 					(reg_q113 AND symb_decoder(16#4d#)) OR
 					(reg_q113 AND symb_decoder(16#7d#)) OR
 					(reg_q113 AND symb_decoder(16#b4#)) OR
 					(reg_q113 AND symb_decoder(16#9e#)) OR
 					(reg_q113 AND symb_decoder(16#cf#)) OR
 					(reg_q113 AND symb_decoder(16#eb#)) OR
 					(reg_q113 AND symb_decoder(16#5f#)) OR
 					(reg_q113 AND symb_decoder(16#1f#)) OR
 					(reg_q113 AND symb_decoder(16#9c#)) OR
 					(reg_q113 AND symb_decoder(16#04#)) OR
 					(reg_q113 AND symb_decoder(16#09#)) OR
 					(reg_q113 AND symb_decoder(16#b5#)) OR
 					(reg_q113 AND symb_decoder(16#23#)) OR
 					(reg_q113 AND symb_decoder(16#fd#)) OR
 					(reg_q113 AND symb_decoder(16#81#)) OR
 					(reg_q113 AND symb_decoder(16#b2#)) OR
 					(reg_q113 AND symb_decoder(16#46#)) OR
 					(reg_q113 AND symb_decoder(16#a3#)) OR
 					(reg_q113 AND symb_decoder(16#2f#)) OR
 					(reg_q113 AND symb_decoder(16#c6#)) OR
 					(reg_q113 AND symb_decoder(16#cd#)) OR
 					(reg_q113 AND symb_decoder(16#2c#)) OR
 					(reg_q113 AND symb_decoder(16#dc#)) OR
 					(reg_q113 AND symb_decoder(16#87#)) OR
 					(reg_q113 AND symb_decoder(16#30#)) OR
 					(reg_q113 AND symb_decoder(16#ee#)) OR
 					(reg_q113 AND symb_decoder(16#73#)) OR
 					(reg_q113 AND symb_decoder(16#2e#)) OR
 					(reg_q113 AND symb_decoder(16#a6#)) OR
 					(reg_q113 AND symb_decoder(16#e1#)) OR
 					(reg_q113 AND symb_decoder(16#5b#)) OR
 					(reg_q113 AND symb_decoder(16#39#)) OR
 					(reg_q113 AND symb_decoder(16#75#)) OR
 					(reg_q113 AND symb_decoder(16#44#)) OR
 					(reg_q113 AND symb_decoder(16#6d#)) OR
 					(reg_q113 AND symb_decoder(16#80#)) OR
 					(reg_q113 AND symb_decoder(16#76#)) OR
 					(reg_q113 AND symb_decoder(16#be#)) OR
 					(reg_q113 AND symb_decoder(16#d4#)) OR
 					(reg_q113 AND symb_decoder(16#f8#)) OR
 					(reg_q113 AND symb_decoder(16#b9#)) OR
 					(reg_q113 AND symb_decoder(16#5e#)) OR
 					(reg_q113 AND symb_decoder(16#67#)) OR
 					(reg_q113 AND symb_decoder(16#28#)) OR
 					(reg_q113 AND symb_decoder(16#85#)) OR
 					(reg_q113 AND symb_decoder(16#05#)) OR
 					(reg_q113 AND symb_decoder(16#96#)) OR
 					(reg_q113 AND symb_decoder(16#50#)) OR
 					(reg_q113 AND symb_decoder(16#53#)) OR
 					(reg_q113 AND symb_decoder(16#f9#)) OR
 					(reg_q113 AND symb_decoder(16#40#)) OR
 					(reg_q113 AND symb_decoder(16#78#)) OR
 					(reg_q113 AND symb_decoder(16#70#)) OR
 					(reg_q113 AND symb_decoder(16#f4#)) OR
 					(reg_q113 AND symb_decoder(16#94#)) OR
 					(reg_q113 AND symb_decoder(16#0e#)) OR
 					(reg_q113 AND symb_decoder(16#54#)) OR
 					(reg_q113 AND symb_decoder(16#61#)) OR
 					(reg_q113 AND symb_decoder(16#ba#)) OR
 					(reg_q113 AND symb_decoder(16#5a#)) OR
 					(reg_q113 AND symb_decoder(16#88#)) OR
 					(reg_q113 AND symb_decoder(16#99#)) OR
 					(reg_q113 AND symb_decoder(16#a0#)) OR
 					(reg_q113 AND symb_decoder(16#7a#)) OR
 					(reg_q113 AND symb_decoder(16#ff#)) OR
 					(reg_q113 AND symb_decoder(16#47#)) OR
 					(reg_q113 AND symb_decoder(16#43#)) OR
 					(reg_q113 AND symb_decoder(16#6c#)) OR
 					(reg_q113 AND symb_decoder(16#02#)) OR
 					(reg_q113 AND symb_decoder(16#37#)) OR
 					(reg_q113 AND symb_decoder(16#64#)) OR
 					(reg_q113 AND symb_decoder(16#6b#)) OR
 					(reg_q113 AND symb_decoder(16#32#)) OR
 					(reg_q113 AND symb_decoder(16#9a#)) OR
 					(reg_q113 AND symb_decoder(16#1a#)) OR
 					(reg_q113 AND symb_decoder(16#b0#)) OR
 					(reg_q113 AND symb_decoder(16#e8#)) OR
 					(reg_q113 AND symb_decoder(16#71#)) OR
 					(reg_q113 AND symb_decoder(16#29#)) OR
 					(reg_q113 AND symb_decoder(16#8c#)) OR
 					(reg_q113 AND symb_decoder(16#c1#)) OR
 					(reg_q113 AND symb_decoder(16#49#)) OR
 					(reg_q113 AND symb_decoder(16#60#)) OR
 					(reg_q113 AND symb_decoder(16#16#)) OR
 					(reg_q113 AND symb_decoder(16#84#)) OR
 					(reg_q113 AND symb_decoder(16#98#)) OR
 					(reg_q113 AND symb_decoder(16#26#)) OR
 					(reg_q113 AND symb_decoder(16#52#)) OR
 					(reg_q113 AND symb_decoder(16#93#)) OR
 					(reg_q113 AND symb_decoder(16#bb#)) OR
 					(reg_q113 AND symb_decoder(16#ab#)) OR
 					(reg_q113 AND symb_decoder(16#31#)) OR
 					(reg_q113 AND symb_decoder(16#b3#)) OR
 					(reg_q113 AND symb_decoder(16#77#)) OR
 					(reg_q113 AND symb_decoder(16#8d#)) OR
 					(reg_q113 AND symb_decoder(16#dd#)) OR
 					(reg_q113 AND symb_decoder(16#1d#)) OR
 					(reg_q113 AND symb_decoder(16#a1#)) OR
 					(reg_q113 AND symb_decoder(16#55#)) OR
 					(reg_q113 AND symb_decoder(16#34#)) OR
 					(reg_q113 AND symb_decoder(16#c4#)) OR
 					(reg_q113 AND symb_decoder(16#63#)) OR
 					(reg_q113 AND symb_decoder(16#9b#)) OR
 					(reg_q113 AND symb_decoder(16#6f#)) OR
 					(reg_q113 AND symb_decoder(16#68#)) OR
 					(reg_q113 AND symb_decoder(16#a4#)) OR
 					(reg_q113 AND symb_decoder(16#41#)) OR
 					(reg_q113 AND symb_decoder(16#d7#)) OR
 					(reg_q113 AND symb_decoder(16#f7#)) OR
 					(reg_q113 AND symb_decoder(16#cb#)) OR
 					(reg_q113 AND symb_decoder(16#17#)) OR
 					(reg_q113 AND symb_decoder(16#3e#)) OR
 					(reg_q113 AND symb_decoder(16#ef#)) OR
 					(reg_q113 AND symb_decoder(16#2a#)) OR
 					(reg_q113 AND symb_decoder(16#bf#)) OR
 					(reg_q113 AND symb_decoder(16#95#)) OR
 					(reg_q113 AND symb_decoder(16#0c#)) OR
 					(reg_q113 AND symb_decoder(16#f2#)) OR
 					(reg_q113 AND symb_decoder(16#72#)) OR
 					(reg_q113 AND symb_decoder(16#36#)) OR
 					(reg_q113 AND symb_decoder(16#ac#)) OR
 					(reg_q113 AND symb_decoder(16#92#)) OR
 					(reg_q113 AND symb_decoder(16#1c#)) OR
 					(reg_q113 AND symb_decoder(16#c0#)) OR
 					(reg_q113 AND symb_decoder(16#d8#)) OR
 					(reg_q113 AND symb_decoder(16#3a#)) OR
 					(reg_q113 AND symb_decoder(16#df#)) OR
 					(reg_q113 AND symb_decoder(16#35#)) OR
 					(reg_q113 AND symb_decoder(16#3c#)) OR
 					(reg_q113 AND symb_decoder(16#2b#)) OR
 					(reg_q113 AND symb_decoder(16#01#)) OR
 					(reg_q113 AND symb_decoder(16#bc#)) OR
 					(reg_q113 AND symb_decoder(16#af#)) OR
 					(reg_q113 AND symb_decoder(16#de#)) OR
 					(reg_q113 AND symb_decoder(16#c8#)) OR
 					(reg_q113 AND symb_decoder(16#57#)) OR
 					(reg_q113 AND symb_decoder(16#3f#)) OR
 					(reg_q113 AND symb_decoder(16#59#)) OR
 					(reg_q113 AND symb_decoder(16#b8#)) OR
 					(reg_q113 AND symb_decoder(16#f1#)) OR
 					(reg_q113 AND symb_decoder(16#4b#)) OR
 					(reg_q113 AND symb_decoder(16#03#)) OR
 					(reg_q113 AND symb_decoder(16#bd#)) OR
 					(reg_q113 AND symb_decoder(16#a9#)) OR
 					(reg_q113 AND symb_decoder(16#fe#)) OR
 					(reg_q113 AND symb_decoder(16#3d#)) OR
 					(reg_q113 AND symb_decoder(16#6a#)) OR
 					(reg_q113 AND symb_decoder(16#8e#)) OR
 					(reg_q113 AND symb_decoder(16#19#)) OR
 					(reg_q113 AND symb_decoder(16#20#)) OR
 					(reg_q113 AND symb_decoder(16#74#)) OR
 					(reg_q113 AND symb_decoder(16#c7#)) OR
 					(reg_q113 AND symb_decoder(16#f0#)) OR
 					(reg_q113 AND symb_decoder(16#ae#)) OR
 					(reg_q113 AND symb_decoder(16#58#)) OR
 					(reg_q113 AND symb_decoder(16#51#)) OR
 					(reg_q113 AND symb_decoder(16#e7#)) OR
 					(reg_q113 AND symb_decoder(16#48#)) OR
 					(reg_q113 AND symb_decoder(16#90#)) OR
 					(reg_q113 AND symb_decoder(16#0b#)) OR
 					(reg_q113 AND symb_decoder(16#1e#)) OR
 					(reg_q113 AND symb_decoder(16#06#)) OR
 					(reg_q113 AND symb_decoder(16#fa#)) OR
 					(reg_q113 AND symb_decoder(16#9f#)) OR
 					(reg_q113 AND symb_decoder(16#65#)) OR
 					(reg_q113 AND symb_decoder(16#97#)) OR
 					(reg_q113 AND symb_decoder(16#5c#)) OR
 					(reg_q113 AND symb_decoder(16#7b#)) OR
 					(reg_q113 AND symb_decoder(16#8a#)) OR
 					(reg_q113 AND symb_decoder(16#83#)) OR
 					(reg_q113 AND symb_decoder(16#4c#)) OR
 					(reg_q113 AND symb_decoder(16#8b#)) OR
 					(reg_q113 AND symb_decoder(16#e4#)) OR
 					(reg_q113 AND symb_decoder(16#10#)) OR
 					(reg_q113 AND symb_decoder(16#e3#)) OR
 					(reg_q113 AND symb_decoder(16#24#)) OR
 					(reg_q113 AND symb_decoder(16#42#)) OR
 					(reg_q113 AND symb_decoder(16#b6#)) OR
 					(reg_q113 AND symb_decoder(16#62#)) OR
 					(reg_q113 AND symb_decoder(16#3b#)) OR
 					(reg_q113 AND symb_decoder(16#1b#)) OR
 					(reg_q113 AND symb_decoder(16#cc#)) OR
 					(reg_q113 AND symb_decoder(16#86#)) OR
 					(reg_q113 AND symb_decoder(16#9d#)) OR
 					(reg_q113 AND symb_decoder(16#b1#)) OR
 					(reg_q113 AND symb_decoder(16#07#)) OR
 					(reg_q113 AND symb_decoder(16#fb#)) OR
 					(reg_q113 AND symb_decoder(16#a8#)) OR
 					(reg_q113 AND symb_decoder(16#4f#)) OR
 					(reg_q113 AND symb_decoder(16#12#)) OR
 					(reg_q113 AND symb_decoder(16#c9#)) OR
 					(reg_q113 AND symb_decoder(16#ec#)) OR
 					(reg_q113 AND symb_decoder(16#b7#)) OR
 					(reg_q113 AND symb_decoder(16#d3#)) OR
 					(reg_q113 AND symb_decoder(16#22#)) OR
 					(reg_q113 AND symb_decoder(16#7f#)) OR
 					(reg_q113 AND symb_decoder(16#d0#)) OR
 					(reg_q113 AND symb_decoder(16#ad#)) OR
 					(reg_q113 AND symb_decoder(16#89#)) OR
 					(reg_q113 AND symb_decoder(16#56#)) OR
 					(reg_q113 AND symb_decoder(16#e9#)) OR
 					(reg_q113 AND symb_decoder(16#11#)) OR
 					(reg_q113 AND symb_decoder(16#ce#)) OR
 					(reg_q113 AND symb_decoder(16#e0#)) OR
 					(reg_q113 AND symb_decoder(16#08#));
reg_q498_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q497 AND symb_decoder(16#0d#)) OR
 					(reg_q497 AND symb_decoder(16#0a#));
reg_fullgraph62_init <= "00";

reg_fullgraph62_sel <= "00" & reg_q498_in & reg_q113_in;

	--coder fullgraph62
with reg_fullgraph62_sel select
reg_fullgraph62_in <=
	"01" when "0001",
	"10" when "0010",
	"00" when others;
 --end coder

	p_reg_fullgraph62: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph62 <= reg_fullgraph62_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph62 <= reg_fullgraph62_init;
        else
          reg_fullgraph62 <= reg_fullgraph62_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph62

		reg_q113 <= '1' when reg_fullgraph62 = "01" else '0'; 
		reg_q498 <= '1' when reg_fullgraph62 = "10" else '0'; 
--end decoder 

reg_q116_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q116 AND symb_decoder(16#16#)) OR
 					(reg_q116 AND symb_decoder(16#93#)) OR
 					(reg_q116 AND symb_decoder(16#4b#)) OR
 					(reg_q116 AND symb_decoder(16#9e#)) OR
 					(reg_q116 AND symb_decoder(16#03#)) OR
 					(reg_q116 AND symb_decoder(16#f1#)) OR
 					(reg_q116 AND symb_decoder(16#ca#)) OR
 					(reg_q116 AND symb_decoder(16#9a#)) OR
 					(reg_q116 AND symb_decoder(16#22#)) OR
 					(reg_q116 AND symb_decoder(16#46#)) OR
 					(reg_q116 AND symb_decoder(16#cd#)) OR
 					(reg_q116 AND symb_decoder(16#71#)) OR
 					(reg_q116 AND symb_decoder(16#6d#)) OR
 					(reg_q116 AND symb_decoder(16#14#)) OR
 					(reg_q116 AND symb_decoder(16#31#)) OR
 					(reg_q116 AND symb_decoder(16#0a#)) OR
 					(reg_q116 AND symb_decoder(16#27#)) OR
 					(reg_q116 AND symb_decoder(16#05#)) OR
 					(reg_q116 AND symb_decoder(16#59#)) OR
 					(reg_q116 AND symb_decoder(16#88#)) OR
 					(reg_q116 AND symb_decoder(16#1f#)) OR
 					(reg_q116 AND symb_decoder(16#c7#)) OR
 					(reg_q116 AND symb_decoder(16#d5#)) OR
 					(reg_q116 AND symb_decoder(16#aa#)) OR
 					(reg_q116 AND symb_decoder(16#8e#)) OR
 					(reg_q116 AND symb_decoder(16#df#)) OR
 					(reg_q116 AND symb_decoder(16#42#)) OR
 					(reg_q116 AND symb_decoder(16#b0#)) OR
 					(reg_q116 AND symb_decoder(16#19#)) OR
 					(reg_q116 AND symb_decoder(16#32#)) OR
 					(reg_q116 AND symb_decoder(16#4d#)) OR
 					(reg_q116 AND symb_decoder(16#55#)) OR
 					(reg_q116 AND symb_decoder(16#8d#)) OR
 					(reg_q116 AND symb_decoder(16#3b#)) OR
 					(reg_q116 AND symb_decoder(16#e2#)) OR
 					(reg_q116 AND symb_decoder(16#76#)) OR
 					(reg_q116 AND symb_decoder(16#a6#)) OR
 					(reg_q116 AND symb_decoder(16#e0#)) OR
 					(reg_q116 AND symb_decoder(16#63#)) OR
 					(reg_q116 AND symb_decoder(16#35#)) OR
 					(reg_q116 AND symb_decoder(16#b2#)) OR
 					(reg_q116 AND symb_decoder(16#fe#)) OR
 					(reg_q116 AND symb_decoder(16#74#)) OR
 					(reg_q116 AND symb_decoder(16#9c#)) OR
 					(reg_q116 AND symb_decoder(16#e3#)) OR
 					(reg_q116 AND symb_decoder(16#f9#)) OR
 					(reg_q116 AND symb_decoder(16#92#)) OR
 					(reg_q116 AND symb_decoder(16#5c#)) OR
 					(reg_q116 AND symb_decoder(16#dc#)) OR
 					(reg_q116 AND symb_decoder(16#5d#)) OR
 					(reg_q116 AND symb_decoder(16#13#)) OR
 					(reg_q116 AND symb_decoder(16#c5#)) OR
 					(reg_q116 AND symb_decoder(16#4f#)) OR
 					(reg_q116 AND symb_decoder(16#1e#)) OR
 					(reg_q116 AND symb_decoder(16#0f#)) OR
 					(reg_q116 AND symb_decoder(16#67#)) OR
 					(reg_q116 AND symb_decoder(16#c1#)) OR
 					(reg_q116 AND symb_decoder(16#20#)) OR
 					(reg_q116 AND symb_decoder(16#ec#)) OR
 					(reg_q116 AND symb_decoder(16#f5#)) OR
 					(reg_q116 AND symb_decoder(16#d3#)) OR
 					(reg_q116 AND symb_decoder(16#f8#)) OR
 					(reg_q116 AND symb_decoder(16#0e#)) OR
 					(reg_q116 AND symb_decoder(16#8b#)) OR
 					(reg_q116 AND symb_decoder(16#40#)) OR
 					(reg_q116 AND symb_decoder(16#07#)) OR
 					(reg_q116 AND symb_decoder(16#ee#)) OR
 					(reg_q116 AND symb_decoder(16#6c#)) OR
 					(reg_q116 AND symb_decoder(16#bb#)) OR
 					(reg_q116 AND symb_decoder(16#e5#)) OR
 					(reg_q116 AND symb_decoder(16#69#)) OR
 					(reg_q116 AND symb_decoder(16#6a#)) OR
 					(reg_q116 AND symb_decoder(16#5e#)) OR
 					(reg_q116 AND symb_decoder(16#70#)) OR
 					(reg_q116 AND symb_decoder(16#95#)) OR
 					(reg_q116 AND symb_decoder(16#c3#)) OR
 					(reg_q116 AND symb_decoder(16#7e#)) OR
 					(reg_q116 AND symb_decoder(16#f6#)) OR
 					(reg_q116 AND symb_decoder(16#73#)) OR
 					(reg_q116 AND symb_decoder(16#e4#)) OR
 					(reg_q116 AND symb_decoder(16#7c#)) OR
 					(reg_q116 AND symb_decoder(16#79#)) OR
 					(reg_q116 AND symb_decoder(16#cb#)) OR
 					(reg_q116 AND symb_decoder(16#12#)) OR
 					(reg_q116 AND symb_decoder(16#3a#)) OR
 					(reg_q116 AND symb_decoder(16#d6#)) OR
 					(reg_q116 AND symb_decoder(16#41#)) OR
 					(reg_q116 AND symb_decoder(16#34#)) OR
 					(reg_q116 AND symb_decoder(16#39#)) OR
 					(reg_q116 AND symb_decoder(16#7a#)) OR
 					(reg_q116 AND symb_decoder(16#2b#)) OR
 					(reg_q116 AND symb_decoder(16#a0#)) OR
 					(reg_q116 AND symb_decoder(16#2a#)) OR
 					(reg_q116 AND symb_decoder(16#a7#)) OR
 					(reg_q116 AND symb_decoder(16#57#)) OR
 					(reg_q116 AND symb_decoder(16#d0#)) OR
 					(reg_q116 AND symb_decoder(16#00#)) OR
 					(reg_q116 AND symb_decoder(16#62#)) OR
 					(reg_q116 AND symb_decoder(16#fc#)) OR
 					(reg_q116 AND symb_decoder(16#c2#)) OR
 					(reg_q116 AND symb_decoder(16#43#)) OR
 					(reg_q116 AND symb_decoder(16#7d#)) OR
 					(reg_q116 AND symb_decoder(16#82#)) OR
 					(reg_q116 AND symb_decoder(16#30#)) OR
 					(reg_q116 AND symb_decoder(16#a1#)) OR
 					(reg_q116 AND symb_decoder(16#18#)) OR
 					(reg_q116 AND symb_decoder(16#50#)) OR
 					(reg_q116 AND symb_decoder(16#a3#)) OR
 					(reg_q116 AND symb_decoder(16#29#)) OR
 					(reg_q116 AND symb_decoder(16#26#)) OR
 					(reg_q116 AND symb_decoder(16#a5#)) OR
 					(reg_q116 AND symb_decoder(16#77#)) OR
 					(reg_q116 AND symb_decoder(16#3e#)) OR
 					(reg_q116 AND symb_decoder(16#47#)) OR
 					(reg_q116 AND symb_decoder(16#b4#)) OR
 					(reg_q116 AND symb_decoder(16#fb#)) OR
 					(reg_q116 AND symb_decoder(16#bf#)) OR
 					(reg_q116 AND symb_decoder(16#e6#)) OR
 					(reg_q116 AND symb_decoder(16#a2#)) OR
 					(reg_q116 AND symb_decoder(16#24#)) OR
 					(reg_q116 AND symb_decoder(16#65#)) OR
 					(reg_q116 AND symb_decoder(16#10#)) OR
 					(reg_q116 AND symb_decoder(16#c8#)) OR
 					(reg_q116 AND symb_decoder(16#fa#)) OR
 					(reg_q116 AND symb_decoder(16#d8#)) OR
 					(reg_q116 AND symb_decoder(16#64#)) OR
 					(reg_q116 AND symb_decoder(16#fd#)) OR
 					(reg_q116 AND symb_decoder(16#ce#)) OR
 					(reg_q116 AND symb_decoder(16#84#)) OR
 					(reg_q116 AND symb_decoder(16#2f#)) OR
 					(reg_q116 AND symb_decoder(16#8a#)) OR
 					(reg_q116 AND symb_decoder(16#61#)) OR
 					(reg_q116 AND symb_decoder(16#ed#)) OR
 					(reg_q116 AND symb_decoder(16#6e#)) OR
 					(reg_q116 AND symb_decoder(16#72#)) OR
 					(reg_q116 AND symb_decoder(16#dd#)) OR
 					(reg_q116 AND symb_decoder(16#3c#)) OR
 					(reg_q116 AND symb_decoder(16#44#)) OR
 					(reg_q116 AND symb_decoder(16#c6#)) OR
 					(reg_q116 AND symb_decoder(16#6b#)) OR
 					(reg_q116 AND symb_decoder(16#01#)) OR
 					(reg_q116 AND symb_decoder(16#08#)) OR
 					(reg_q116 AND symb_decoder(16#ab#)) OR
 					(reg_q116 AND symb_decoder(16#75#)) OR
 					(reg_q116 AND symb_decoder(16#cf#)) OR
 					(reg_q116 AND symb_decoder(16#f3#)) OR
 					(reg_q116 AND symb_decoder(16#1d#)) OR
 					(reg_q116 AND symb_decoder(16#b6#)) OR
 					(reg_q116 AND symb_decoder(16#ac#)) OR
 					(reg_q116 AND symb_decoder(16#04#)) OR
 					(reg_q116 AND symb_decoder(16#d1#)) OR
 					(reg_q116 AND symb_decoder(16#5b#)) OR
 					(reg_q116 AND symb_decoder(16#d9#)) OR
 					(reg_q116 AND symb_decoder(16#56#)) OR
 					(reg_q116 AND symb_decoder(16#ae#)) OR
 					(reg_q116 AND symb_decoder(16#09#)) OR
 					(reg_q116 AND symb_decoder(16#11#)) OR
 					(reg_q116 AND symb_decoder(16#89#)) OR
 					(reg_q116 AND symb_decoder(16#85#)) OR
 					(reg_q116 AND symb_decoder(16#ad#)) OR
 					(reg_q116 AND symb_decoder(16#ba#)) OR
 					(reg_q116 AND symb_decoder(16#78#)) OR
 					(reg_q116 AND symb_decoder(16#94#)) OR
 					(reg_q116 AND symb_decoder(16#4e#)) OR
 					(reg_q116 AND symb_decoder(16#c0#)) OR
 					(reg_q116 AND symb_decoder(16#17#)) OR
 					(reg_q116 AND symb_decoder(16#1c#)) OR
 					(reg_q116 AND symb_decoder(16#81#)) OR
 					(reg_q116 AND symb_decoder(16#cc#)) OR
 					(reg_q116 AND symb_decoder(16#c4#)) OR
 					(reg_q116 AND symb_decoder(16#bc#)) OR
 					(reg_q116 AND symb_decoder(16#5f#)) OR
 					(reg_q116 AND symb_decoder(16#eb#)) OR
 					(reg_q116 AND symb_decoder(16#23#)) OR
 					(reg_q116 AND symb_decoder(16#80#)) OR
 					(reg_q116 AND symb_decoder(16#9d#)) OR
 					(reg_q116 AND symb_decoder(16#60#)) OR
 					(reg_q116 AND symb_decoder(16#b9#)) OR
 					(reg_q116 AND symb_decoder(16#d2#)) OR
 					(reg_q116 AND symb_decoder(16#a9#)) OR
 					(reg_q116 AND symb_decoder(16#a8#)) OR
 					(reg_q116 AND symb_decoder(16#e1#)) OR
 					(reg_q116 AND symb_decoder(16#06#)) OR
 					(reg_q116 AND symb_decoder(16#a4#)) OR
 					(reg_q116 AND symb_decoder(16#0c#)) OR
 					(reg_q116 AND symb_decoder(16#86#)) OR
 					(reg_q116 AND symb_decoder(16#97#)) OR
 					(reg_q116 AND symb_decoder(16#48#)) OR
 					(reg_q116 AND symb_decoder(16#21#)) OR
 					(reg_q116 AND symb_decoder(16#af#)) OR
 					(reg_q116 AND symb_decoder(16#02#)) OR
 					(reg_q116 AND symb_decoder(16#52#)) OR
 					(reg_q116 AND symb_decoder(16#b7#)) OR
 					(reg_q116 AND symb_decoder(16#54#)) OR
 					(reg_q116 AND symb_decoder(16#91#)) OR
 					(reg_q116 AND symb_decoder(16#da#)) OR
 					(reg_q116 AND symb_decoder(16#2c#)) OR
 					(reg_q116 AND symb_decoder(16#58#)) OR
 					(reg_q116 AND symb_decoder(16#f0#)) OR
 					(reg_q116 AND symb_decoder(16#b1#)) OR
 					(reg_q116 AND symb_decoder(16#b3#)) OR
 					(reg_q116 AND symb_decoder(16#68#)) OR
 					(reg_q116 AND symb_decoder(16#96#)) OR
 					(reg_q116 AND symb_decoder(16#51#)) OR
 					(reg_q116 AND symb_decoder(16#99#)) OR
 					(reg_q116 AND symb_decoder(16#2d#)) OR
 					(reg_q116 AND symb_decoder(16#83#)) OR
 					(reg_q116 AND symb_decoder(16#36#)) OR
 					(reg_q116 AND symb_decoder(16#66#)) OR
 					(reg_q116 AND symb_decoder(16#b5#)) OR
 					(reg_q116 AND symb_decoder(16#8c#)) OR
 					(reg_q116 AND symb_decoder(16#87#)) OR
 					(reg_q116 AND symb_decoder(16#b8#)) OR
 					(reg_q116 AND symb_decoder(16#4a#)) OR
 					(reg_q116 AND symb_decoder(16#7f#)) OR
 					(reg_q116 AND symb_decoder(16#25#)) OR
 					(reg_q116 AND symb_decoder(16#0b#)) OR
 					(reg_q116 AND symb_decoder(16#49#)) OR
 					(reg_q116 AND symb_decoder(16#53#)) OR
 					(reg_q116 AND symb_decoder(16#28#)) OR
 					(reg_q116 AND symb_decoder(16#6f#)) OR
 					(reg_q116 AND symb_decoder(16#db#)) OR
 					(reg_q116 AND symb_decoder(16#ef#)) OR
 					(reg_q116 AND symb_decoder(16#7b#)) OR
 					(reg_q116 AND symb_decoder(16#f2#)) OR
 					(reg_q116 AND symb_decoder(16#3d#)) OR
 					(reg_q116 AND symb_decoder(16#0d#)) OR
 					(reg_q116 AND symb_decoder(16#45#)) OR
 					(reg_q116 AND symb_decoder(16#3f#)) OR
 					(reg_q116 AND symb_decoder(16#be#)) OR
 					(reg_q116 AND symb_decoder(16#9b#)) OR
 					(reg_q116 AND symb_decoder(16#ff#)) OR
 					(reg_q116 AND symb_decoder(16#c9#)) OR
 					(reg_q116 AND symb_decoder(16#1a#)) OR
 					(reg_q116 AND symb_decoder(16#90#)) OR
 					(reg_q116 AND symb_decoder(16#e9#)) OR
 					(reg_q116 AND symb_decoder(16#de#)) OR
 					(reg_q116 AND symb_decoder(16#2e#)) OR
 					(reg_q116 AND symb_decoder(16#bd#)) OR
 					(reg_q116 AND symb_decoder(16#f4#)) OR
 					(reg_q116 AND symb_decoder(16#e7#)) OR
 					(reg_q116 AND symb_decoder(16#f7#)) OR
 					(reg_q116 AND symb_decoder(16#37#)) OR
 					(reg_q116 AND symb_decoder(16#1b#)) OR
 					(reg_q116 AND symb_decoder(16#38#)) OR
 					(reg_q116 AND symb_decoder(16#33#)) OR
 					(reg_q116 AND symb_decoder(16#98#)) OR
 					(reg_q116 AND symb_decoder(16#e8#)) OR
 					(reg_q116 AND symb_decoder(16#4c#)) OR
 					(reg_q116 AND symb_decoder(16#15#)) OR
 					(reg_q116 AND symb_decoder(16#ea#)) OR
 					(reg_q116 AND symb_decoder(16#8f#)) OR
 					(reg_q116 AND symb_decoder(16#9f#)) OR
 					(reg_q116 AND symb_decoder(16#5a#)) OR
 					(reg_q116 AND symb_decoder(16#d4#)) OR
 					(reg_q116 AND symb_decoder(16#d7#));
reg_q116_init <= '0' ;
	p_reg_q116: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q116 <= reg_q116_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q116 <= reg_q116_init;
        else
          reg_q116 <= reg_q116_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph64

reg_q2326_in <= (reg_q2290 AND symb_decoder(16#10#)) OR
 					(reg_q2290 AND symb_decoder(16#1e#)) OR
 					(reg_q2290 AND symb_decoder(16#f8#)) OR
 					(reg_q2290 AND symb_decoder(16#1f#)) OR
 					(reg_q2290 AND symb_decoder(16#36#)) OR
 					(reg_q2290 AND symb_decoder(16#67#)) OR
 					(reg_q2290 AND symb_decoder(16#c8#)) OR
 					(reg_q2290 AND symb_decoder(16#f4#)) OR
 					(reg_q2290 AND symb_decoder(16#49#)) OR
 					(reg_q2290 AND symb_decoder(16#97#)) OR
 					(reg_q2290 AND symb_decoder(16#64#)) OR
 					(reg_q2290 AND symb_decoder(16#a7#)) OR
 					(reg_q2290 AND symb_decoder(16#cb#)) OR
 					(reg_q2290 AND symb_decoder(16#04#)) OR
 					(reg_q2290 AND symb_decoder(16#ae#)) OR
 					(reg_q2290 AND symb_decoder(16#e5#)) OR
 					(reg_q2290 AND symb_decoder(16#57#)) OR
 					(reg_q2290 AND symb_decoder(16#54#)) OR
 					(reg_q2290 AND symb_decoder(16#be#)) OR
 					(reg_q2290 AND symb_decoder(16#1d#)) OR
 					(reg_q2290 AND symb_decoder(16#b8#)) OR
 					(reg_q2290 AND symb_decoder(16#e6#)) OR
 					(reg_q2290 AND symb_decoder(16#c1#)) OR
 					(reg_q2290 AND symb_decoder(16#a5#)) OR
 					(reg_q2290 AND symb_decoder(16#8e#)) OR
 					(reg_q2290 AND symb_decoder(16#e1#)) OR
 					(reg_q2290 AND symb_decoder(16#bb#)) OR
 					(reg_q2290 AND symb_decoder(16#e9#)) OR
 					(reg_q2290 AND symb_decoder(16#8a#)) OR
 					(reg_q2290 AND symb_decoder(16#98#)) OR
 					(reg_q2290 AND symb_decoder(16#a0#)) OR
 					(reg_q2290 AND symb_decoder(16#94#)) OR
 					(reg_q2290 AND symb_decoder(16#00#)) OR
 					(reg_q2290 AND symb_decoder(16#9c#)) OR
 					(reg_q2290 AND symb_decoder(16#66#)) OR
 					(reg_q2290 AND symb_decoder(16#4b#)) OR
 					(reg_q2290 AND symb_decoder(16#ca#)) OR
 					(reg_q2290 AND symb_decoder(16#d2#)) OR
 					(reg_q2290 AND symb_decoder(16#2f#)) OR
 					(reg_q2290 AND symb_decoder(16#e2#)) OR
 					(reg_q2290 AND symb_decoder(16#6f#)) OR
 					(reg_q2290 AND symb_decoder(16#ea#)) OR
 					(reg_q2290 AND symb_decoder(16#86#)) OR
 					(reg_q2290 AND symb_decoder(16#ad#)) OR
 					(reg_q2290 AND symb_decoder(16#50#)) OR
 					(reg_q2290 AND symb_decoder(16#c7#)) OR
 					(reg_q2290 AND symb_decoder(16#32#)) OR
 					(reg_q2290 AND symb_decoder(16#44#)) OR
 					(reg_q2290 AND symb_decoder(16#ce#)) OR
 					(reg_q2290 AND symb_decoder(16#0c#)) OR
 					(reg_q2290 AND symb_decoder(16#11#)) OR
 					(reg_q2290 AND symb_decoder(16#39#)) OR
 					(reg_q2290 AND symb_decoder(16#2e#)) OR
 					(reg_q2290 AND symb_decoder(16#6c#)) OR
 					(reg_q2290 AND symb_decoder(16#28#)) OR
 					(reg_q2290 AND symb_decoder(16#12#)) OR
 					(reg_q2290 AND symb_decoder(16#9e#)) OR
 					(reg_q2290 AND symb_decoder(16#2a#)) OR
 					(reg_q2290 AND symb_decoder(16#60#)) OR
 					(reg_q2290 AND symb_decoder(16#15#)) OR
 					(reg_q2290 AND symb_decoder(16#68#)) OR
 					(reg_q2290 AND symb_decoder(16#aa#)) OR
 					(reg_q2290 AND symb_decoder(16#70#)) OR
 					(reg_q2290 AND symb_decoder(16#31#)) OR
 					(reg_q2290 AND symb_decoder(16#0b#)) OR
 					(reg_q2290 AND symb_decoder(16#fa#)) OR
 					(reg_q2290 AND symb_decoder(16#47#)) OR
 					(reg_q2290 AND symb_decoder(16#0f#)) OR
 					(reg_q2290 AND symb_decoder(16#85#)) OR
 					(reg_q2290 AND symb_decoder(16#06#)) OR
 					(reg_q2290 AND symb_decoder(16#a6#)) OR
 					(reg_q2290 AND symb_decoder(16#a2#)) OR
 					(reg_q2290 AND symb_decoder(16#20#)) OR
 					(reg_q2290 AND symb_decoder(16#cc#)) OR
 					(reg_q2290 AND symb_decoder(16#a9#)) OR
 					(reg_q2290 AND symb_decoder(16#a3#)) OR
 					(reg_q2290 AND symb_decoder(16#83#)) OR
 					(reg_q2290 AND symb_decoder(16#76#)) OR
 					(reg_q2290 AND symb_decoder(16#51#)) OR
 					(reg_q2290 AND symb_decoder(16#d3#)) OR
 					(reg_q2290 AND symb_decoder(16#41#)) OR
 					(reg_q2290 AND symb_decoder(16#d6#)) OR
 					(reg_q2290 AND symb_decoder(16#d7#)) OR
 					(reg_q2290 AND symb_decoder(16#d5#)) OR
 					(reg_q2290 AND symb_decoder(16#13#)) OR
 					(reg_q2290 AND symb_decoder(16#22#)) OR
 					(reg_q2290 AND symb_decoder(16#27#)) OR
 					(reg_q2290 AND symb_decoder(16#05#)) OR
 					(reg_q2290 AND symb_decoder(16#b6#)) OR
 					(reg_q2290 AND symb_decoder(16#55#)) OR
 					(reg_q2290 AND symb_decoder(16#e4#)) OR
 					(reg_q2290 AND symb_decoder(16#35#)) OR
 					(reg_q2290 AND symb_decoder(16#88#)) OR
 					(reg_q2290 AND symb_decoder(16#df#)) OR
 					(reg_q2290 AND symb_decoder(16#87#)) OR
 					(reg_q2290 AND symb_decoder(16#9b#)) OR
 					(reg_q2290 AND symb_decoder(16#fc#)) OR
 					(reg_q2290 AND symb_decoder(16#7e#)) OR
 					(reg_q2290 AND symb_decoder(16#c9#)) OR
 					(reg_q2290 AND symb_decoder(16#93#)) OR
 					(reg_q2290 AND symb_decoder(16#8d#)) OR
 					(reg_q2290 AND symb_decoder(16#cd#)) OR
 					(reg_q2290 AND symb_decoder(16#cf#)) OR
 					(reg_q2290 AND symb_decoder(16#24#)) OR
 					(reg_q2290 AND symb_decoder(16#7f#)) OR
 					(reg_q2290 AND symb_decoder(16#4d#)) OR
 					(reg_q2290 AND symb_decoder(16#1c#)) OR
 					(reg_q2290 AND symb_decoder(16#b9#)) OR
 					(reg_q2290 AND symb_decoder(16#da#)) OR
 					(reg_q2290 AND symb_decoder(16#4f#)) OR
 					(reg_q2290 AND symb_decoder(16#25#)) OR
 					(reg_q2290 AND symb_decoder(16#6a#)) OR
 					(reg_q2290 AND symb_decoder(16#07#)) OR
 					(reg_q2290 AND symb_decoder(16#fd#)) OR
 					(reg_q2290 AND symb_decoder(16#26#)) OR
 					(reg_q2290 AND symb_decoder(16#5c#)) OR
 					(reg_q2290 AND symb_decoder(16#ab#)) OR
 					(reg_q2290 AND symb_decoder(16#e7#)) OR
 					(reg_q2290 AND symb_decoder(16#b2#)) OR
 					(reg_q2290 AND symb_decoder(16#95#)) OR
 					(reg_q2290 AND symb_decoder(16#dd#)) OR
 					(reg_q2290 AND symb_decoder(16#d1#)) OR
 					(reg_q2290 AND symb_decoder(16#a8#)) OR
 					(reg_q2290 AND symb_decoder(16#eb#)) OR
 					(reg_q2290 AND symb_decoder(16#a1#)) OR
 					(reg_q2290 AND symb_decoder(16#3a#)) OR
 					(reg_q2290 AND symb_decoder(16#ef#)) OR
 					(reg_q2290 AND symb_decoder(16#77#)) OR
 					(reg_q2290 AND symb_decoder(16#ee#)) OR
 					(reg_q2290 AND symb_decoder(16#b1#)) OR
 					(reg_q2290 AND symb_decoder(16#37#)) OR
 					(reg_q2290 AND symb_decoder(16#4e#)) OR
 					(reg_q2290 AND symb_decoder(16#38#)) OR
 					(reg_q2290 AND symb_decoder(16#61#)) OR
 					(reg_q2290 AND symb_decoder(16#f7#)) OR
 					(reg_q2290 AND symb_decoder(16#3c#)) OR
 					(reg_q2290 AND symb_decoder(16#82#)) OR
 					(reg_q2290 AND symb_decoder(16#2c#)) OR
 					(reg_q2290 AND symb_decoder(16#53#)) OR
 					(reg_q2290 AND symb_decoder(16#17#)) OR
 					(reg_q2290 AND symb_decoder(16#09#)) OR
 					(reg_q2290 AND symb_decoder(16#7a#)) OR
 					(reg_q2290 AND symb_decoder(16#99#)) OR
 					(reg_q2290 AND symb_decoder(16#8b#)) OR
 					(reg_q2290 AND symb_decoder(16#21#)) OR
 					(reg_q2290 AND symb_decoder(16#5a#)) OR
 					(reg_q2290 AND symb_decoder(16#0e#)) OR
 					(reg_q2290 AND symb_decoder(16#16#)) OR
 					(reg_q2290 AND symb_decoder(16#fb#)) OR
 					(reg_q2290 AND symb_decoder(16#02#)) OR
 					(reg_q2290 AND symb_decoder(16#b7#)) OR
 					(reg_q2290 AND symb_decoder(16#75#)) OR
 					(reg_q2290 AND symb_decoder(16#45#)) OR
 					(reg_q2290 AND symb_decoder(16#29#)) OR
 					(reg_q2290 AND symb_decoder(16#bf#)) OR
 					(reg_q2290 AND symb_decoder(16#01#)) OR
 					(reg_q2290 AND symb_decoder(16#1a#)) OR
 					(reg_q2290 AND symb_decoder(16#af#)) OR
 					(reg_q2290 AND symb_decoder(16#84#)) OR
 					(reg_q2290 AND symb_decoder(16#7b#)) OR
 					(reg_q2290 AND symb_decoder(16#f5#)) OR
 					(reg_q2290 AND symb_decoder(16#4a#)) OR
 					(reg_q2290 AND symb_decoder(16#bc#)) OR
 					(reg_q2290 AND symb_decoder(16#59#)) OR
 					(reg_q2290 AND symb_decoder(16#2b#)) OR
 					(reg_q2290 AND symb_decoder(16#72#)) OR
 					(reg_q2290 AND symb_decoder(16#80#)) OR
 					(reg_q2290 AND symb_decoder(16#23#)) OR
 					(reg_q2290 AND symb_decoder(16#db#)) OR
 					(reg_q2290 AND symb_decoder(16#08#)) OR
 					(reg_q2290 AND symb_decoder(16#81#)) OR
 					(reg_q2290 AND symb_decoder(16#f0#)) OR
 					(reg_q2290 AND symb_decoder(16#92#)) OR
 					(reg_q2290 AND symb_decoder(16#74#)) OR
 					(reg_q2290 AND symb_decoder(16#3e#)) OR
 					(reg_q2290 AND symb_decoder(16#8f#)) OR
 					(reg_q2290 AND symb_decoder(16#73#)) OR
 					(reg_q2290 AND symb_decoder(16#03#)) OR
 					(reg_q2290 AND symb_decoder(16#d0#)) OR
 					(reg_q2290 AND symb_decoder(16#ac#)) OR
 					(reg_q2290 AND symb_decoder(16#bd#)) OR
 					(reg_q2290 AND symb_decoder(16#6b#)) OR
 					(reg_q2290 AND symb_decoder(16#46#)) OR
 					(reg_q2290 AND symb_decoder(16#5e#)) OR
 					(reg_q2290 AND symb_decoder(16#18#)) OR
 					(reg_q2290 AND symb_decoder(16#5d#)) OR
 					(reg_q2290 AND symb_decoder(16#c0#)) OR
 					(reg_q2290 AND symb_decoder(16#9d#)) OR
 					(reg_q2290 AND symb_decoder(16#f1#)) OR
 					(reg_q2290 AND symb_decoder(16#8c#)) OR
 					(reg_q2290 AND symb_decoder(16#ba#)) OR
 					(reg_q2290 AND symb_decoder(16#f2#)) OR
 					(reg_q2290 AND symb_decoder(16#3b#)) OR
 					(reg_q2290 AND symb_decoder(16#fe#)) OR
 					(reg_q2290 AND symb_decoder(16#dc#)) OR
 					(reg_q2290 AND symb_decoder(16#1b#)) OR
 					(reg_q2290 AND symb_decoder(16#91#)) OR
 					(reg_q2290 AND symb_decoder(16#69#)) OR
 					(reg_q2290 AND symb_decoder(16#30#)) OR
 					(reg_q2290 AND symb_decoder(16#c5#)) OR
 					(reg_q2290 AND symb_decoder(16#89#)) OR
 					(reg_q2290 AND symb_decoder(16#ec#)) OR
 					(reg_q2290 AND symb_decoder(16#9f#)) OR
 					(reg_q2290 AND symb_decoder(16#d9#)) OR
 					(reg_q2290 AND symb_decoder(16#14#)) OR
 					(reg_q2290 AND symb_decoder(16#71#)) OR
 					(reg_q2290 AND symb_decoder(16#e3#)) OR
 					(reg_q2290 AND symb_decoder(16#6e#)) OR
 					(reg_q2290 AND symb_decoder(16#65#)) OR
 					(reg_q2290 AND symb_decoder(16#f3#)) OR
 					(reg_q2290 AND symb_decoder(16#b3#)) OR
 					(reg_q2290 AND symb_decoder(16#d8#)) OR
 					(reg_q2290 AND symb_decoder(16#c3#)) OR
 					(reg_q2290 AND symb_decoder(16#6d#)) OR
 					(reg_q2290 AND symb_decoder(16#33#)) OR
 					(reg_q2290 AND symb_decoder(16#40#)) OR
 					(reg_q2290 AND symb_decoder(16#42#)) OR
 					(reg_q2290 AND symb_decoder(16#56#)) OR
 					(reg_q2290 AND symb_decoder(16#5f#)) OR
 					(reg_q2290 AND symb_decoder(16#f9#)) OR
 					(reg_q2290 AND symb_decoder(16#62#)) OR
 					(reg_q2290 AND symb_decoder(16#ff#)) OR
 					(reg_q2290 AND symb_decoder(16#a4#)) OR
 					(reg_q2290 AND symb_decoder(16#3d#)) OR
 					(reg_q2290 AND symb_decoder(16#7c#)) OR
 					(reg_q2290 AND symb_decoder(16#52#)) OR
 					(reg_q2290 AND symb_decoder(16#de#)) OR
 					(reg_q2290 AND symb_decoder(16#4c#)) OR
 					(reg_q2290 AND symb_decoder(16#34#)) OR
 					(reg_q2290 AND symb_decoder(16#c6#)) OR
 					(reg_q2290 AND symb_decoder(16#78#)) OR
 					(reg_q2290 AND symb_decoder(16#e0#)) OR
 					(reg_q2290 AND symb_decoder(16#b4#)) OR
 					(reg_q2290 AND symb_decoder(16#ed#)) OR
 					(reg_q2290 AND symb_decoder(16#5b#)) OR
 					(reg_q2290 AND symb_decoder(16#d4#)) OR
 					(reg_q2290 AND symb_decoder(16#f6#)) OR
 					(reg_q2290 AND symb_decoder(16#58#)) OR
 					(reg_q2290 AND symb_decoder(16#43#)) OR
 					(reg_q2290 AND symb_decoder(16#7d#)) OR
 					(reg_q2290 AND symb_decoder(16#79#)) OR
 					(reg_q2290 AND symb_decoder(16#c2#)) OR
 					(reg_q2290 AND symb_decoder(16#19#)) OR
 					(reg_q2290 AND symb_decoder(16#63#)) OR
 					(reg_q2290 AND symb_decoder(16#b5#)) OR
 					(reg_q2290 AND symb_decoder(16#c4#)) OR
 					(reg_q2290 AND symb_decoder(16#2d#)) OR
 					(reg_q2290 AND symb_decoder(16#b0#)) OR
 					(reg_q2290 AND symb_decoder(16#e8#)) OR
 					(reg_q2290 AND symb_decoder(16#96#)) OR
 					(reg_q2290 AND symb_decoder(16#48#)) OR
 					(reg_q2290 AND symb_decoder(16#90#)) OR
 					(reg_q2290 AND symb_decoder(16#3f#)) OR
 					(reg_q2290 AND symb_decoder(16#9a#)) OR
 					(reg_q2326 AND symb_decoder(16#5f#)) OR
 					(reg_q2326 AND symb_decoder(16#65#)) OR
 					(reg_q2326 AND symb_decoder(16#7f#)) OR
 					(reg_q2326 AND symb_decoder(16#01#)) OR
 					(reg_q2326 AND symb_decoder(16#5d#)) OR
 					(reg_q2326 AND symb_decoder(16#f9#)) OR
 					(reg_q2326 AND symb_decoder(16#5e#)) OR
 					(reg_q2326 AND symb_decoder(16#b4#)) OR
 					(reg_q2326 AND symb_decoder(16#ed#)) OR
 					(reg_q2326 AND symb_decoder(16#93#)) OR
 					(reg_q2326 AND symb_decoder(16#1d#)) OR
 					(reg_q2326 AND symb_decoder(16#b8#)) OR
 					(reg_q2326 AND symb_decoder(16#dd#)) OR
 					(reg_q2326 AND symb_decoder(16#98#)) OR
 					(reg_q2326 AND symb_decoder(16#6b#)) OR
 					(reg_q2326 AND symb_decoder(16#d9#)) OR
 					(reg_q2326 AND symb_decoder(16#fe#)) OR
 					(reg_q2326 AND symb_decoder(16#7d#)) OR
 					(reg_q2326 AND symb_decoder(16#bc#)) OR
 					(reg_q2326 AND symb_decoder(16#47#)) OR
 					(reg_q2326 AND symb_decoder(16#41#)) OR
 					(reg_q2326 AND symb_decoder(16#95#)) OR
 					(reg_q2326 AND symb_decoder(16#51#)) OR
 					(reg_q2326 AND symb_decoder(16#cd#)) OR
 					(reg_q2326 AND symb_decoder(16#92#)) OR
 					(reg_q2326 AND symb_decoder(16#f8#)) OR
 					(reg_q2326 AND symb_decoder(16#a0#)) OR
 					(reg_q2326 AND symb_decoder(16#a1#)) OR
 					(reg_q2326 AND symb_decoder(16#e9#)) OR
 					(reg_q2326 AND symb_decoder(16#91#)) OR
 					(reg_q2326 AND symb_decoder(16#09#)) OR
 					(reg_q2326 AND symb_decoder(16#24#)) OR
 					(reg_q2326 AND symb_decoder(16#3d#)) OR
 					(reg_q2326 AND symb_decoder(16#9e#)) OR
 					(reg_q2326 AND symb_decoder(16#7b#)) OR
 					(reg_q2326 AND symb_decoder(16#ea#)) OR
 					(reg_q2326 AND symb_decoder(16#9a#)) OR
 					(reg_q2326 AND symb_decoder(16#1c#)) OR
 					(reg_q2326 AND symb_decoder(16#67#)) OR
 					(reg_q2326 AND symb_decoder(16#71#)) OR
 					(reg_q2326 AND symb_decoder(16#30#)) OR
 					(reg_q2326 AND symb_decoder(16#b7#)) OR
 					(reg_q2326 AND symb_decoder(16#66#)) OR
 					(reg_q2326 AND symb_decoder(16#4f#)) OR
 					(reg_q2326 AND symb_decoder(16#1f#)) OR
 					(reg_q2326 AND symb_decoder(16#3e#)) OR
 					(reg_q2326 AND symb_decoder(16#b9#)) OR
 					(reg_q2326 AND symb_decoder(16#d7#)) OR
 					(reg_q2326 AND symb_decoder(16#b6#)) OR
 					(reg_q2326 AND symb_decoder(16#86#)) OR
 					(reg_q2326 AND symb_decoder(16#b0#)) OR
 					(reg_q2326 AND symb_decoder(16#db#)) OR
 					(reg_q2326 AND symb_decoder(16#21#)) OR
 					(reg_q2326 AND symb_decoder(16#0f#)) OR
 					(reg_q2326 AND symb_decoder(16#49#)) OR
 					(reg_q2326 AND symb_decoder(16#16#)) OR
 					(reg_q2326 AND symb_decoder(16#55#)) OR
 					(reg_q2326 AND symb_decoder(16#5b#)) OR
 					(reg_q2326 AND symb_decoder(16#34#)) OR
 					(reg_q2326 AND symb_decoder(16#2f#)) OR
 					(reg_q2326 AND symb_decoder(16#14#)) OR
 					(reg_q2326 AND symb_decoder(16#e1#)) OR
 					(reg_q2326 AND symb_decoder(16#52#)) OR
 					(reg_q2326 AND symb_decoder(16#05#)) OR
 					(reg_q2326 AND symb_decoder(16#1e#)) OR
 					(reg_q2326 AND symb_decoder(16#43#)) OR
 					(reg_q2326 AND symb_decoder(16#d0#)) OR
 					(reg_q2326 AND symb_decoder(16#28#)) OR
 					(reg_q2326 AND symb_decoder(16#a8#)) OR
 					(reg_q2326 AND symb_decoder(16#18#)) OR
 					(reg_q2326 AND symb_decoder(16#7a#)) OR
 					(reg_q2326 AND symb_decoder(16#c0#)) OR
 					(reg_q2326 AND symb_decoder(16#f6#)) OR
 					(reg_q2326 AND symb_decoder(16#56#)) OR
 					(reg_q2326 AND symb_decoder(16#17#)) OR
 					(reg_q2326 AND symb_decoder(16#5c#)) OR
 					(reg_q2326 AND symb_decoder(16#80#)) OR
 					(reg_q2326 AND symb_decoder(16#ec#)) OR
 					(reg_q2326 AND symb_decoder(16#33#)) OR
 					(reg_q2326 AND symb_decoder(16#3a#)) OR
 					(reg_q2326 AND symb_decoder(16#0c#)) OR
 					(reg_q2326 AND symb_decoder(16#7c#)) OR
 					(reg_q2326 AND symb_decoder(16#37#)) OR
 					(reg_q2326 AND symb_decoder(16#69#)) OR
 					(reg_q2326 AND symb_decoder(16#f7#)) OR
 					(reg_q2326 AND symb_decoder(16#ef#)) OR
 					(reg_q2326 AND symb_decoder(16#53#)) OR
 					(reg_q2326 AND symb_decoder(16#af#)) OR
 					(reg_q2326 AND symb_decoder(16#97#)) OR
 					(reg_q2326 AND symb_decoder(16#94#)) OR
 					(reg_q2326 AND symb_decoder(16#df#)) OR
 					(reg_q2326 AND symb_decoder(16#d3#)) OR
 					(reg_q2326 AND symb_decoder(16#fa#)) OR
 					(reg_q2326 AND symb_decoder(16#9d#)) OR
 					(reg_q2326 AND symb_decoder(16#88#)) OR
 					(reg_q2326 AND symb_decoder(16#57#)) OR
 					(reg_q2326 AND symb_decoder(16#2c#)) OR
 					(reg_q2326 AND symb_decoder(16#68#)) OR
 					(reg_q2326 AND symb_decoder(16#81#)) OR
 					(reg_q2326 AND symb_decoder(16#62#)) OR
 					(reg_q2326 AND symb_decoder(16#96#)) OR
 					(reg_q2326 AND symb_decoder(16#89#)) OR
 					(reg_q2326 AND symb_decoder(16#03#)) OR
 					(reg_q2326 AND symb_decoder(16#06#)) OR
 					(reg_q2326 AND symb_decoder(16#fb#)) OR
 					(reg_q2326 AND symb_decoder(16#e2#)) OR
 					(reg_q2326 AND symb_decoder(16#c2#)) OR
 					(reg_q2326 AND symb_decoder(16#bd#)) OR
 					(reg_q2326 AND symb_decoder(16#ba#)) OR
 					(reg_q2326 AND symb_decoder(16#f1#)) OR
 					(reg_q2326 AND symb_decoder(16#f5#)) OR
 					(reg_q2326 AND symb_decoder(16#00#)) OR
 					(reg_q2326 AND symb_decoder(16#4a#)) OR
 					(reg_q2326 AND symb_decoder(16#44#)) OR
 					(reg_q2326 AND symb_decoder(16#bf#)) OR
 					(reg_q2326 AND symb_decoder(16#e7#)) OR
 					(reg_q2326 AND symb_decoder(16#e6#)) OR
 					(reg_q2326 AND symb_decoder(16#4b#)) OR
 					(reg_q2326 AND symb_decoder(16#cf#)) OR
 					(reg_q2326 AND symb_decoder(16#e0#)) OR
 					(reg_q2326 AND symb_decoder(16#77#)) OR
 					(reg_q2326 AND symb_decoder(16#a2#)) OR
 					(reg_q2326 AND symb_decoder(16#40#)) OR
 					(reg_q2326 AND symb_decoder(16#74#)) OR
 					(reg_q2326 AND symb_decoder(16#c6#)) OR
 					(reg_q2326 AND symb_decoder(16#83#)) OR
 					(reg_q2326 AND symb_decoder(16#ff#)) OR
 					(reg_q2326 AND symb_decoder(16#72#)) OR
 					(reg_q2326 AND symb_decoder(16#2b#)) OR
 					(reg_q2326 AND symb_decoder(16#8c#)) OR
 					(reg_q2326 AND symb_decoder(16#be#)) OR
 					(reg_q2326 AND symb_decoder(16#9c#)) OR
 					(reg_q2326 AND symb_decoder(16#fc#)) OR
 					(reg_q2326 AND symb_decoder(16#8a#)) OR
 					(reg_q2326 AND symb_decoder(16#f3#)) OR
 					(reg_q2326 AND symb_decoder(16#f2#)) OR
 					(reg_q2326 AND symb_decoder(16#82#)) OR
 					(reg_q2326 AND symb_decoder(16#b3#)) OR
 					(reg_q2326 AND symb_decoder(16#dc#)) OR
 					(reg_q2326 AND symb_decoder(16#35#)) OR
 					(reg_q2326 AND symb_decoder(16#63#)) OR
 					(reg_q2326 AND symb_decoder(16#2d#)) OR
 					(reg_q2326 AND symb_decoder(16#b1#)) OR
 					(reg_q2326 AND symb_decoder(16#ab#)) OR
 					(reg_q2326 AND symb_decoder(16#23#)) OR
 					(reg_q2326 AND symb_decoder(16#04#)) OR
 					(reg_q2326 AND symb_decoder(16#a4#)) OR
 					(reg_q2326 AND symb_decoder(16#76#)) OR
 					(reg_q2326 AND symb_decoder(16#27#)) OR
 					(reg_q2326 AND symb_decoder(16#60#)) OR
 					(reg_q2326 AND symb_decoder(16#de#)) OR
 					(reg_q2326 AND symb_decoder(16#50#)) OR
 					(reg_q2326 AND symb_decoder(16#36#)) OR
 					(reg_q2326 AND symb_decoder(16#c5#)) OR
 					(reg_q2326 AND symb_decoder(16#bb#)) OR
 					(reg_q2326 AND symb_decoder(16#58#)) OR
 					(reg_q2326 AND symb_decoder(16#6e#)) OR
 					(reg_q2326 AND symb_decoder(16#d5#)) OR
 					(reg_q2326 AND symb_decoder(16#5a#)) OR
 					(reg_q2326 AND symb_decoder(16#29#)) OR
 					(reg_q2326 AND symb_decoder(16#54#)) OR
 					(reg_q2326 AND symb_decoder(16#c7#)) OR
 					(reg_q2326 AND symb_decoder(16#7e#)) OR
 					(reg_q2326 AND symb_decoder(16#6a#)) OR
 					(reg_q2326 AND symb_decoder(16#c8#)) OR
 					(reg_q2326 AND symb_decoder(16#08#)) OR
 					(reg_q2326 AND symb_decoder(16#eb#)) OR
 					(reg_q2326 AND symb_decoder(16#ce#)) OR
 					(reg_q2326 AND symb_decoder(16#a9#)) OR
 					(reg_q2326 AND symb_decoder(16#10#)) OR
 					(reg_q2326 AND symb_decoder(16#22#)) OR
 					(reg_q2326 AND symb_decoder(16#02#)) OR
 					(reg_q2326 AND symb_decoder(16#a3#)) OR
 					(reg_q2326 AND symb_decoder(16#e3#)) OR
 					(reg_q2326 AND symb_decoder(16#4e#)) OR
 					(reg_q2326 AND symb_decoder(16#85#)) OR
 					(reg_q2326 AND symb_decoder(16#c4#)) OR
 					(reg_q2326 AND symb_decoder(16#6c#)) OR
 					(reg_q2326 AND symb_decoder(16#8e#)) OR
 					(reg_q2326 AND symb_decoder(16#9f#)) OR
 					(reg_q2326 AND symb_decoder(16#d4#)) OR
 					(reg_q2326 AND symb_decoder(16#75#)) OR
 					(reg_q2326 AND symb_decoder(16#6f#)) OR
 					(reg_q2326 AND symb_decoder(16#da#)) OR
 					(reg_q2326 AND symb_decoder(16#90#)) OR
 					(reg_q2326 AND symb_decoder(16#07#)) OR
 					(reg_q2326 AND symb_decoder(16#8f#)) OR
 					(reg_q2326 AND symb_decoder(16#12#)) OR
 					(reg_q2326 AND symb_decoder(16#a7#)) OR
 					(reg_q2326 AND symb_decoder(16#39#)) OR
 					(reg_q2326 AND symb_decoder(16#70#)) OR
 					(reg_q2326 AND symb_decoder(16#d2#)) OR
 					(reg_q2326 AND symb_decoder(16#a6#)) OR
 					(reg_q2326 AND symb_decoder(16#e4#)) OR
 					(reg_q2326 AND symb_decoder(16#f4#)) OR
 					(reg_q2326 AND symb_decoder(16#0e#)) OR
 					(reg_q2326 AND symb_decoder(16#e8#)) OR
 					(reg_q2326 AND symb_decoder(16#d1#)) OR
 					(reg_q2326 AND symb_decoder(16#78#)) OR
 					(reg_q2326 AND symb_decoder(16#c9#)) OR
 					(reg_q2326 AND symb_decoder(16#3f#)) OR
 					(reg_q2326 AND symb_decoder(16#13#)) OR
 					(reg_q2326 AND symb_decoder(16#26#)) OR
 					(reg_q2326 AND symb_decoder(16#64#)) OR
 					(reg_q2326 AND symb_decoder(16#87#)) OR
 					(reg_q2326 AND symb_decoder(16#99#)) OR
 					(reg_q2326 AND symb_decoder(16#aa#)) OR
 					(reg_q2326 AND symb_decoder(16#ee#)) OR
 					(reg_q2326 AND symb_decoder(16#48#)) OR
 					(reg_q2326 AND symb_decoder(16#25#)) OR
 					(reg_q2326 AND symb_decoder(16#19#)) OR
 					(reg_q2326 AND symb_decoder(16#cb#)) OR
 					(reg_q2326 AND symb_decoder(16#1b#)) OR
 					(reg_q2326 AND symb_decoder(16#ac#)) OR
 					(reg_q2326 AND symb_decoder(16#d6#)) OR
 					(reg_q2326 AND symb_decoder(16#fd#)) OR
 					(reg_q2326 AND symb_decoder(16#84#)) OR
 					(reg_q2326 AND symb_decoder(16#cc#)) OR
 					(reg_q2326 AND symb_decoder(16#59#)) OR
 					(reg_q2326 AND symb_decoder(16#32#)) OR
 					(reg_q2326 AND symb_decoder(16#79#)) OR
 					(reg_q2326 AND symb_decoder(16#3b#)) OR
 					(reg_q2326 AND symb_decoder(16#6d#)) OR
 					(reg_q2326 AND symb_decoder(16#c3#)) OR
 					(reg_q2326 AND symb_decoder(16#11#)) OR
 					(reg_q2326 AND symb_decoder(16#9b#)) OR
 					(reg_q2326 AND symb_decoder(16#e5#)) OR
 					(reg_q2326 AND symb_decoder(16#31#)) OR
 					(reg_q2326 AND symb_decoder(16#2e#)) OR
 					(reg_q2326 AND symb_decoder(16#8b#)) OR
 					(reg_q2326 AND symb_decoder(16#b5#)) OR
 					(reg_q2326 AND symb_decoder(16#d8#)) OR
 					(reg_q2326 AND symb_decoder(16#1a#)) OR
 					(reg_q2326 AND symb_decoder(16#ae#)) OR
 					(reg_q2326 AND symb_decoder(16#61#)) OR
 					(reg_q2326 AND symb_decoder(16#8d#)) OR
 					(reg_q2326 AND symb_decoder(16#2a#)) OR
 					(reg_q2326 AND symb_decoder(16#4c#)) OR
 					(reg_q2326 AND symb_decoder(16#0b#)) OR
 					(reg_q2326 AND symb_decoder(16#b2#)) OR
 					(reg_q2326 AND symb_decoder(16#ca#)) OR
 					(reg_q2326 AND symb_decoder(16#45#)) OR
 					(reg_q2326 AND symb_decoder(16#ad#)) OR
 					(reg_q2326 AND symb_decoder(16#38#)) OR
 					(reg_q2326 AND symb_decoder(16#20#)) OR
 					(reg_q2326 AND symb_decoder(16#f0#)) OR
 					(reg_q2326 AND symb_decoder(16#46#)) OR
 					(reg_q2326 AND symb_decoder(16#15#)) OR
 					(reg_q2326 AND symb_decoder(16#73#)) OR
 					(reg_q2326 AND symb_decoder(16#c1#)) OR
 					(reg_q2326 AND symb_decoder(16#4d#)) OR
 					(reg_q2326 AND symb_decoder(16#a5#)) OR
 					(reg_q2326 AND symb_decoder(16#3c#)) OR
 					(reg_q2326 AND symb_decoder(16#42#));
reg_q2584_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2583 AND symb_decoder(16#0a#)) OR
 					(reg_q2583 AND symb_decoder(16#0d#));
reg_fullgraph64_init <= "00";

reg_fullgraph64_sel <= "00" & reg_q2584_in & reg_q2326_in;

	--coder fullgraph64
with reg_fullgraph64_sel select
reg_fullgraph64_in <=
	"01" when "0001",
	"10" when "0010",
	"00" when others;
 --end coder

	p_reg_fullgraph64: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph64 <= reg_fullgraph64_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph64 <= reg_fullgraph64_init;
        else
          reg_fullgraph64 <= reg_fullgraph64_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph64

		reg_q2326 <= '1' when reg_fullgraph64 = "01" else '0'; 
		reg_q2584 <= '1' when reg_fullgraph64 = "10" else '0'; 
--end decoder 

reg_q1022_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1022 AND symb_decoder(16#42#)) OR
 					(reg_q1022 AND symb_decoder(16#3a#)) OR
 					(reg_q1022 AND symb_decoder(16#73#)) OR
 					(reg_q1022 AND symb_decoder(16#0e#)) OR
 					(reg_q1022 AND symb_decoder(16#8e#)) OR
 					(reg_q1022 AND symb_decoder(16#1b#)) OR
 					(reg_q1022 AND symb_decoder(16#51#)) OR
 					(reg_q1022 AND symb_decoder(16#65#)) OR
 					(reg_q1022 AND symb_decoder(16#a8#)) OR
 					(reg_q1022 AND symb_decoder(16#eb#)) OR
 					(reg_q1022 AND symb_decoder(16#32#)) OR
 					(reg_q1022 AND symb_decoder(16#53#)) OR
 					(reg_q1022 AND symb_decoder(16#87#)) OR
 					(reg_q1022 AND symb_decoder(16#de#)) OR
 					(reg_q1022 AND symb_decoder(16#e3#)) OR
 					(reg_q1022 AND symb_decoder(16#b7#)) OR
 					(reg_q1022 AND symb_decoder(16#03#)) OR
 					(reg_q1022 AND symb_decoder(16#59#)) OR
 					(reg_q1022 AND symb_decoder(16#ad#)) OR
 					(reg_q1022 AND symb_decoder(16#6c#)) OR
 					(reg_q1022 AND symb_decoder(16#58#)) OR
 					(reg_q1022 AND symb_decoder(16#d0#)) OR
 					(reg_q1022 AND symb_decoder(16#d1#)) OR
 					(reg_q1022 AND symb_decoder(16#21#)) OR
 					(reg_q1022 AND symb_decoder(16#d7#)) OR
 					(reg_q1022 AND symb_decoder(16#22#)) OR
 					(reg_q1022 AND symb_decoder(16#43#)) OR
 					(reg_q1022 AND symb_decoder(16#16#)) OR
 					(reg_q1022 AND symb_decoder(16#ba#)) OR
 					(reg_q1022 AND symb_decoder(16#40#)) OR
 					(reg_q1022 AND symb_decoder(16#f9#)) OR
 					(reg_q1022 AND symb_decoder(16#bb#)) OR
 					(reg_q1022 AND symb_decoder(16#bc#)) OR
 					(reg_q1022 AND symb_decoder(16#88#)) OR
 					(reg_q1022 AND symb_decoder(16#34#)) OR
 					(reg_q1022 AND symb_decoder(16#d3#)) OR
 					(reg_q1022 AND symb_decoder(16#6b#)) OR
 					(reg_q1022 AND symb_decoder(16#75#)) OR
 					(reg_q1022 AND symb_decoder(16#c6#)) OR
 					(reg_q1022 AND symb_decoder(16#79#)) OR
 					(reg_q1022 AND symb_decoder(16#0d#)) OR
 					(reg_q1022 AND symb_decoder(16#39#)) OR
 					(reg_q1022 AND symb_decoder(16#31#)) OR
 					(reg_q1022 AND symb_decoder(16#47#)) OR
 					(reg_q1022 AND symb_decoder(16#5b#)) OR
 					(reg_q1022 AND symb_decoder(16#b0#)) OR
 					(reg_q1022 AND symb_decoder(16#7e#)) OR
 					(reg_q1022 AND symb_decoder(16#a6#)) OR
 					(reg_q1022 AND symb_decoder(16#12#)) OR
 					(reg_q1022 AND symb_decoder(16#61#)) OR
 					(reg_q1022 AND symb_decoder(16#66#)) OR
 					(reg_q1022 AND symb_decoder(16#8a#)) OR
 					(reg_q1022 AND symb_decoder(16#4a#)) OR
 					(reg_q1022 AND symb_decoder(16#7a#)) OR
 					(reg_q1022 AND symb_decoder(16#f5#)) OR
 					(reg_q1022 AND symb_decoder(16#18#)) OR
 					(reg_q1022 AND symb_decoder(16#8c#)) OR
 					(reg_q1022 AND symb_decoder(16#d4#)) OR
 					(reg_q1022 AND symb_decoder(16#dd#)) OR
 					(reg_q1022 AND symb_decoder(16#67#)) OR
 					(reg_q1022 AND symb_decoder(16#3d#)) OR
 					(reg_q1022 AND symb_decoder(16#13#)) OR
 					(reg_q1022 AND symb_decoder(16#df#)) OR
 					(reg_q1022 AND symb_decoder(16#c5#)) OR
 					(reg_q1022 AND symb_decoder(16#ae#)) OR
 					(reg_q1022 AND symb_decoder(16#3c#)) OR
 					(reg_q1022 AND symb_decoder(16#af#)) OR
 					(reg_q1022 AND symb_decoder(16#24#)) OR
 					(reg_q1022 AND symb_decoder(16#dc#)) OR
 					(reg_q1022 AND symb_decoder(16#60#)) OR
 					(reg_q1022 AND symb_decoder(16#69#)) OR
 					(reg_q1022 AND symb_decoder(16#71#)) OR
 					(reg_q1022 AND symb_decoder(16#e4#)) OR
 					(reg_q1022 AND symb_decoder(16#e7#)) OR
 					(reg_q1022 AND symb_decoder(16#c8#)) OR
 					(reg_q1022 AND symb_decoder(16#ca#)) OR
 					(reg_q1022 AND symb_decoder(16#1c#)) OR
 					(reg_q1022 AND symb_decoder(16#48#)) OR
 					(reg_q1022 AND symb_decoder(16#17#)) OR
 					(reg_q1022 AND symb_decoder(16#08#)) OR
 					(reg_q1022 AND symb_decoder(16#fa#)) OR
 					(reg_q1022 AND symb_decoder(16#a7#)) OR
 					(reg_q1022 AND symb_decoder(16#4b#)) OR
 					(reg_q1022 AND symb_decoder(16#ed#)) OR
 					(reg_q1022 AND symb_decoder(16#11#)) OR
 					(reg_q1022 AND symb_decoder(16#74#)) OR
 					(reg_q1022 AND symb_decoder(16#c0#)) OR
 					(reg_q1022 AND symb_decoder(16#b5#)) OR
 					(reg_q1022 AND symb_decoder(16#a1#)) OR
 					(reg_q1022 AND symb_decoder(16#14#)) OR
 					(reg_q1022 AND symb_decoder(16#30#)) OR
 					(reg_q1022 AND symb_decoder(16#e2#)) OR
 					(reg_q1022 AND symb_decoder(16#f0#)) OR
 					(reg_q1022 AND symb_decoder(16#84#)) OR
 					(reg_q1022 AND symb_decoder(16#9f#)) OR
 					(reg_q1022 AND symb_decoder(16#ec#)) OR
 					(reg_q1022 AND symb_decoder(16#27#)) OR
 					(reg_q1022 AND symb_decoder(16#cd#)) OR
 					(reg_q1022 AND symb_decoder(16#9d#)) OR
 					(reg_q1022 AND symb_decoder(16#b8#)) OR
 					(reg_q1022 AND symb_decoder(16#82#)) OR
 					(reg_q1022 AND symb_decoder(16#c9#)) OR
 					(reg_q1022 AND symb_decoder(16#89#)) OR
 					(reg_q1022 AND symb_decoder(16#2c#)) OR
 					(reg_q1022 AND symb_decoder(16#6f#)) OR
 					(reg_q1022 AND symb_decoder(16#68#)) OR
 					(reg_q1022 AND symb_decoder(16#9b#)) OR
 					(reg_q1022 AND symb_decoder(16#50#)) OR
 					(reg_q1022 AND symb_decoder(16#98#)) OR
 					(reg_q1022 AND symb_decoder(16#c2#)) OR
 					(reg_q1022 AND symb_decoder(16#19#)) OR
 					(reg_q1022 AND symb_decoder(16#2f#)) OR
 					(reg_q1022 AND symb_decoder(16#0b#)) OR
 					(reg_q1022 AND symb_decoder(16#fe#)) OR
 					(reg_q1022 AND symb_decoder(16#46#)) OR
 					(reg_q1022 AND symb_decoder(16#95#)) OR
 					(reg_q1022 AND symb_decoder(16#ce#)) OR
 					(reg_q1022 AND symb_decoder(16#91#)) OR
 					(reg_q1022 AND symb_decoder(16#49#)) OR
 					(reg_q1022 AND symb_decoder(16#9e#)) OR
 					(reg_q1022 AND symb_decoder(16#15#)) OR
 					(reg_q1022 AND symb_decoder(16#ee#)) OR
 					(reg_q1022 AND symb_decoder(16#54#)) OR
 					(reg_q1022 AND symb_decoder(16#bd#)) OR
 					(reg_q1022 AND symb_decoder(16#0f#)) OR
 					(reg_q1022 AND symb_decoder(16#99#)) OR
 					(reg_q1022 AND symb_decoder(16#76#)) OR
 					(reg_q1022 AND symb_decoder(16#6d#)) OR
 					(reg_q1022 AND symb_decoder(16#f3#)) OR
 					(reg_q1022 AND symb_decoder(16#a0#)) OR
 					(reg_q1022 AND symb_decoder(16#4e#)) OR
 					(reg_q1022 AND symb_decoder(16#b3#)) OR
 					(reg_q1022 AND symb_decoder(16#10#)) OR
 					(reg_q1022 AND symb_decoder(16#9c#)) OR
 					(reg_q1022 AND symb_decoder(16#77#)) OR
 					(reg_q1022 AND symb_decoder(16#04#)) OR
 					(reg_q1022 AND symb_decoder(16#0c#)) OR
 					(reg_q1022 AND symb_decoder(16#f2#)) OR
 					(reg_q1022 AND symb_decoder(16#5a#)) OR
 					(reg_q1022 AND symb_decoder(16#55#)) OR
 					(reg_q1022 AND symb_decoder(16#5f#)) OR
 					(reg_q1022 AND symb_decoder(16#38#)) OR
 					(reg_q1022 AND symb_decoder(16#1e#)) OR
 					(reg_q1022 AND symb_decoder(16#96#)) OR
 					(reg_q1022 AND symb_decoder(16#e8#)) OR
 					(reg_q1022 AND symb_decoder(16#c1#)) OR
 					(reg_q1022 AND symb_decoder(16#a2#)) OR
 					(reg_q1022 AND symb_decoder(16#b2#)) OR
 					(reg_q1022 AND symb_decoder(16#3e#)) OR
 					(reg_q1022 AND symb_decoder(16#fb#)) OR
 					(reg_q1022 AND symb_decoder(16#b4#)) OR
 					(reg_q1022 AND symb_decoder(16#37#)) OR
 					(reg_q1022 AND symb_decoder(16#2e#)) OR
 					(reg_q1022 AND symb_decoder(16#6a#)) OR
 					(reg_q1022 AND symb_decoder(16#e5#)) OR
 					(reg_q1022 AND symb_decoder(16#e9#)) OR
 					(reg_q1022 AND symb_decoder(16#1a#)) OR
 					(reg_q1022 AND symb_decoder(16#fd#)) OR
 					(reg_q1022 AND symb_decoder(16#33#)) OR
 					(reg_q1022 AND symb_decoder(16#01#)) OR
 					(reg_q1022 AND symb_decoder(16#ab#)) OR
 					(reg_q1022 AND symb_decoder(16#b1#)) OR
 					(reg_q1022 AND symb_decoder(16#f6#)) OR
 					(reg_q1022 AND symb_decoder(16#70#)) OR
 					(reg_q1022 AND symb_decoder(16#c7#)) OR
 					(reg_q1022 AND symb_decoder(16#2b#)) OR
 					(reg_q1022 AND symb_decoder(16#a3#)) OR
 					(reg_q1022 AND symb_decoder(16#56#)) OR
 					(reg_q1022 AND symb_decoder(16#90#)) OR
 					(reg_q1022 AND symb_decoder(16#d6#)) OR
 					(reg_q1022 AND symb_decoder(16#be#)) OR
 					(reg_q1022 AND symb_decoder(16#5c#)) OR
 					(reg_q1022 AND symb_decoder(16#5d#)) OR
 					(reg_q1022 AND symb_decoder(16#b6#)) OR
 					(reg_q1022 AND symb_decoder(16#e6#)) OR
 					(reg_q1022 AND symb_decoder(16#f4#)) OR
 					(reg_q1022 AND symb_decoder(16#bf#)) OR
 					(reg_q1022 AND symb_decoder(16#4f#)) OR
 					(reg_q1022 AND symb_decoder(16#fc#)) OR
 					(reg_q1022 AND symb_decoder(16#c4#)) OR
 					(reg_q1022 AND symb_decoder(16#b9#)) OR
 					(reg_q1022 AND symb_decoder(16#ef#)) OR
 					(reg_q1022 AND symb_decoder(16#93#)) OR
 					(reg_q1022 AND symb_decoder(16#85#)) OR
 					(reg_q1022 AND symb_decoder(16#80#)) OR
 					(reg_q1022 AND symb_decoder(16#02#)) OR
 					(reg_q1022 AND symb_decoder(16#a5#)) OR
 					(reg_q1022 AND symb_decoder(16#1f#)) OR
 					(reg_q1022 AND symb_decoder(16#da#)) OR
 					(reg_q1022 AND symb_decoder(16#07#)) OR
 					(reg_q1022 AND symb_decoder(16#2a#)) OR
 					(reg_q1022 AND symb_decoder(16#d9#)) OR
 					(reg_q1022 AND symb_decoder(16#4c#)) OR
 					(reg_q1022 AND symb_decoder(16#d5#)) OR
 					(reg_q1022 AND symb_decoder(16#7f#)) OR
 					(reg_q1022 AND symb_decoder(16#a9#)) OR
 					(reg_q1022 AND symb_decoder(16#35#)) OR
 					(reg_q1022 AND symb_decoder(16#97#)) OR
 					(reg_q1022 AND symb_decoder(16#86#)) OR
 					(reg_q1022 AND symb_decoder(16#aa#)) OR
 					(reg_q1022 AND symb_decoder(16#00#)) OR
 					(reg_q1022 AND symb_decoder(16#29#)) OR
 					(reg_q1022 AND symb_decoder(16#52#)) OR
 					(reg_q1022 AND symb_decoder(16#36#)) OR
 					(reg_q1022 AND symb_decoder(16#d8#)) OR
 					(reg_q1022 AND symb_decoder(16#7c#)) OR
 					(reg_q1022 AND symb_decoder(16#81#)) OR
 					(reg_q1022 AND symb_decoder(16#63#)) OR
 					(reg_q1022 AND symb_decoder(16#5e#)) OR
 					(reg_q1022 AND symb_decoder(16#d2#)) OR
 					(reg_q1022 AND symb_decoder(16#94#)) OR
 					(reg_q1022 AND symb_decoder(16#28#)) OR
 					(reg_q1022 AND symb_decoder(16#0a#)) OR
 					(reg_q1022 AND symb_decoder(16#83#)) OR
 					(reg_q1022 AND symb_decoder(16#7d#)) OR
 					(reg_q1022 AND symb_decoder(16#cb#)) OR
 					(reg_q1022 AND symb_decoder(16#06#)) OR
 					(reg_q1022 AND symb_decoder(16#8b#)) OR
 					(reg_q1022 AND symb_decoder(16#e0#)) OR
 					(reg_q1022 AND symb_decoder(16#8f#)) OR
 					(reg_q1022 AND symb_decoder(16#25#)) OR
 					(reg_q1022 AND symb_decoder(16#4d#)) OR
 					(reg_q1022 AND symb_decoder(16#20#)) OR
 					(reg_q1022 AND symb_decoder(16#9a#)) OR
 					(reg_q1022 AND symb_decoder(16#c3#)) OR
 					(reg_q1022 AND symb_decoder(16#23#)) OR
 					(reg_q1022 AND symb_decoder(16#db#)) OR
 					(reg_q1022 AND symb_decoder(16#3f#)) OR
 					(reg_q1022 AND symb_decoder(16#f8#)) OR
 					(reg_q1022 AND symb_decoder(16#26#)) OR
 					(reg_q1022 AND symb_decoder(16#72#)) OR
 					(reg_q1022 AND symb_decoder(16#ac#)) OR
 					(reg_q1022 AND symb_decoder(16#05#)) OR
 					(reg_q1022 AND symb_decoder(16#f1#)) OR
 					(reg_q1022 AND symb_decoder(16#8d#)) OR
 					(reg_q1022 AND symb_decoder(16#2d#)) OR
 					(reg_q1022 AND symb_decoder(16#ff#)) OR
 					(reg_q1022 AND symb_decoder(16#44#)) OR
 					(reg_q1022 AND symb_decoder(16#e1#)) OR
 					(reg_q1022 AND symb_decoder(16#cc#)) OR
 					(reg_q1022 AND symb_decoder(16#62#)) OR
 					(reg_q1022 AND symb_decoder(16#cf#)) OR
 					(reg_q1022 AND symb_decoder(16#45#)) OR
 					(reg_q1022 AND symb_decoder(16#64#)) OR
 					(reg_q1022 AND symb_decoder(16#09#)) OR
 					(reg_q1022 AND symb_decoder(16#57#)) OR
 					(reg_q1022 AND symb_decoder(16#3b#)) OR
 					(reg_q1022 AND symb_decoder(16#41#)) OR
 					(reg_q1022 AND symb_decoder(16#f7#)) OR
 					(reg_q1022 AND symb_decoder(16#ea#)) OR
 					(reg_q1022 AND symb_decoder(16#92#)) OR
 					(reg_q1022 AND symb_decoder(16#1d#)) OR
 					(reg_q1022 AND symb_decoder(16#78#)) OR
 					(reg_q1022 AND symb_decoder(16#a4#)) OR
 					(reg_q1022 AND symb_decoder(16#6e#)) OR
 					(reg_q1022 AND symb_decoder(16#7b#));
reg_q1022_init <= '0' ;
	p_reg_q1022: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1022 <= reg_q1022_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1022 <= reg_q1022_init;
        else
          reg_q1022 <= reg_q1022_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2221_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q2221 AND symb_decoder(16#47#)) OR
 					(reg_q2221 AND symb_decoder(16#37#)) OR
 					(reg_q2221 AND symb_decoder(16#48#)) OR
 					(reg_q2221 AND symb_decoder(16#df#)) OR
 					(reg_q2221 AND symb_decoder(16#3f#)) OR
 					(reg_q2221 AND symb_decoder(16#62#)) OR
 					(reg_q2221 AND symb_decoder(16#ee#)) OR
 					(reg_q2221 AND symb_decoder(16#68#)) OR
 					(reg_q2221 AND symb_decoder(16#ef#)) OR
 					(reg_q2221 AND symb_decoder(16#5e#)) OR
 					(reg_q2221 AND symb_decoder(16#52#)) OR
 					(reg_q2221 AND symb_decoder(16#d3#)) OR
 					(reg_q2221 AND symb_decoder(16#65#)) OR
 					(reg_q2221 AND symb_decoder(16#28#)) OR
 					(reg_q2221 AND symb_decoder(16#b7#)) OR
 					(reg_q2221 AND symb_decoder(16#cc#)) OR
 					(reg_q2221 AND symb_decoder(16#da#)) OR
 					(reg_q2221 AND symb_decoder(16#cb#)) OR
 					(reg_q2221 AND symb_decoder(16#f3#)) OR
 					(reg_q2221 AND symb_decoder(16#8b#)) OR
 					(reg_q2221 AND symb_decoder(16#81#)) OR
 					(reg_q2221 AND symb_decoder(16#04#)) OR
 					(reg_q2221 AND symb_decoder(16#fc#)) OR
 					(reg_q2221 AND symb_decoder(16#fb#)) OR
 					(reg_q2221 AND symb_decoder(16#c6#)) OR
 					(reg_q2221 AND symb_decoder(16#8c#)) OR
 					(reg_q2221 AND symb_decoder(16#59#)) OR
 					(reg_q2221 AND symb_decoder(16#b4#)) OR
 					(reg_q2221 AND symb_decoder(16#d7#)) OR
 					(reg_q2221 AND symb_decoder(16#75#)) OR
 					(reg_q2221 AND symb_decoder(16#02#)) OR
 					(reg_q2221 AND symb_decoder(16#8a#)) OR
 					(reg_q2221 AND symb_decoder(16#bd#)) OR
 					(reg_q2221 AND symb_decoder(16#18#)) OR
 					(reg_q2221 AND symb_decoder(16#1e#)) OR
 					(reg_q2221 AND symb_decoder(16#79#)) OR
 					(reg_q2221 AND symb_decoder(16#a3#)) OR
 					(reg_q2221 AND symb_decoder(16#49#)) OR
 					(reg_q2221 AND symb_decoder(16#57#)) OR
 					(reg_q2221 AND symb_decoder(16#1d#)) OR
 					(reg_q2221 AND symb_decoder(16#b1#)) OR
 					(reg_q2221 AND symb_decoder(16#85#)) OR
 					(reg_q2221 AND symb_decoder(16#1a#)) OR
 					(reg_q2221 AND symb_decoder(16#b6#)) OR
 					(reg_q2221 AND symb_decoder(16#96#)) OR
 					(reg_q2221 AND symb_decoder(16#4f#)) OR
 					(reg_q2221 AND symb_decoder(16#a6#)) OR
 					(reg_q2221 AND symb_decoder(16#89#)) OR
 					(reg_q2221 AND symb_decoder(16#03#)) OR
 					(reg_q2221 AND symb_decoder(16#3b#)) OR
 					(reg_q2221 AND symb_decoder(16#ab#)) OR
 					(reg_q2221 AND symb_decoder(16#ac#)) OR
 					(reg_q2221 AND symb_decoder(16#6c#)) OR
 					(reg_q2221 AND symb_decoder(16#0f#)) OR
 					(reg_q2221 AND symb_decoder(16#b0#)) OR
 					(reg_q2221 AND symb_decoder(16#11#)) OR
 					(reg_q2221 AND symb_decoder(16#3e#)) OR
 					(reg_q2221 AND symb_decoder(16#e8#)) OR
 					(reg_q2221 AND symb_decoder(16#a9#)) OR
 					(reg_q2221 AND symb_decoder(16#4e#)) OR
 					(reg_q2221 AND symb_decoder(16#cd#)) OR
 					(reg_q2221 AND symb_decoder(16#15#)) OR
 					(reg_q2221 AND symb_decoder(16#ba#)) OR
 					(reg_q2221 AND symb_decoder(16#db#)) OR
 					(reg_q2221 AND symb_decoder(16#22#)) OR
 					(reg_q2221 AND symb_decoder(16#5d#)) OR
 					(reg_q2221 AND symb_decoder(16#de#)) OR
 					(reg_q2221 AND symb_decoder(16#93#)) OR
 					(reg_q2221 AND symb_decoder(16#6e#)) OR
 					(reg_q2221 AND symb_decoder(16#00#)) OR
 					(reg_q2221 AND symb_decoder(16#14#)) OR
 					(reg_q2221 AND symb_decoder(16#c9#)) OR
 					(reg_q2221 AND symb_decoder(16#9c#)) OR
 					(reg_q2221 AND symb_decoder(16#b8#)) OR
 					(reg_q2221 AND symb_decoder(16#9f#)) OR
 					(reg_q2221 AND symb_decoder(16#4c#)) OR
 					(reg_q2221 AND symb_decoder(16#50#)) OR
 					(reg_q2221 AND symb_decoder(16#b5#)) OR
 					(reg_q2221 AND symb_decoder(16#bc#)) OR
 					(reg_q2221 AND symb_decoder(16#fa#)) OR
 					(reg_q2221 AND symb_decoder(16#9d#)) OR
 					(reg_q2221 AND symb_decoder(16#e6#)) OR
 					(reg_q2221 AND symb_decoder(16#71#)) OR
 					(reg_q2221 AND symb_decoder(16#0d#)) OR
 					(reg_q2221 AND symb_decoder(16#6f#)) OR
 					(reg_q2221 AND symb_decoder(16#56#)) OR
 					(reg_q2221 AND symb_decoder(16#f9#)) OR
 					(reg_q2221 AND symb_decoder(16#f1#)) OR
 					(reg_q2221 AND symb_decoder(16#0a#)) OR
 					(reg_q2221 AND symb_decoder(16#1c#)) OR
 					(reg_q2221 AND symb_decoder(16#44#)) OR
 					(reg_q2221 AND symb_decoder(16#b9#)) OR
 					(reg_q2221 AND symb_decoder(16#dd#)) OR
 					(reg_q2221 AND symb_decoder(16#8f#)) OR
 					(reg_q2221 AND symb_decoder(16#33#)) OR
 					(reg_q2221 AND symb_decoder(16#3d#)) OR
 					(reg_q2221 AND symb_decoder(16#e2#)) OR
 					(reg_q2221 AND symb_decoder(16#8e#)) OR
 					(reg_q2221 AND symb_decoder(16#8d#)) OR
 					(reg_q2221 AND symb_decoder(16#5f#)) OR
 					(reg_q2221 AND symb_decoder(16#26#)) OR
 					(reg_q2221 AND symb_decoder(16#a2#)) OR
 					(reg_q2221 AND symb_decoder(16#86#)) OR
 					(reg_q2221 AND symb_decoder(16#5c#)) OR
 					(reg_q2221 AND symb_decoder(16#38#)) OR
 					(reg_q2221 AND symb_decoder(16#f7#)) OR
 					(reg_q2221 AND symb_decoder(16#b2#)) OR
 					(reg_q2221 AND symb_decoder(16#6b#)) OR
 					(reg_q2221 AND symb_decoder(16#36#)) OR
 					(reg_q2221 AND symb_decoder(16#13#)) OR
 					(reg_q2221 AND symb_decoder(16#b3#)) OR
 					(reg_q2221 AND symb_decoder(16#16#)) OR
 					(reg_q2221 AND symb_decoder(16#39#)) OR
 					(reg_q2221 AND symb_decoder(16#94#)) OR
 					(reg_q2221 AND symb_decoder(16#07#)) OR
 					(reg_q2221 AND symb_decoder(16#a8#)) OR
 					(reg_q2221 AND symb_decoder(16#63#)) OR
 					(reg_q2221 AND symb_decoder(16#20#)) OR
 					(reg_q2221 AND symb_decoder(16#d8#)) OR
 					(reg_q2221 AND symb_decoder(16#05#)) OR
 					(reg_q2221 AND symb_decoder(16#ff#)) OR
 					(reg_q2221 AND symb_decoder(16#53#)) OR
 					(reg_q2221 AND symb_decoder(16#4d#)) OR
 					(reg_q2221 AND symb_decoder(16#3a#)) OR
 					(reg_q2221 AND symb_decoder(16#fd#)) OR
 					(reg_q2221 AND symb_decoder(16#98#)) OR
 					(reg_q2221 AND symb_decoder(16#97#)) OR
 					(reg_q2221 AND symb_decoder(16#d9#)) OR
 					(reg_q2221 AND symb_decoder(16#6d#)) OR
 					(reg_q2221 AND symb_decoder(16#51#)) OR
 					(reg_q2221 AND symb_decoder(16#5a#)) OR
 					(reg_q2221 AND symb_decoder(16#3c#)) OR
 					(reg_q2221 AND symb_decoder(16#41#)) OR
 					(reg_q2221 AND symb_decoder(16#f6#)) OR
 					(reg_q2221 AND symb_decoder(16#25#)) OR
 					(reg_q2221 AND symb_decoder(16#e7#)) OR
 					(reg_q2221 AND symb_decoder(16#aa#)) OR
 					(reg_q2221 AND symb_decoder(16#23#)) OR
 					(reg_q2221 AND symb_decoder(16#01#)) OR
 					(reg_q2221 AND symb_decoder(16#0b#)) OR
 					(reg_q2221 AND symb_decoder(16#ad#)) OR
 					(reg_q2221 AND symb_decoder(16#ca#)) OR
 					(reg_q2221 AND symb_decoder(16#7d#)) OR
 					(reg_q2221 AND symb_decoder(16#46#)) OR
 					(reg_q2221 AND symb_decoder(16#c5#)) OR
 					(reg_q2221 AND symb_decoder(16#c7#)) OR
 					(reg_q2221 AND symb_decoder(16#1b#)) OR
 					(reg_q2221 AND symb_decoder(16#fe#)) OR
 					(reg_q2221 AND symb_decoder(16#a1#)) OR
 					(reg_q2221 AND symb_decoder(16#08#)) OR
 					(reg_q2221 AND symb_decoder(16#c1#)) OR
 					(reg_q2221 AND symb_decoder(16#7b#)) OR
 					(reg_q2221 AND symb_decoder(16#7e#)) OR
 					(reg_q2221 AND symb_decoder(16#2c#)) OR
 					(reg_q2221 AND symb_decoder(16#e0#)) OR
 					(reg_q2221 AND symb_decoder(16#60#)) OR
 					(reg_q2221 AND symb_decoder(16#12#)) OR
 					(reg_q2221 AND symb_decoder(16#a5#)) OR
 					(reg_q2221 AND symb_decoder(16#7c#)) OR
 					(reg_q2221 AND symb_decoder(16#0c#)) OR
 					(reg_q2221 AND symb_decoder(16#24#)) OR
 					(reg_q2221 AND symb_decoder(16#90#)) OR
 					(reg_q2221 AND symb_decoder(16#dc#)) OR
 					(reg_q2221 AND symb_decoder(16#27#)) OR
 					(reg_q2221 AND symb_decoder(16#35#)) OR
 					(reg_q2221 AND symb_decoder(16#9b#)) OR
 					(reg_q2221 AND symb_decoder(16#99#)) OR
 					(reg_q2221 AND symb_decoder(16#ae#)) OR
 					(reg_q2221 AND symb_decoder(16#f0#)) OR
 					(reg_q2221 AND symb_decoder(16#d6#)) OR
 					(reg_q2221 AND symb_decoder(16#66#)) OR
 					(reg_q2221 AND symb_decoder(16#f5#)) OR
 					(reg_q2221 AND symb_decoder(16#17#)) OR
 					(reg_q2221 AND symb_decoder(16#eb#)) OR
 					(reg_q2221 AND symb_decoder(16#a7#)) OR
 					(reg_q2221 AND symb_decoder(16#30#)) OR
 					(reg_q2221 AND symb_decoder(16#80#)) OR
 					(reg_q2221 AND symb_decoder(16#a0#)) OR
 					(reg_q2221 AND symb_decoder(16#ed#)) OR
 					(reg_q2221 AND symb_decoder(16#cf#)) OR
 					(reg_q2221 AND symb_decoder(16#92#)) OR
 					(reg_q2221 AND symb_decoder(16#4b#)) OR
 					(reg_q2221 AND symb_decoder(16#c8#)) OR
 					(reg_q2221 AND symb_decoder(16#42#)) OR
 					(reg_q2221 AND symb_decoder(16#72#)) OR
 					(reg_q2221 AND symb_decoder(16#54#)) OR
 					(reg_q2221 AND symb_decoder(16#87#)) OR
 					(reg_q2221 AND symb_decoder(16#45#)) OR
 					(reg_q2221 AND symb_decoder(16#73#)) OR
 					(reg_q2221 AND symb_decoder(16#43#)) OR
 					(reg_q2221 AND symb_decoder(16#10#)) OR
 					(reg_q2221 AND symb_decoder(16#21#)) OR
 					(reg_q2221 AND symb_decoder(16#83#)) OR
 					(reg_q2221 AND symb_decoder(16#76#)) OR
 					(reg_q2221 AND symb_decoder(16#29#)) OR
 					(reg_q2221 AND symb_decoder(16#ce#)) OR
 					(reg_q2221 AND symb_decoder(16#4a#)) OR
 					(reg_q2221 AND symb_decoder(16#e4#)) OR
 					(reg_q2221 AND symb_decoder(16#31#)) OR
 					(reg_q2221 AND symb_decoder(16#06#)) OR
 					(reg_q2221 AND symb_decoder(16#82#)) OR
 					(reg_q2221 AND symb_decoder(16#2e#)) OR
 					(reg_q2221 AND symb_decoder(16#91#)) OR
 					(reg_q2221 AND symb_decoder(16#61#)) OR
 					(reg_q2221 AND symb_decoder(16#a4#)) OR
 					(reg_q2221 AND symb_decoder(16#5b#)) OR
 					(reg_q2221 AND symb_decoder(16#c0#)) OR
 					(reg_q2221 AND symb_decoder(16#e3#)) OR
 					(reg_q2221 AND symb_decoder(16#c2#)) OR
 					(reg_q2221 AND symb_decoder(16#e1#)) OR
 					(reg_q2221 AND symb_decoder(16#d1#)) OR
 					(reg_q2221 AND symb_decoder(16#e9#)) OR
 					(reg_q2221 AND symb_decoder(16#55#)) OR
 					(reg_q2221 AND symb_decoder(16#af#)) OR
 					(reg_q2221 AND symb_decoder(16#67#)) OR
 					(reg_q2221 AND symb_decoder(16#ec#)) OR
 					(reg_q2221 AND symb_decoder(16#69#)) OR
 					(reg_q2221 AND symb_decoder(16#d2#)) OR
 					(reg_q2221 AND symb_decoder(16#09#)) OR
 					(reg_q2221 AND symb_decoder(16#78#)) OR
 					(reg_q2221 AND symb_decoder(16#c3#)) OR
 					(reg_q2221 AND symb_decoder(16#7f#)) OR
 					(reg_q2221 AND symb_decoder(16#be#)) OR
 					(reg_q2221 AND symb_decoder(16#6a#)) OR
 					(reg_q2221 AND symb_decoder(16#c4#)) OR
 					(reg_q2221 AND symb_decoder(16#95#)) OR
 					(reg_q2221 AND symb_decoder(16#f2#)) OR
 					(reg_q2221 AND symb_decoder(16#32#)) OR
 					(reg_q2221 AND symb_decoder(16#bf#)) OR
 					(reg_q2221 AND symb_decoder(16#84#)) OR
 					(reg_q2221 AND symb_decoder(16#2d#)) OR
 					(reg_q2221 AND symb_decoder(16#9e#)) OR
 					(reg_q2221 AND symb_decoder(16#64#)) OR
 					(reg_q2221 AND symb_decoder(16#1f#)) OR
 					(reg_q2221 AND symb_decoder(16#f8#)) OR
 					(reg_q2221 AND symb_decoder(16#9a#)) OR
 					(reg_q2221 AND symb_decoder(16#2b#)) OR
 					(reg_q2221 AND symb_decoder(16#74#)) OR
 					(reg_q2221 AND symb_decoder(16#58#)) OR
 					(reg_q2221 AND symb_decoder(16#70#)) OR
 					(reg_q2221 AND symb_decoder(16#88#)) OR
 					(reg_q2221 AND symb_decoder(16#2f#)) OR
 					(reg_q2221 AND symb_decoder(16#7a#)) OR
 					(reg_q2221 AND symb_decoder(16#77#)) OR
 					(reg_q2221 AND symb_decoder(16#e5#)) OR
 					(reg_q2221 AND symb_decoder(16#34#)) OR
 					(reg_q2221 AND symb_decoder(16#d5#)) OR
 					(reg_q2221 AND symb_decoder(16#2a#)) OR
 					(reg_q2221 AND symb_decoder(16#bb#)) OR
 					(reg_q2221 AND symb_decoder(16#0e#)) OR
 					(reg_q2221 AND symb_decoder(16#40#)) OR
 					(reg_q2221 AND symb_decoder(16#d4#)) OR
 					(reg_q2221 AND symb_decoder(16#19#)) OR
 					(reg_q2221 AND symb_decoder(16#d0#)) OR
 					(reg_q2221 AND symb_decoder(16#f4#)) OR
 					(reg_q2221 AND symb_decoder(16#ea#));
reg_q2221_init <= '0' ;
	p_reg_q2221: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2221 <= reg_q2221_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2221 <= reg_q2221_init;
        else
          reg_q2221 <= reg_q2221_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q188_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q188 AND symb_decoder(16#e0#)) OR
 					(reg_q188 AND symb_decoder(16#63#)) OR
 					(reg_q188 AND symb_decoder(16#e8#)) OR
 					(reg_q188 AND symb_decoder(16#f4#)) OR
 					(reg_q188 AND symb_decoder(16#55#)) OR
 					(reg_q188 AND symb_decoder(16#ab#)) OR
 					(reg_q188 AND symb_decoder(16#10#)) OR
 					(reg_q188 AND symb_decoder(16#e7#)) OR
 					(reg_q188 AND symb_decoder(16#9f#)) OR
 					(reg_q188 AND symb_decoder(16#e2#)) OR
 					(reg_q188 AND symb_decoder(16#8a#)) OR
 					(reg_q188 AND symb_decoder(16#ef#)) OR
 					(reg_q188 AND symb_decoder(16#ce#)) OR
 					(reg_q188 AND symb_decoder(16#d6#)) OR
 					(reg_q188 AND symb_decoder(16#b2#)) OR
 					(reg_q188 AND symb_decoder(16#56#)) OR
 					(reg_q188 AND symb_decoder(16#2b#)) OR
 					(reg_q188 AND symb_decoder(16#58#)) OR
 					(reg_q188 AND symb_decoder(16#15#)) OR
 					(reg_q188 AND symb_decoder(16#43#)) OR
 					(reg_q188 AND symb_decoder(16#37#)) OR
 					(reg_q188 AND symb_decoder(16#54#)) OR
 					(reg_q188 AND symb_decoder(16#b0#)) OR
 					(reg_q188 AND symb_decoder(16#02#)) OR
 					(reg_q188 AND symb_decoder(16#39#)) OR
 					(reg_q188 AND symb_decoder(16#0c#)) OR
 					(reg_q188 AND symb_decoder(16#f1#)) OR
 					(reg_q188 AND symb_decoder(16#4e#)) OR
 					(reg_q188 AND symb_decoder(16#77#)) OR
 					(reg_q188 AND symb_decoder(16#81#)) OR
 					(reg_q188 AND symb_decoder(16#0a#)) OR
 					(reg_q188 AND symb_decoder(16#44#)) OR
 					(reg_q188 AND symb_decoder(16#a1#)) OR
 					(reg_q188 AND symb_decoder(16#07#)) OR
 					(reg_q188 AND symb_decoder(16#41#)) OR
 					(reg_q188 AND symb_decoder(16#b5#)) OR
 					(reg_q188 AND symb_decoder(16#23#)) OR
 					(reg_q188 AND symb_decoder(16#5b#)) OR
 					(reg_q188 AND symb_decoder(16#ec#)) OR
 					(reg_q188 AND symb_decoder(16#30#)) OR
 					(reg_q188 AND symb_decoder(16#b7#)) OR
 					(reg_q188 AND symb_decoder(16#76#)) OR
 					(reg_q188 AND symb_decoder(16#65#)) OR
 					(reg_q188 AND symb_decoder(16#59#)) OR
 					(reg_q188 AND symb_decoder(16#9a#)) OR
 					(reg_q188 AND symb_decoder(16#e4#)) OR
 					(reg_q188 AND symb_decoder(16#3b#)) OR
 					(reg_q188 AND symb_decoder(16#ae#)) OR
 					(reg_q188 AND symb_decoder(16#d0#)) OR
 					(reg_q188 AND symb_decoder(16#ee#)) OR
 					(reg_q188 AND symb_decoder(16#6d#)) OR
 					(reg_q188 AND symb_decoder(16#66#)) OR
 					(reg_q188 AND symb_decoder(16#c2#)) OR
 					(reg_q188 AND symb_decoder(16#b3#)) OR
 					(reg_q188 AND symb_decoder(16#33#)) OR
 					(reg_q188 AND symb_decoder(16#97#)) OR
 					(reg_q188 AND symb_decoder(16#0d#)) OR
 					(reg_q188 AND symb_decoder(16#4f#)) OR
 					(reg_q188 AND symb_decoder(16#cd#)) OR
 					(reg_q188 AND symb_decoder(16#eb#)) OR
 					(reg_q188 AND symb_decoder(16#1e#)) OR
 					(reg_q188 AND symb_decoder(16#27#)) OR
 					(reg_q188 AND symb_decoder(16#8e#)) OR
 					(reg_q188 AND symb_decoder(16#dd#)) OR
 					(reg_q188 AND symb_decoder(16#5e#)) OR
 					(reg_q188 AND symb_decoder(16#96#)) OR
 					(reg_q188 AND symb_decoder(16#6b#)) OR
 					(reg_q188 AND symb_decoder(16#a6#)) OR
 					(reg_q188 AND symb_decoder(16#af#)) OR
 					(reg_q188 AND symb_decoder(16#f6#)) OR
 					(reg_q188 AND symb_decoder(16#7e#)) OR
 					(reg_q188 AND symb_decoder(16#d1#)) OR
 					(reg_q188 AND symb_decoder(16#fb#)) OR
 					(reg_q188 AND symb_decoder(16#f0#)) OR
 					(reg_q188 AND symb_decoder(16#d3#)) OR
 					(reg_q188 AND symb_decoder(16#14#)) OR
 					(reg_q188 AND symb_decoder(16#6a#)) OR
 					(reg_q188 AND symb_decoder(16#4d#)) OR
 					(reg_q188 AND symb_decoder(16#62#)) OR
 					(reg_q188 AND symb_decoder(16#be#)) OR
 					(reg_q188 AND symb_decoder(16#b1#)) OR
 					(reg_q188 AND symb_decoder(16#a3#)) OR
 					(reg_q188 AND symb_decoder(16#c3#)) OR
 					(reg_q188 AND symb_decoder(16#78#)) OR
 					(reg_q188 AND symb_decoder(16#2e#)) OR
 					(reg_q188 AND symb_decoder(16#b8#)) OR
 					(reg_q188 AND symb_decoder(16#46#)) OR
 					(reg_q188 AND symb_decoder(16#e9#)) OR
 					(reg_q188 AND symb_decoder(16#2a#)) OR
 					(reg_q188 AND symb_decoder(16#83#)) OR
 					(reg_q188 AND symb_decoder(16#da#)) OR
 					(reg_q188 AND symb_decoder(16#0b#)) OR
 					(reg_q188 AND symb_decoder(16#7b#)) OR
 					(reg_q188 AND symb_decoder(16#38#)) OR
 					(reg_q188 AND symb_decoder(16#7d#)) OR
 					(reg_q188 AND symb_decoder(16#2c#)) OR
 					(reg_q188 AND symb_decoder(16#c4#)) OR
 					(reg_q188 AND symb_decoder(16#16#)) OR
 					(reg_q188 AND symb_decoder(16#29#)) OR
 					(reg_q188 AND symb_decoder(16#8f#)) OR
 					(reg_q188 AND symb_decoder(16#db#)) OR
 					(reg_q188 AND symb_decoder(16#d5#)) OR
 					(reg_q188 AND symb_decoder(16#5a#)) OR
 					(reg_q188 AND symb_decoder(16#9c#)) OR
 					(reg_q188 AND symb_decoder(16#d2#)) OR
 					(reg_q188 AND symb_decoder(16#03#)) OR
 					(reg_q188 AND symb_decoder(16#18#)) OR
 					(reg_q188 AND symb_decoder(16#1f#)) OR
 					(reg_q188 AND symb_decoder(16#87#)) OR
 					(reg_q188 AND symb_decoder(16#fe#)) OR
 					(reg_q188 AND symb_decoder(16#5f#)) OR
 					(reg_q188 AND symb_decoder(16#f9#)) OR
 					(reg_q188 AND symb_decoder(16#20#)) OR
 					(reg_q188 AND symb_decoder(16#2f#)) OR
 					(reg_q188 AND symb_decoder(16#36#)) OR
 					(reg_q188 AND symb_decoder(16#a0#)) OR
 					(reg_q188 AND symb_decoder(16#ff#)) OR
 					(reg_q188 AND symb_decoder(16#85#)) OR
 					(reg_q188 AND symb_decoder(16#b6#)) OR
 					(reg_q188 AND symb_decoder(16#1b#)) OR
 					(reg_q188 AND symb_decoder(16#72#)) OR
 					(reg_q188 AND symb_decoder(16#cb#)) OR
 					(reg_q188 AND symb_decoder(16#01#)) OR
 					(reg_q188 AND symb_decoder(16#6c#)) OR
 					(reg_q188 AND symb_decoder(16#a7#)) OR
 					(reg_q188 AND symb_decoder(16#94#)) OR
 					(reg_q188 AND symb_decoder(16#a9#)) OR
 					(reg_q188 AND symb_decoder(16#91#)) OR
 					(reg_q188 AND symb_decoder(16#32#)) OR
 					(reg_q188 AND symb_decoder(16#7a#)) OR
 					(reg_q188 AND symb_decoder(16#ba#)) OR
 					(reg_q188 AND symb_decoder(16#68#)) OR
 					(reg_q188 AND symb_decoder(16#cc#)) OR
 					(reg_q188 AND symb_decoder(16#8c#)) OR
 					(reg_q188 AND symb_decoder(16#3d#)) OR
 					(reg_q188 AND symb_decoder(16#26#)) OR
 					(reg_q188 AND symb_decoder(16#a4#)) OR
 					(reg_q188 AND symb_decoder(16#e3#)) OR
 					(reg_q188 AND symb_decoder(16#c6#)) OR
 					(reg_q188 AND symb_decoder(16#fa#)) OR
 					(reg_q188 AND symb_decoder(16#60#)) OR
 					(reg_q188 AND symb_decoder(16#f3#)) OR
 					(reg_q188 AND symb_decoder(16#57#)) OR
 					(reg_q188 AND symb_decoder(16#84#)) OR
 					(reg_q188 AND symb_decoder(16#5c#)) OR
 					(reg_q188 AND symb_decoder(16#67#)) OR
 					(reg_q188 AND symb_decoder(16#6f#)) OR
 					(reg_q188 AND symb_decoder(16#11#)) OR
 					(reg_q188 AND symb_decoder(16#3c#)) OR
 					(reg_q188 AND symb_decoder(16#b9#)) OR
 					(reg_q188 AND symb_decoder(16#47#)) OR
 					(reg_q188 AND symb_decoder(16#90#)) OR
 					(reg_q188 AND symb_decoder(16#22#)) OR
 					(reg_q188 AND symb_decoder(16#00#)) OR
 					(reg_q188 AND symb_decoder(16#42#)) OR
 					(reg_q188 AND symb_decoder(16#24#)) OR
 					(reg_q188 AND symb_decoder(16#1c#)) OR
 					(reg_q188 AND symb_decoder(16#3a#)) OR
 					(reg_q188 AND symb_decoder(16#a5#)) OR
 					(reg_q188 AND symb_decoder(16#4c#)) OR
 					(reg_q188 AND symb_decoder(16#93#)) OR
 					(reg_q188 AND symb_decoder(16#ac#)) OR
 					(reg_q188 AND symb_decoder(16#48#)) OR
 					(reg_q188 AND symb_decoder(16#fc#)) OR
 					(reg_q188 AND symb_decoder(16#82#)) OR
 					(reg_q188 AND symb_decoder(16#d7#)) OR
 					(reg_q188 AND symb_decoder(16#8b#)) OR
 					(reg_q188 AND symb_decoder(16#9e#)) OR
 					(reg_q188 AND symb_decoder(16#f7#)) OR
 					(reg_q188 AND symb_decoder(16#1d#)) OR
 					(reg_q188 AND symb_decoder(16#69#)) OR
 					(reg_q188 AND symb_decoder(16#9b#)) OR
 					(reg_q188 AND symb_decoder(16#50#)) OR
 					(reg_q188 AND symb_decoder(16#04#)) OR
 					(reg_q188 AND symb_decoder(16#7c#)) OR
 					(reg_q188 AND symb_decoder(16#25#)) OR
 					(reg_q188 AND symb_decoder(16#35#)) OR
 					(reg_q188 AND symb_decoder(16#45#)) OR
 					(reg_q188 AND symb_decoder(16#64#)) OR
 					(reg_q188 AND symb_decoder(16#a2#)) OR
 					(reg_q188 AND symb_decoder(16#e5#)) OR
 					(reg_q188 AND symb_decoder(16#75#)) OR
 					(reg_q188 AND symb_decoder(16#8d#)) OR
 					(reg_q188 AND symb_decoder(16#7f#)) OR
 					(reg_q188 AND symb_decoder(16#ca#)) OR
 					(reg_q188 AND symb_decoder(16#ad#)) OR
 					(reg_q188 AND symb_decoder(16#2d#)) OR
 					(reg_q188 AND symb_decoder(16#31#)) OR
 					(reg_q188 AND symb_decoder(16#fd#)) OR
 					(reg_q188 AND symb_decoder(16#c5#)) OR
 					(reg_q188 AND symb_decoder(16#34#)) OR
 					(reg_q188 AND symb_decoder(16#71#)) OR
 					(reg_q188 AND symb_decoder(16#89#)) OR
 					(reg_q188 AND symb_decoder(16#e1#)) OR
 					(reg_q188 AND symb_decoder(16#0f#)) OR
 					(reg_q188 AND symb_decoder(16#49#)) OR
 					(reg_q188 AND symb_decoder(16#a8#)) OR
 					(reg_q188 AND symb_decoder(16#4b#)) OR
 					(reg_q188 AND symb_decoder(16#19#)) OR
 					(reg_q188 AND symb_decoder(16#9d#)) OR
 					(reg_q188 AND symb_decoder(16#28#)) OR
 					(reg_q188 AND symb_decoder(16#f5#)) OR
 					(reg_q188 AND symb_decoder(16#06#)) OR
 					(reg_q188 AND symb_decoder(16#ea#)) OR
 					(reg_q188 AND symb_decoder(16#98#)) OR
 					(reg_q188 AND symb_decoder(16#3f#)) OR
 					(reg_q188 AND symb_decoder(16#b4#)) OR
 					(reg_q188 AND symb_decoder(16#c7#)) OR
 					(reg_q188 AND symb_decoder(16#df#)) OR
 					(reg_q188 AND symb_decoder(16#51#)) OR
 					(reg_q188 AND symb_decoder(16#0e#)) OR
 					(reg_q188 AND symb_decoder(16#5d#)) OR
 					(reg_q188 AND symb_decoder(16#74#)) OR
 					(reg_q188 AND symb_decoder(16#21#)) OR
 					(reg_q188 AND symb_decoder(16#79#)) OR
 					(reg_q188 AND symb_decoder(16#bf#)) OR
 					(reg_q188 AND symb_decoder(16#53#)) OR
 					(reg_q188 AND symb_decoder(16#40#)) OR
 					(reg_q188 AND symb_decoder(16#52#)) OR
 					(reg_q188 AND symb_decoder(16#3e#)) OR
 					(reg_q188 AND symb_decoder(16#70#)) OR
 					(reg_q188 AND symb_decoder(16#dc#)) OR
 					(reg_q188 AND symb_decoder(16#95#)) OR
 					(reg_q188 AND symb_decoder(16#bd#)) OR
 					(reg_q188 AND symb_decoder(16#d8#)) OR
 					(reg_q188 AND symb_decoder(16#ed#)) OR
 					(reg_q188 AND symb_decoder(16#73#)) OR
 					(reg_q188 AND symb_decoder(16#d9#)) OR
 					(reg_q188 AND symb_decoder(16#12#)) OR
 					(reg_q188 AND symb_decoder(16#bc#)) OR
 					(reg_q188 AND symb_decoder(16#f2#)) OR
 					(reg_q188 AND symb_decoder(16#d4#)) OR
 					(reg_q188 AND symb_decoder(16#09#)) OR
 					(reg_q188 AND symb_decoder(16#e6#)) OR
 					(reg_q188 AND symb_decoder(16#92#)) OR
 					(reg_q188 AND symb_decoder(16#c1#)) OR
 					(reg_q188 AND symb_decoder(16#17#)) OR
 					(reg_q188 AND symb_decoder(16#c8#)) OR
 					(reg_q188 AND symb_decoder(16#13#)) OR
 					(reg_q188 AND symb_decoder(16#86#)) OR
 					(reg_q188 AND symb_decoder(16#08#)) OR
 					(reg_q188 AND symb_decoder(16#61#)) OR
 					(reg_q188 AND symb_decoder(16#6e#)) OR
 					(reg_q188 AND symb_decoder(16#80#)) OR
 					(reg_q188 AND symb_decoder(16#bb#)) OR
 					(reg_q188 AND symb_decoder(16#cf#)) OR
 					(reg_q188 AND symb_decoder(16#c9#)) OR
 					(reg_q188 AND symb_decoder(16#05#)) OR
 					(reg_q188 AND symb_decoder(16#aa#)) OR
 					(reg_q188 AND symb_decoder(16#4a#)) OR
 					(reg_q188 AND symb_decoder(16#c0#)) OR
 					(reg_q188 AND symb_decoder(16#de#)) OR
 					(reg_q188 AND symb_decoder(16#99#)) OR
 					(reg_q188 AND symb_decoder(16#88#)) OR
 					(reg_q188 AND symb_decoder(16#f8#)) OR
 					(reg_q188 AND symb_decoder(16#1a#));
reg_q188_init <= '0' ;
	p_reg_q188: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q188 <= reg_q188_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q188 <= reg_q188_init;
        else
          reg_q188 <= reg_q188_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1816_in <= (reg_q2757 AND symb_decoder(16#52#)) OR
 					(reg_q2757 AND symb_decoder(16#d0#)) OR
 					(reg_q2757 AND symb_decoder(16#71#)) OR
 					(reg_q2757 AND symb_decoder(16#56#)) OR
 					(reg_q2757 AND symb_decoder(16#44#)) OR
 					(reg_q2757 AND symb_decoder(16#47#)) OR
 					(reg_q2757 AND symb_decoder(16#bf#)) OR
 					(reg_q2757 AND symb_decoder(16#40#)) OR
 					(reg_q2757 AND symb_decoder(16#b6#)) OR
 					(reg_q2757 AND symb_decoder(16#ea#)) OR
 					(reg_q2757 AND symb_decoder(16#86#)) OR
 					(reg_q2757 AND symb_decoder(16#2d#)) OR
 					(reg_q2757 AND symb_decoder(16#fc#)) OR
 					(reg_q2757 AND symb_decoder(16#5a#)) OR
 					(reg_q2757 AND symb_decoder(16#4c#)) OR
 					(reg_q2757 AND symb_decoder(16#46#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#01#)) OR
 					(reg_q2757 AND symb_decoder(16#db#)) OR
 					(reg_q2757 AND symb_decoder(16#72#)) OR
 					(reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q2757 AND symb_decoder(16#85#)) OR
 					(reg_q2757 AND symb_decoder(16#b7#)) OR
 					(reg_q2757 AND symb_decoder(16#02#)) OR
 					(reg_q2757 AND symb_decoder(16#28#)) OR
 					(reg_q2757 AND symb_decoder(16#4d#)) OR
 					(reg_q2757 AND symb_decoder(16#9b#)) OR
 					(reg_q2757 AND symb_decoder(16#7e#)) OR
 					(reg_q2757 AND symb_decoder(16#eb#)) OR
 					(reg_q2757 AND symb_decoder(16#a0#)) OR
 					(reg_q2757 AND symb_decoder(16#5b#)) OR
 					(reg_q2757 AND symb_decoder(16#8c#)) OR
 					(reg_q2757 AND symb_decoder(16#cf#)) OR
 					(reg_q2757 AND symb_decoder(16#5c#)) OR
 					(reg_q2757 AND symb_decoder(16#70#)) OR
 					(reg_q2757 AND symb_decoder(16#9d#)) OR
 					(reg_q2757 AND symb_decoder(16#84#)) OR
 					(reg_q2757 AND symb_decoder(16#f6#)) OR
 					(reg_q2757 AND symb_decoder(16#f8#)) OR
 					(reg_q2757 AND symb_decoder(16#27#)) OR
 					(reg_q2757 AND symb_decoder(16#af#)) OR
 					(reg_q2757 AND symb_decoder(16#39#)) OR
 					(reg_q2757 AND symb_decoder(16#91#)) OR
 					(reg_q2757 AND symb_decoder(16#9e#)) OR
 					(reg_q2757 AND symb_decoder(16#d5#)) OR
 					(reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#2c#)) OR
 					(reg_q2757 AND symb_decoder(16#5f#)) OR
 					(reg_q2757 AND symb_decoder(16#97#)) OR
 					(reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2757 AND symb_decoder(16#92#)) OR
 					(reg_q2757 AND symb_decoder(16#f2#)) OR
 					(reg_q2757 AND symb_decoder(16#68#)) OR
 					(reg_q2757 AND symb_decoder(16#d8#)) OR
 					(reg_q2757 AND symb_decoder(16#6e#)) OR
 					(reg_q2757 AND symb_decoder(16#50#)) OR
 					(reg_q2757 AND symb_decoder(16#00#)) OR
 					(reg_q2757 AND symb_decoder(16#ed#)) OR
 					(reg_q2757 AND symb_decoder(16#15#)) OR
 					(reg_q2757 AND symb_decoder(16#a8#)) OR
 					(reg_q2757 AND symb_decoder(16#63#)) OR
 					(reg_q2757 AND symb_decoder(16#06#)) OR
 					(reg_q2757 AND symb_decoder(16#c9#)) OR
 					(reg_q2757 AND symb_decoder(16#ce#)) OR
 					(reg_q2757 AND symb_decoder(16#be#)) OR
 					(reg_q2757 AND symb_decoder(16#59#)) OR
 					(reg_q2757 AND symb_decoder(16#55#)) OR
 					(reg_q2757 AND symb_decoder(16#75#)) OR
 					(reg_q2757 AND symb_decoder(16#e8#)) OR
 					(reg_q2757 AND symb_decoder(16#04#)) OR
 					(reg_q2757 AND symb_decoder(16#e3#)) OR
 					(reg_q2757 AND symb_decoder(16#6a#)) OR
 					(reg_q2757 AND symb_decoder(16#c0#)) OR
 					(reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#67#)) OR
 					(reg_q2757 AND symb_decoder(16#d1#)) OR
 					(reg_q2757 AND symb_decoder(16#31#)) OR
 					(reg_q2757 AND symb_decoder(16#1b#)) OR
 					(reg_q2757 AND symb_decoder(16#b3#)) OR
 					(reg_q2757 AND symb_decoder(16#a9#)) OR
 					(reg_q2757 AND symb_decoder(16#ff#)) OR
 					(reg_q2757 AND symb_decoder(16#98#)) OR
 					(reg_q2757 AND symb_decoder(16#7f#)) OR
 					(reg_q2757 AND symb_decoder(16#61#)) OR
 					(reg_q2757 AND symb_decoder(16#da#)) OR
 					(reg_q2757 AND symb_decoder(16#94#)) OR
 					(reg_q2757 AND symb_decoder(16#99#)) OR
 					(reg_q2757 AND symb_decoder(16#20#)) OR
 					(reg_q2757 AND symb_decoder(16#79#)) OR
 					(reg_q2757 AND symb_decoder(16#a3#)) OR
 					(reg_q2757 AND symb_decoder(16#22#)) OR
 					(reg_q2757 AND symb_decoder(16#90#)) OR
 					(reg_q2757 AND symb_decoder(16#41#)) OR
 					(reg_q2757 AND symb_decoder(16#d6#)) OR
 					(reg_q2757 AND symb_decoder(16#df#)) OR
 					(reg_q2757 AND symb_decoder(16#b5#)) OR
 					(reg_q2757 AND symb_decoder(16#65#)) OR
 					(reg_q2757 AND symb_decoder(16#69#)) OR
 					(reg_q2757 AND symb_decoder(16#7d#)) OR
 					(reg_q2757 AND symb_decoder(16#9a#)) OR
 					(reg_q2757 AND symb_decoder(16#de#)) OR
 					(reg_q2757 AND symb_decoder(16#48#)) OR
 					(reg_q2757 AND symb_decoder(16#10#)) OR
 					(reg_q2757 AND symb_decoder(16#4e#)) OR
 					(reg_q2757 AND symb_decoder(16#8a#)) OR
 					(reg_q2757 AND symb_decoder(16#b4#)) OR
 					(reg_q2757 AND symb_decoder(16#26#)) OR
 					(reg_q2757 AND symb_decoder(16#12#)) OR
 					(reg_q2757 AND symb_decoder(16#f7#)) OR
 					(reg_q2757 AND symb_decoder(16#24#)) OR
 					(reg_q2757 AND symb_decoder(16#a1#)) OR
 					(reg_q2757 AND symb_decoder(16#7b#)) OR
 					(reg_q2757 AND symb_decoder(16#0f#)) OR
 					(reg_q2757 AND symb_decoder(16#80#)) OR
 					(reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2757 AND symb_decoder(16#07#)) OR
 					(reg_q2757 AND symb_decoder(16#c8#)) OR
 					(reg_q2757 AND symb_decoder(16#3f#)) OR
 					(reg_q2757 AND symb_decoder(16#e7#)) OR
 					(reg_q2757 AND symb_decoder(16#93#)) OR
 					(reg_q2757 AND symb_decoder(16#58#)) OR
 					(reg_q2757 AND symb_decoder(16#8f#)) OR
 					(reg_q2757 AND symb_decoder(16#cb#)) OR
 					(reg_q2757 AND symb_decoder(16#b2#)) OR
 					(reg_q2757 AND symb_decoder(16#64#)) OR
 					(reg_q2757 AND symb_decoder(16#e2#)) OR
 					(reg_q2757 AND symb_decoder(16#36#)) OR
 					(reg_q2757 AND symb_decoder(16#25#)) OR
 					(reg_q2757 AND symb_decoder(16#a2#)) OR
 					(reg_q2757 AND symb_decoder(16#b9#)) OR
 					(reg_q2757 AND symb_decoder(16#fb#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q2757 AND symb_decoder(16#bc#)) OR
 					(reg_q2757 AND symb_decoder(16#23#)) OR
 					(reg_q2757 AND symb_decoder(16#fa#)) OR
 					(reg_q2757 AND symb_decoder(16#1a#)) OR
 					(reg_q2757 AND symb_decoder(16#2e#)) OR
 					(reg_q2757 AND symb_decoder(16#09#)) OR
 					(reg_q2757 AND symb_decoder(16#11#)) OR
 					(reg_q2757 AND symb_decoder(16#ec#)) OR
 					(reg_q2757 AND symb_decoder(16#d9#)) OR
 					(reg_q2757 AND symb_decoder(16#74#)) OR
 					(reg_q2757 AND symb_decoder(16#5d#)) OR
 					(reg_q2757 AND symb_decoder(16#7a#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q2757 AND symb_decoder(16#17#)) OR
 					(reg_q2757 AND symb_decoder(16#88#)) OR
 					(reg_q2757 AND symb_decoder(16#e0#)) OR
 					(reg_q2757 AND symb_decoder(16#fd#)) OR
 					(reg_q2757 AND symb_decoder(16#ae#)) OR
 					(reg_q2757 AND symb_decoder(16#83#)) OR
 					(reg_q2757 AND symb_decoder(16#13#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#8d#)) OR
 					(reg_q2757 AND symb_decoder(16#f3#)) OR
 					(reg_q2757 AND symb_decoder(16#95#)) OR
 					(reg_q2757 AND symb_decoder(16#dc#)) OR
 					(reg_q2757 AND symb_decoder(16#76#)) OR
 					(reg_q2757 AND symb_decoder(16#34#)) OR
 					(reg_q2757 AND symb_decoder(16#03#)) OR
 					(reg_q2757 AND symb_decoder(16#0e#)) OR
 					(reg_q2757 AND symb_decoder(16#21#)) OR
 					(reg_q2757 AND symb_decoder(16#42#)) OR
 					(reg_q2757 AND symb_decoder(16#d2#)) OR
 					(reg_q2757 AND symb_decoder(16#82#)) OR
 					(reg_q2757 AND symb_decoder(16#60#)) OR
 					(reg_q2757 AND symb_decoder(16#37#)) OR
 					(reg_q2757 AND symb_decoder(16#3a#)) OR
 					(reg_q2757 AND symb_decoder(16#66#)) OR
 					(reg_q2757 AND symb_decoder(16#cc#)) OR
 					(reg_q2757 AND symb_decoder(16#45#)) OR
 					(reg_q2757 AND symb_decoder(16#e1#)) OR
 					(reg_q2757 AND symb_decoder(16#c4#)) OR
 					(reg_q2757 AND symb_decoder(16#b1#)) OR
 					(reg_q2757 AND symb_decoder(16#0b#)) OR
 					(reg_q2757 AND symb_decoder(16#8e#)) OR
 					(reg_q2757 AND symb_decoder(16#ba#)) OR
 					(reg_q2757 AND symb_decoder(16#ac#)) OR
 					(reg_q2757 AND symb_decoder(16#4f#)) OR
 					(reg_q2757 AND symb_decoder(16#3e#)) OR
 					(reg_q2757 AND symb_decoder(16#32#)) OR
 					(reg_q2757 AND symb_decoder(16#19#)) OR
 					(reg_q2757 AND symb_decoder(16#d7#)) OR
 					(reg_q2757 AND symb_decoder(16#5e#)) OR
 					(reg_q2757 AND symb_decoder(16#87#)) OR
 					(reg_q2757 AND symb_decoder(16#35#)) OR
 					(reg_q2757 AND symb_decoder(16#7c#)) OR
 					(reg_q2757 AND symb_decoder(16#f1#)) OR
 					(reg_q2757 AND symb_decoder(16#6d#)) OR
 					(reg_q2757 AND symb_decoder(16#4b#)) OR
 					(reg_q2757 AND symb_decoder(16#a7#)) OR
 					(reg_q2757 AND symb_decoder(16#78#)) OR
 					(reg_q2757 AND symb_decoder(16#6c#)) OR
 					(reg_q2757 AND symb_decoder(16#30#)) OR
 					(reg_q2757 AND symb_decoder(16#b8#)) OR
 					(reg_q2757 AND symb_decoder(16#0c#)) OR
 					(reg_q2757 AND symb_decoder(16#d4#)) OR
 					(reg_q2757 AND symb_decoder(16#e4#)) OR
 					(reg_q2757 AND symb_decoder(16#08#)) OR
 					(reg_q2757 AND symb_decoder(16#14#)) OR
 					(reg_q2757 AND symb_decoder(16#c6#)) OR
 					(reg_q2757 AND symb_decoder(16#6f#)) OR
 					(reg_q2757 AND symb_decoder(16#51#)) OR
 					(reg_q2757 AND symb_decoder(16#c5#)) OR
 					(reg_q2757 AND symb_decoder(16#bd#)) OR
 					(reg_q2757 AND symb_decoder(16#3b#)) OR
 					(reg_q2757 AND symb_decoder(16#81#)) OR
 					(reg_q2757 AND symb_decoder(16#b0#)) OR
 					(reg_q2757 AND symb_decoder(16#33#)) OR
 					(reg_q2757 AND symb_decoder(16#8b#)) OR
 					(reg_q2757 AND symb_decoder(16#16#)) OR
 					(reg_q2757 AND symb_decoder(16#c7#)) OR
 					(reg_q2757 AND symb_decoder(16#c3#)) OR
 					(reg_q2757 AND symb_decoder(16#1d#)) OR
 					(reg_q2757 AND symb_decoder(16#ab#)) OR
 					(reg_q2757 AND symb_decoder(16#bb#)) OR
 					(reg_q2757 AND symb_decoder(16#2b#)) OR
 					(reg_q2757 AND symb_decoder(16#3d#)) OR
 					(reg_q2757 AND symb_decoder(16#ad#)) OR
 					(reg_q2757 AND symb_decoder(16#1c#)) OR
 					(reg_q2757 AND symb_decoder(16#e9#)) OR
 					(reg_q2757 AND symb_decoder(16#49#)) OR
 					(reg_q2757 AND symb_decoder(16#fe#)) OR
 					(reg_q2757 AND symb_decoder(16#cd#)) OR
 					(reg_q2757 AND symb_decoder(16#a4#)) OR
 					(reg_q2757 AND symb_decoder(16#d3#)) OR
 					(reg_q2757 AND symb_decoder(16#1e#)) OR
 					(reg_q2757 AND symb_decoder(16#e6#)) OR
 					(reg_q2757 AND symb_decoder(16#ca#)) OR
 					(reg_q2757 AND symb_decoder(16#a5#)) OR
 					(reg_q2757 AND symb_decoder(16#62#)) OR
 					(reg_q2757 AND symb_decoder(16#2a#)) OR
 					(reg_q2757 AND symb_decoder(16#89#)) OR
 					(reg_q2757 AND symb_decoder(16#ef#)) OR
 					(reg_q2757 AND symb_decoder(16#f5#)) OR
 					(reg_q2757 AND symb_decoder(16#43#)) OR
 					(reg_q2757 AND symb_decoder(16#c1#)) OR
 					(reg_q2757 AND symb_decoder(16#9f#)) OR
 					(reg_q2757 AND symb_decoder(16#c2#)) OR
 					(reg_q2757 AND symb_decoder(16#6b#)) OR
 					(reg_q2757 AND symb_decoder(16#96#)) OR
 					(reg_q2757 AND symb_decoder(16#ee#)) OR
 					(reg_q2757 AND symb_decoder(16#29#)) OR
 					(reg_q2757 AND symb_decoder(16#dd#)) OR
 					(reg_q2757 AND symb_decoder(16#9c#)) OR
 					(reg_q2757 AND symb_decoder(16#4a#)) OR
 					(reg_q2757 AND symb_decoder(16#1f#)) OR
 					(reg_q2757 AND symb_decoder(16#e5#)) OR
 					(reg_q2757 AND symb_decoder(16#aa#)) OR
 					(reg_q2757 AND symb_decoder(16#05#)) OR
 					(reg_q2757 AND symb_decoder(16#f9#)) OR
 					(reg_q2757 AND symb_decoder(16#18#)) OR
 					(reg_q2757 AND symb_decoder(16#f4#)) OR
 					(reg_q2757 AND symb_decoder(16#38#)) OR
 					(reg_q2757 AND symb_decoder(16#a6#)) OR
 					(reg_q2757 AND symb_decoder(16#f0#)) OR
 					(reg_q1816 AND symb_decoder(16#ec#)) OR
 					(reg_q1816 AND symb_decoder(16#1c#)) OR
 					(reg_q1816 AND symb_decoder(16#89#)) OR
 					(reg_q1816 AND symb_decoder(16#d0#)) OR
 					(reg_q1816 AND symb_decoder(16#19#)) OR
 					(reg_q1816 AND symb_decoder(16#6f#)) OR
 					(reg_q1816 AND symb_decoder(16#7f#)) OR
 					(reg_q1816 AND symb_decoder(16#f4#)) OR
 					(reg_q1816 AND symb_decoder(16#18#)) OR
 					(reg_q1816 AND symb_decoder(16#3b#)) OR
 					(reg_q1816 AND symb_decoder(16#84#)) OR
 					(reg_q1816 AND symb_decoder(16#45#)) OR
 					(reg_q1816 AND symb_decoder(16#29#)) OR
 					(reg_q1816 AND symb_decoder(16#e7#)) OR
 					(reg_q1816 AND symb_decoder(16#33#)) OR
 					(reg_q1816 AND symb_decoder(16#72#)) OR
 					(reg_q1816 AND symb_decoder(16#d2#)) OR
 					(reg_q1816 AND symb_decoder(16#d5#)) OR
 					(reg_q1816 AND symb_decoder(16#35#)) OR
 					(reg_q1816 AND symb_decoder(16#e0#)) OR
 					(reg_q1816 AND symb_decoder(16#c0#)) OR
 					(reg_q1816 AND symb_decoder(16#37#)) OR
 					(reg_q1816 AND symb_decoder(16#de#)) OR
 					(reg_q1816 AND symb_decoder(16#bc#)) OR
 					(reg_q1816 AND symb_decoder(16#56#)) OR
 					(reg_q1816 AND symb_decoder(16#c3#)) OR
 					(reg_q1816 AND symb_decoder(16#96#)) OR
 					(reg_q1816 AND symb_decoder(16#0c#)) OR
 					(reg_q1816 AND symb_decoder(16#5e#)) OR
 					(reg_q1816 AND symb_decoder(16#63#)) OR
 					(reg_q1816 AND symb_decoder(16#12#)) OR
 					(reg_q1816 AND symb_decoder(16#d8#)) OR
 					(reg_q1816 AND symb_decoder(16#dd#)) OR
 					(reg_q1816 AND symb_decoder(16#bd#)) OR
 					(reg_q1816 AND symb_decoder(16#e1#)) OR
 					(reg_q1816 AND symb_decoder(16#1f#)) OR
 					(reg_q1816 AND symb_decoder(16#a8#)) OR
 					(reg_q1816 AND symb_decoder(16#06#)) OR
 					(reg_q1816 AND symb_decoder(16#8f#)) OR
 					(reg_q1816 AND symb_decoder(16#47#)) OR
 					(reg_q1816 AND symb_decoder(16#ac#)) OR
 					(reg_q1816 AND symb_decoder(16#6e#)) OR
 					(reg_q1816 AND symb_decoder(16#59#)) OR
 					(reg_q1816 AND symb_decoder(16#3f#)) OR
 					(reg_q1816 AND symb_decoder(16#42#)) OR
 					(reg_q1816 AND symb_decoder(16#8e#)) OR
 					(reg_q1816 AND symb_decoder(16#e8#)) OR
 					(reg_q1816 AND symb_decoder(16#46#)) OR
 					(reg_q1816 AND symb_decoder(16#61#)) OR
 					(reg_q1816 AND symb_decoder(16#80#)) OR
 					(reg_q1816 AND symb_decoder(16#08#)) OR
 					(reg_q1816 AND symb_decoder(16#39#)) OR
 					(reg_q1816 AND symb_decoder(16#6a#)) OR
 					(reg_q1816 AND symb_decoder(16#cb#)) OR
 					(reg_q1816 AND symb_decoder(16#62#)) OR
 					(reg_q1816 AND symb_decoder(16#6b#)) OR
 					(reg_q1816 AND symb_decoder(16#1e#)) OR
 					(reg_q1816 AND symb_decoder(16#5f#)) OR
 					(reg_q1816 AND symb_decoder(16#66#)) OR
 					(reg_q1816 AND symb_decoder(16#1b#)) OR
 					(reg_q1816 AND symb_decoder(16#50#)) OR
 					(reg_q1816 AND symb_decoder(16#1a#)) OR
 					(reg_q1816 AND symb_decoder(16#fe#)) OR
 					(reg_q1816 AND symb_decoder(16#ad#)) OR
 					(reg_q1816 AND symb_decoder(16#94#)) OR
 					(reg_q1816 AND symb_decoder(16#05#)) OR
 					(reg_q1816 AND symb_decoder(16#9b#)) OR
 					(reg_q1816 AND symb_decoder(16#5c#)) OR
 					(reg_q1816 AND symb_decoder(16#8b#)) OR
 					(reg_q1816 AND symb_decoder(16#14#)) OR
 					(reg_q1816 AND symb_decoder(16#b1#)) OR
 					(reg_q1816 AND symb_decoder(16#34#)) OR
 					(reg_q1816 AND symb_decoder(16#4b#)) OR
 					(reg_q1816 AND symb_decoder(16#7a#)) OR
 					(reg_q1816 AND symb_decoder(16#81#)) OR
 					(reg_q1816 AND symb_decoder(16#2b#)) OR
 					(reg_q1816 AND symb_decoder(16#70#)) OR
 					(reg_q1816 AND symb_decoder(16#60#)) OR
 					(reg_q1816 AND symb_decoder(16#00#)) OR
 					(reg_q1816 AND symb_decoder(16#17#)) OR
 					(reg_q1816 AND symb_decoder(16#c9#)) OR
 					(reg_q1816 AND symb_decoder(16#15#)) OR
 					(reg_q1816 AND symb_decoder(16#aa#)) OR
 					(reg_q1816 AND symb_decoder(16#f8#)) OR
 					(reg_q1816 AND symb_decoder(16#4a#)) OR
 					(reg_q1816 AND symb_decoder(16#13#)) OR
 					(reg_q1816 AND symb_decoder(16#31#)) OR
 					(reg_q1816 AND symb_decoder(16#48#)) OR
 					(reg_q1816 AND symb_decoder(16#3d#)) OR
 					(reg_q1816 AND symb_decoder(16#75#)) OR
 					(reg_q1816 AND symb_decoder(16#69#)) OR
 					(reg_q1816 AND symb_decoder(16#d3#)) OR
 					(reg_q1816 AND symb_decoder(16#bf#)) OR
 					(reg_q1816 AND symb_decoder(16#78#)) OR
 					(reg_q1816 AND symb_decoder(16#e2#)) OR
 					(reg_q1816 AND symb_decoder(16#e6#)) OR
 					(reg_q1816 AND symb_decoder(16#3c#)) OR
 					(reg_q1816 AND symb_decoder(16#dc#)) OR
 					(reg_q1816 AND symb_decoder(16#10#)) OR
 					(reg_q1816 AND symb_decoder(16#88#)) OR
 					(reg_q1816 AND symb_decoder(16#65#)) OR
 					(reg_q1816 AND symb_decoder(16#d7#)) OR
 					(reg_q1816 AND symb_decoder(16#a6#)) OR
 					(reg_q1816 AND symb_decoder(16#76#)) OR
 					(reg_q1816 AND symb_decoder(16#fc#)) OR
 					(reg_q1816 AND symb_decoder(16#a0#)) OR
 					(reg_q1816 AND symb_decoder(16#07#)) OR
 					(reg_q1816 AND symb_decoder(16#a7#)) OR
 					(reg_q1816 AND symb_decoder(16#57#)) OR
 					(reg_q1816 AND symb_decoder(16#fd#)) OR
 					(reg_q1816 AND symb_decoder(16#52#)) OR
 					(reg_q1816 AND symb_decoder(16#a3#)) OR
 					(reg_q1816 AND symb_decoder(16#22#)) OR
 					(reg_q1816 AND symb_decoder(16#2e#)) OR
 					(reg_q1816 AND symb_decoder(16#5d#)) OR
 					(reg_q1816 AND symb_decoder(16#d4#)) OR
 					(reg_q1816 AND symb_decoder(16#0d#)) OR
 					(reg_q1816 AND symb_decoder(16#f6#)) OR
 					(reg_q1816 AND symb_decoder(16#74#)) OR
 					(reg_q1816 AND symb_decoder(16#16#)) OR
 					(reg_q1816 AND symb_decoder(16#eb#)) OR
 					(reg_q1816 AND symb_decoder(16#f2#)) OR
 					(reg_q1816 AND symb_decoder(16#ae#)) OR
 					(reg_q1816 AND symb_decoder(16#20#)) OR
 					(reg_q1816 AND symb_decoder(16#91#)) OR
 					(reg_q1816 AND symb_decoder(16#01#)) OR
 					(reg_q1816 AND symb_decoder(16#23#)) OR
 					(reg_q1816 AND symb_decoder(16#4d#)) OR
 					(reg_q1816 AND symb_decoder(16#40#)) OR
 					(reg_q1816 AND symb_decoder(16#32#)) OR
 					(reg_q1816 AND symb_decoder(16#b7#)) OR
 					(reg_q1816 AND symb_decoder(16#98#)) OR
 					(reg_q1816 AND symb_decoder(16#c5#)) OR
 					(reg_q1816 AND symb_decoder(16#be#)) OR
 					(reg_q1816 AND symb_decoder(16#cc#)) OR
 					(reg_q1816 AND symb_decoder(16#25#)) OR
 					(reg_q1816 AND symb_decoder(16#cf#)) OR
 					(reg_q1816 AND symb_decoder(16#a4#)) OR
 					(reg_q1816 AND symb_decoder(16#73#)) OR
 					(reg_q1816 AND symb_decoder(16#ab#)) OR
 					(reg_q1816 AND symb_decoder(16#9c#)) OR
 					(reg_q1816 AND symb_decoder(16#83#)) OR
 					(reg_q1816 AND symb_decoder(16#21#)) OR
 					(reg_q1816 AND symb_decoder(16#41#)) OR
 					(reg_q1816 AND symb_decoder(16#49#)) OR
 					(reg_q1816 AND symb_decoder(16#a9#)) OR
 					(reg_q1816 AND symb_decoder(16#f5#)) OR
 					(reg_q1816 AND symb_decoder(16#ed#)) OR
 					(reg_q1816 AND symb_decoder(16#68#)) OR
 					(reg_q1816 AND symb_decoder(16#3e#)) OR
 					(reg_q1816 AND symb_decoder(16#26#)) OR
 					(reg_q1816 AND symb_decoder(16#c4#)) OR
 					(reg_q1816 AND symb_decoder(16#6d#)) OR
 					(reg_q1816 AND symb_decoder(16#7b#)) OR
 					(reg_q1816 AND symb_decoder(16#64#)) OR
 					(reg_q1816 AND symb_decoder(16#e5#)) OR
 					(reg_q1816 AND symb_decoder(16#7d#)) OR
 					(reg_q1816 AND symb_decoder(16#b3#)) OR
 					(reg_q1816 AND symb_decoder(16#a1#)) OR
 					(reg_q1816 AND symb_decoder(16#d1#)) OR
 					(reg_q1816 AND symb_decoder(16#55#)) OR
 					(reg_q1816 AND symb_decoder(16#77#)) OR
 					(reg_q1816 AND symb_decoder(16#04#)) OR
 					(reg_q1816 AND symb_decoder(16#2c#)) OR
 					(reg_q1816 AND symb_decoder(16#f1#)) OR
 					(reg_q1816 AND symb_decoder(16#9e#)) OR
 					(reg_q1816 AND symb_decoder(16#fa#)) OR
 					(reg_q1816 AND symb_decoder(16#1d#)) OR
 					(reg_q1816 AND symb_decoder(16#b0#)) OR
 					(reg_q1816 AND symb_decoder(16#ca#)) OR
 					(reg_q1816 AND symb_decoder(16#ea#)) OR
 					(reg_q1816 AND symb_decoder(16#82#)) OR
 					(reg_q1816 AND symb_decoder(16#9f#)) OR
 					(reg_q1816 AND symb_decoder(16#51#)) OR
 					(reg_q1816 AND symb_decoder(16#71#)) OR
 					(reg_q1816 AND symb_decoder(16#9a#)) OR
 					(reg_q1816 AND symb_decoder(16#0a#)) OR
 					(reg_q1816 AND symb_decoder(16#5a#)) OR
 					(reg_q1816 AND symb_decoder(16#79#)) OR
 					(reg_q1816 AND symb_decoder(16#db#)) OR
 					(reg_q1816 AND symb_decoder(16#95#)) OR
 					(reg_q1816 AND symb_decoder(16#e4#)) OR
 					(reg_q1816 AND symb_decoder(16#53#)) OR
 					(reg_q1816 AND symb_decoder(16#c1#)) OR
 					(reg_q1816 AND symb_decoder(16#c7#)) OR
 					(reg_q1816 AND symb_decoder(16#6c#)) OR
 					(reg_q1816 AND symb_decoder(16#bb#)) OR
 					(reg_q1816 AND symb_decoder(16#97#)) OR
 					(reg_q1816 AND symb_decoder(16#67#)) OR
 					(reg_q1816 AND symb_decoder(16#ee#)) OR
 					(reg_q1816 AND symb_decoder(16#d6#)) OR
 					(reg_q1816 AND symb_decoder(16#43#)) OR
 					(reg_q1816 AND symb_decoder(16#9d#)) OR
 					(reg_q1816 AND symb_decoder(16#09#)) OR
 					(reg_q1816 AND symb_decoder(16#c8#)) OR
 					(reg_q1816 AND symb_decoder(16#2f#)) OR
 					(reg_q1816 AND symb_decoder(16#b6#)) OR
 					(reg_q1816 AND symb_decoder(16#7c#)) OR
 					(reg_q1816 AND symb_decoder(16#a5#)) OR
 					(reg_q1816 AND symb_decoder(16#85#)) OR
 					(reg_q1816 AND symb_decoder(16#b5#)) OR
 					(reg_q1816 AND symb_decoder(16#4f#)) OR
 					(reg_q1816 AND symb_decoder(16#ff#)) OR
 					(reg_q1816 AND symb_decoder(16#03#)) OR
 					(reg_q1816 AND symb_decoder(16#4c#)) OR
 					(reg_q1816 AND symb_decoder(16#7e#)) OR
 					(reg_q1816 AND symb_decoder(16#c6#)) OR
 					(reg_q1816 AND symb_decoder(16#58#)) OR
 					(reg_q1816 AND symb_decoder(16#0f#)) OR
 					(reg_q1816 AND symb_decoder(16#f3#)) OR
 					(reg_q1816 AND symb_decoder(16#e9#)) OR
 					(reg_q1816 AND symb_decoder(16#f9#)) OR
 					(reg_q1816 AND symb_decoder(16#3a#)) OR
 					(reg_q1816 AND symb_decoder(16#0b#)) OR
 					(reg_q1816 AND symb_decoder(16#93#)) OR
 					(reg_q1816 AND symb_decoder(16#ef#)) OR
 					(reg_q1816 AND symb_decoder(16#8c#)) OR
 					(reg_q1816 AND symb_decoder(16#d9#)) OR
 					(reg_q1816 AND symb_decoder(16#11#)) OR
 					(reg_q1816 AND symb_decoder(16#99#)) OR
 					(reg_q1816 AND symb_decoder(16#30#)) OR
 					(reg_q1816 AND symb_decoder(16#ce#)) OR
 					(reg_q1816 AND symb_decoder(16#28#)) OR
 					(reg_q1816 AND symb_decoder(16#38#)) OR
 					(reg_q1816 AND symb_decoder(16#fb#)) OR
 					(reg_q1816 AND symb_decoder(16#ba#)) OR
 					(reg_q1816 AND symb_decoder(16#da#)) OR
 					(reg_q1816 AND symb_decoder(16#87#)) OR
 					(reg_q1816 AND symb_decoder(16#02#)) OR
 					(reg_q1816 AND symb_decoder(16#8d#)) OR
 					(reg_q1816 AND symb_decoder(16#f0#)) OR
 					(reg_q1816 AND symb_decoder(16#92#)) OR
 					(reg_q1816 AND symb_decoder(16#b9#)) OR
 					(reg_q1816 AND symb_decoder(16#a2#)) OR
 					(reg_q1816 AND symb_decoder(16#0e#)) OR
 					(reg_q1816 AND symb_decoder(16#27#)) OR
 					(reg_q1816 AND symb_decoder(16#c2#)) OR
 					(reg_q1816 AND symb_decoder(16#af#)) OR
 					(reg_q1816 AND symb_decoder(16#b2#)) OR
 					(reg_q1816 AND symb_decoder(16#2a#)) OR
 					(reg_q1816 AND symb_decoder(16#4e#)) OR
 					(reg_q1816 AND symb_decoder(16#2d#)) OR
 					(reg_q1816 AND symb_decoder(16#e3#)) OR
 					(reg_q1816 AND symb_decoder(16#df#)) OR
 					(reg_q1816 AND symb_decoder(16#8a#)) OR
 					(reg_q1816 AND symb_decoder(16#44#)) OR
 					(reg_q1816 AND symb_decoder(16#5b#)) OR
 					(reg_q1816 AND symb_decoder(16#b4#)) OR
 					(reg_q1816 AND symb_decoder(16#54#)) OR
 					(reg_q1816 AND symb_decoder(16#f7#)) OR
 					(reg_q1816 AND symb_decoder(16#cd#)) OR
 					(reg_q1816 AND symb_decoder(16#86#)) OR
 					(reg_q1816 AND symb_decoder(16#b8#)) OR
 					(reg_q1816 AND symb_decoder(16#90#)) OR
 					(reg_q1816 AND symb_decoder(16#36#)) OR
 					(reg_q1816 AND symb_decoder(16#24#));
reg_q1816_init <= '0' ;
	p_reg_q1816: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1816 <= reg_q1816_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1816 <= reg_q1816_init;
        else
          reg_q1816 <= reg_q1816_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph69

reg_q298_in <= (reg_q296 AND symb_decoder(16#6e#)) OR
 					(reg_q296 AND symb_decoder(16#4e#));
reg_q1620_in <= (reg_q1626 AND symb_decoder(16#69#)) OR
 					(reg_q1626 AND symb_decoder(16#49#)) OR
 					(reg_q1616 AND symb_decoder(16#49#)) OR
 					(reg_q1616 AND symb_decoder(16#69#));
reg_q288_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q286 AND symb_decoder(16#53#)) OR
 					(reg_q286 AND symb_decoder(16#73#));
reg_q2681_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2680 AND symb_decoder(16#0a#)) OR
 					(reg_q2680 AND symb_decoder(16#0d#));
reg_q1965_in <= (reg_q1961 AND symb_decoder(16#7c#)) OR
 					(reg_q1975 AND symb_decoder(16#7c#));
reg_q1630_in <= (reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q1628 AND symb_decoder(16#77#)) OR
 					(reg_q1628 AND symb_decoder(16#57#));
reg_q1361_in <= (reg_q1393 AND symb_decoder(16#66#)) OR
 					(reg_q1393 AND symb_decoder(16#46#)) OR
 					(reg_q1357 AND symb_decoder(16#46#)) OR
 					(reg_q1357 AND symb_decoder(16#66#));
reg_q1391_in <= (reg_q1389 AND symb_decoder(16#4e#)) OR
 					(reg_q1389 AND symb_decoder(16#6e#));
reg_q2058_in <= (reg_q2757 AND symb_decoder(16#2f#)) OR
 					(reg_q2056 AND symb_decoder(16#2f#));
reg_q2419_in <= (reg_q2757 AND symb_decoder(16#3c#)) OR
 					(reg_q2417 AND symb_decoder(16#3c#));
reg_q1584_in <= (reg_q1582 AND symb_decoder(16#4e#)) OR
 					(reg_q1582 AND symb_decoder(16#6e#));
reg_q1222_in <= (reg_q1220 AND symb_decoder(16#45#)) OR
 					(reg_q1220 AND symb_decoder(16#65#));
reg_q1024_in <= (reg_q2757 AND symb_decoder(16#54#)) OR
 					(reg_q1022 AND symb_decoder(16#54#));
reg_q1459_in <= (reg_q1457 AND symb_decoder(16#6e#)) OR
 					(reg_q1457 AND symb_decoder(16#4e#));
reg_q2162_in <= (reg_q2160 AND symb_decoder(16#6e#)) OR
 					(reg_q2160 AND symb_decoder(16#4e#));
reg_fullgraph69_init <= "0000";

reg_fullgraph69_sel <= "0" & reg_q2162_in & reg_q1459_in & reg_q1024_in & reg_q1222_in & reg_q1584_in & reg_q2419_in & reg_q2058_in & reg_q1391_in & reg_q1361_in & reg_q1630_in & reg_q1965_in & reg_q2681_in & reg_q288_in & reg_q1620_in & reg_q298_in;

	--coder fullgraph69
with reg_fullgraph69_sel select
reg_fullgraph69_in <=
	"0001" when "0000000000000001",
	"0010" when "0000000000000010",
	"0011" when "0000000000000100",
	"0100" when "0000000000001000",
	"0101" when "0000000000010000",
	"0110" when "0000000000100000",
	"0111" when "0000000001000000",
	"1000" when "0000000010000000",
	"1001" when "0000000100000000",
	"1010" when "0000001000000000",
	"1011" when "0000010000000000",
	"1100" when "0000100000000000",
	"1101" when "0001000000000000",
	"1110" when "0010000000000000",
	"1111" when "0100000000000000",
	"0000" when others;
 --end coder

	p_reg_fullgraph69: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph69 <= reg_fullgraph69_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph69 <= reg_fullgraph69_init;
        else
          reg_fullgraph69 <= reg_fullgraph69_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph69

		reg_q298 <= '1' when reg_fullgraph69 = "0001" else '0'; 
		reg_q1620 <= '1' when reg_fullgraph69 = "0010" else '0'; 
		reg_q288 <= '1' when reg_fullgraph69 = "0011" else '0'; 
		reg_q2681 <= '1' when reg_fullgraph69 = "0100" else '0'; 
		reg_q1965 <= '1' when reg_fullgraph69 = "0101" else '0'; 
		reg_q1630 <= '1' when reg_fullgraph69 = "0110" else '0'; 
		reg_q1361 <= '1' when reg_fullgraph69 = "0111" else '0'; 
		reg_q1391 <= '1' when reg_fullgraph69 = "1000" else '0'; 
		reg_q2058 <= '1' when reg_fullgraph69 = "1001" else '0'; 
		reg_q2419 <= '1' when reg_fullgraph69 = "1010" else '0'; 
		reg_q1584 <= '1' when reg_fullgraph69 = "1011" else '0'; 
		reg_q1222 <= '1' when reg_fullgraph69 = "1100" else '0'; 
		reg_q1024 <= '1' when reg_fullgraph69 = "1101" else '0'; 
		reg_q1459 <= '1' when reg_fullgraph69 = "1110" else '0'; 
		reg_q2162 <= '1' when reg_fullgraph69 = "1111" else '0'; 
--end decoder 
--######################################################
--fullgraph70

reg_q401_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q399 AND symb_decoder(16#53#)) OR
 					(reg_q399 AND symb_decoder(16#73#));
reg_q695_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q694 AND symb_decoder(16#0a#)) OR
 					(reg_q694 AND symb_decoder(16#0d#));
reg_q1397_in <= (reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q1395 AND symb_decoder(16#57#)) OR
 					(reg_q1395 AND symb_decoder(16#77#));
reg_q1676_in <= (reg_q1672 AND symb_decoder(16#69#)) OR
 					(reg_q1672 AND symb_decoder(16#49#)) OR
 					(reg_q1682 AND symb_decoder(16#69#)) OR
 					(reg_q1682 AND symb_decoder(16#49#));
reg_q2154_in <= (reg_q2216 AND symb_decoder(16#46#)) OR
 					(reg_q2216 AND symb_decoder(16#66#)) OR
 					(reg_q2150 AND symb_decoder(16#66#)) OR
 					(reg_q2150 AND symb_decoder(16#46#));
reg_q2550_in <= (reg_q2548 AND symb_decoder(16#3c#));
reg_q2505_in <= (reg_q2503 AND symb_decoder(16#2f#));
reg_q2655_in <= (reg_q2651 AND symb_decoder(16#7c#)) OR
 					(reg_q2677 AND symb_decoder(16#7c#));
reg_q2503_in <= (reg_q2501 AND symb_decoder(16#3c#));
reg_q1652_in <= (reg_q1650 AND symb_decoder(16#2f#));
reg_fullgraph70_init <= "0000";

reg_fullgraph70_sel <= "000000" & reg_q1652_in & reg_q2503_in & reg_q2655_in & reg_q2505_in & reg_q2550_in & reg_q2154_in & reg_q1676_in & reg_q1397_in & reg_q695_in & reg_q401_in;

	--coder fullgraph70
with reg_fullgraph70_sel select
reg_fullgraph70_in <=
	"0001" when "0000000000000001",
	"0010" when "0000000000000010",
	"0011" when "0000000000000100",
	"0100" when "0000000000001000",
	"0101" when "0000000000010000",
	"0110" when "0000000000100000",
	"0111" when "0000000001000000",
	"1000" when "0000000010000000",
	"1001" when "0000000100000000",
	"1010" when "0000001000000000",
	"0000" when others;
 --end coder

	p_reg_fullgraph70: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph70 <= reg_fullgraph70_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph70 <= reg_fullgraph70_init;
        else
          reg_fullgraph70 <= reg_fullgraph70_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph70

		reg_q401 <= '1' when reg_fullgraph70 = "0001" else '0'; 
		reg_q695 <= '1' when reg_fullgraph70 = "0010" else '0'; 
		reg_q1397 <= '1' when reg_fullgraph70 = "0011" else '0'; 
		reg_q1676 <= '1' when reg_fullgraph70 = "0100" else '0'; 
		reg_q2154 <= '1' when reg_fullgraph70 = "0101" else '0'; 
		reg_q2550 <= '1' when reg_fullgraph70 = "0110" else '0'; 
		reg_q2505 <= '1' when reg_fullgraph70 = "0111" else '0'; 
		reg_q2655 <= '1' when reg_fullgraph70 = "1000" else '0'; 
		reg_q2503 <= '1' when reg_fullgraph70 = "1001" else '0'; 
		reg_q1652 <= '1' when reg_fullgraph70 = "1010" else '0'; 
--end decoder 
--######################################################
--fullgraph71

reg_q2495_in <= (reg_q2493 AND symb_decoder(16#73#)) OR
 					(reg_q2493 AND symb_decoder(16#53#));
reg_q946_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q945 AND symb_decoder(16#0a#)) OR
 					(reg_q945 AND symb_decoder(16#0d#));
reg_q648_in <= (reg_q646 AND symb_decoder(16#73#)) OR
 					(reg_q646 AND symb_decoder(16#53#));
reg_q310_in <= (reg_q308 AND symb_decoder(16#73#)) OR
 					(reg_q308 AND symb_decoder(16#53#));
reg_q1576_in <= (reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q1574 AND symb_decoder(16#57#)) OR
 					(reg_q1574 AND symb_decoder(16#77#));
reg_q1846_in <= (reg_q1844 AND symb_decoder(16#53#)) OR
 					(reg_q1844 AND symb_decoder(16#73#));
reg_q455_in <= (reg_q453 AND symb_decoder(16#73#)) OR
 					(reg_q453 AND symb_decoder(16#53#));
reg_q1447_in <= (reg_q1479 AND symb_decoder(16#46#)) OR
 					(reg_q1479 AND symb_decoder(16#66#)) OR
 					(reg_q1443 AND symb_decoder(16#46#)) OR
 					(reg_q1443 AND symb_decoder(16#66#));
reg_q1296_in <= (reg_q1294 AND symb_decoder(16#73#)) OR
 					(reg_q1294 AND symb_decoder(16#53#));
reg_q894_in <= (reg_q892 AND symb_decoder(16#73#)) OR
 					(reg_q892 AND symb_decoder(16#53#));
reg_q2487_in <= (reg_q2485 AND symb_decoder(16#73#)) OR
 					(reg_q2485 AND symb_decoder(16#53#));
reg_q1046_in <= (reg_q1044 AND symb_decoder(16#53#));
reg_q1596_in <= (reg_q1594 AND symb_decoder(16#53#)) OR
 					(reg_q1594 AND symb_decoder(16#73#));
reg_q1363_in <= (reg_q1361 AND symb_decoder(16#69#)) OR
 					(reg_q1361 AND symb_decoder(16#49#));
reg_fullgraph71_init <= "0000";

reg_fullgraph71_sel <= "00" & reg_q1363_in & reg_q1596_in & reg_q1046_in & reg_q2487_in & reg_q894_in & reg_q1296_in & reg_q1447_in & reg_q455_in & reg_q1846_in & reg_q1576_in & reg_q310_in & reg_q648_in & reg_q946_in & reg_q2495_in;

	--coder fullgraph71
with reg_fullgraph71_sel select
reg_fullgraph71_in <=
	"0001" when "0000000000000001",
	"0010" when "0000000000000010",
	"0011" when "0000000000000100",
	"0100" when "0000000000001000",
	"0101" when "0000000000010000",
	"0110" when "0000000000100000",
	"0111" when "0000000001000000",
	"1000" when "0000000010000000",
	"1001" when "0000000100000000",
	"1010" when "0000001000000000",
	"1011" when "0000010000000000",
	"1100" when "0000100000000000",
	"1101" when "0001000000000000",
	"1110" when "0010000000000000",
	"0000" when others;
 --end coder

	p_reg_fullgraph71: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph71 <= reg_fullgraph71_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph71 <= reg_fullgraph71_init;
        else
          reg_fullgraph71 <= reg_fullgraph71_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph71

		reg_q2495 <= '1' when reg_fullgraph71 = "0001" else '0'; 
		reg_q946 <= '1' when reg_fullgraph71 = "0010" else '0'; 
		reg_q648 <= '1' when reg_fullgraph71 = "0011" else '0'; 
		reg_q310 <= '1' when reg_fullgraph71 = "0100" else '0'; 
		reg_q1576 <= '1' when reg_fullgraph71 = "0101" else '0'; 
		reg_q1846 <= '1' when reg_fullgraph71 = "0110" else '0'; 
		reg_q455 <= '1' when reg_fullgraph71 = "0111" else '0'; 
		reg_q1447 <= '1' when reg_fullgraph71 = "1000" else '0'; 
		reg_q1296 <= '1' when reg_fullgraph71 = "1001" else '0'; 
		reg_q894 <= '1' when reg_fullgraph71 = "1010" else '0'; 
		reg_q2487 <= '1' when reg_fullgraph71 = "1011" else '0'; 
		reg_q1046 <= '1' when reg_fullgraph71 = "1100" else '0'; 
		reg_q1596 <= '1' when reg_fullgraph71 = "1101" else '0'; 
		reg_q1363 <= '1' when reg_fullgraph71 = "1110" else '0'; 
--end decoder 
--######################################################
--fullgraph72

reg_q1483_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q1482 AND symb_decoder(16#0d#)) OR
 					(reg_q1482 AND symb_decoder(16#0a#));
reg_q963_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q946 AND symb_decoder(16#53#));
reg_q1220_in <= (reg_q2757 AND symb_decoder(16#57#)) OR
 					(reg_q2757 AND symb_decoder(16#77#)) OR
 					(reg_q1218 AND symb_decoder(16#57#)) OR
 					(reg_q1218 AND symb_decoder(16#77#));
reg_fullgraph72_init <= "00";

reg_fullgraph72_sel <= "0" & reg_q1220_in & reg_q963_in & reg_q1483_in;

	--coder fullgraph72
with reg_fullgraph72_sel select
reg_fullgraph72_in <=
	"01" when "0001",
	"10" when "0010",
	"11" when "0100",
	"00" when others;
 --end coder

	p_reg_fullgraph72: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph72 <= reg_fullgraph72_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph72 <= reg_fullgraph72_init;
        else
          reg_fullgraph72 <= reg_fullgraph72_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph72

		reg_q1483 <= '1' when reg_fullgraph72 = "01" else '0'; 
		reg_q963 <= '1' when reg_fullgraph72 = "10" else '0'; 
		reg_q1220 <= '1' when reg_fullgraph72 = "11" else '0'; 
--end decoder 
--######################################################
--fullgraph73

reg_q861_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q860 AND symb_decoder(16#0d#)) OR
 					(reg_q860 AND symb_decoder(16#0a#));
reg_q547_in <= (reg_q2757 AND symb_decoder(16#53#)) OR
 					(reg_q2757 AND symb_decoder(16#73#)) OR
 					(reg_q546 AND symb_decoder(16#73#)) OR
 					(reg_q546 AND symb_decoder(16#53#));
reg_fullgraph73_init <= "00";

reg_fullgraph73_sel <= "00" & reg_q547_in & reg_q861_in;

	--coder fullgraph73
with reg_fullgraph73_sel select
reg_fullgraph73_in <=
	"01" when "0001",
	"10" when "0010",
	"00" when others;
 --end coder

	p_reg_fullgraph73: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph73 <= reg_fullgraph73_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph73 <= reg_fullgraph73_init;
        else
          reg_fullgraph73 <= reg_fullgraph73_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph73

		reg_q861 <= '1' when reg_fullgraph73 = "01" else '0'; 
		reg_q547 <= '1' when reg_fullgraph73 = "10" else '0'; 
--end decoder 

reg_q134_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q133 AND symb_decoder(16#0d#)) OR
 					(reg_q133 AND symb_decoder(16#0a#));
reg_q134_init <= '0' ;
	p_reg_q134: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q134 <= reg_q134_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q134 <= reg_q134_init;
        else
          reg_q134 <= reg_q134_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2330_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2329 AND symb_decoder(16#0a#)) OR
 					(reg_q2329 AND symb_decoder(16#0d#));
reg_q2330_init <= '0' ;
	p_reg_q2330: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2330 <= reg_q2330_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2330 <= reg_q2330_init;
        else
          reg_q2330 <= reg_q2330_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q346_in <= (reg_q345 AND symb_decoder(16#0d#)) OR
 					(reg_q345 AND symb_decoder(16#0a#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#));
reg_q346_init <= '0' ;
	p_reg_q346: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q346 <= reg_q346_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q346 <= reg_q346_init;
        else
          reg_q346 <= reg_q346_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph77

reg_q2294_in <= (reg_q2290 AND symb_decoder(16#0d#)) OR
 					(reg_q2326 AND symb_decoder(16#0d#));
reg_q2296_in <= (reg_q2294 AND symb_decoder(16#0a#));
reg_fullgraph77_init <= "00";

reg_fullgraph77_sel <= "00" & reg_q2296_in & reg_q2294_in;

	--coder fullgraph77
with reg_fullgraph77_sel select
reg_fullgraph77_in <=
	"01" when "0001",
	"10" when "0010",
	"00" when others;
 --end coder

	p_reg_fullgraph77: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph77 <= reg_fullgraph77_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph77 <= reg_fullgraph77_init;
        else
          reg_fullgraph77 <= reg_fullgraph77_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph77

		reg_q2294 <= '1' when reg_fullgraph77 = "01" else '0'; 
		reg_q2296 <= '1' when reg_fullgraph77 = "10" else '0'; 
--end decoder 

reg_q2521_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2520 AND symb_decoder(16#0a#)) OR
 					(reg_q2520 AND symb_decoder(16#0d#));
reg_q2521_init <= '0' ;
	p_reg_q2521: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2521 <= reg_q2521_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2521 <= reg_q2521_init;
        else
          reg_q2521 <= reg_q2521_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q662_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q661 AND symb_decoder(16#0d#)) OR
 					(reg_q661 AND symb_decoder(16#0a#));
reg_q662_init <= '0' ;
	p_reg_q662: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q662 <= reg_q662_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q662 <= reg_q662_init;
        else
          reg_q662 <= reg_q662_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q758_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q757 AND symb_decoder(16#0a#)) OR
 					(reg_q757 AND symb_decoder(16#0d#));
reg_q758_init <= '0' ;
	p_reg_q758: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q758 <= reg_q758_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q758 <= reg_q758_init;
        else
          reg_q758 <= reg_q758_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q189_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q188 AND symb_decoder(16#0a#)) OR
 					(reg_q188 AND symb_decoder(16#0d#));
reg_q189_init <= '0' ;
	p_reg_q189: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q189 <= reg_q189_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q189 <= reg_q189_init;
        else
          reg_q189 <= reg_q189_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2245_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2244 AND symb_decoder(16#0a#)) OR
 					(reg_q2244 AND symb_decoder(16#0d#));
reg_q2245_init <= '0' ;
	p_reg_q2245: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2245 <= reg_q2245_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2245 <= reg_q2245_init;
        else
          reg_q2245 <= reg_q2245_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1097_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q1096 AND symb_decoder(16#0a#)) OR
 					(reg_q1096 AND symb_decoder(16#0d#));
reg_q1097_init <= '0' ;
	p_reg_q1097: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1097 <= reg_q1097_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1097 <= reg_q1097_init;
        else
          reg_q1097 <= reg_q1097_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q100_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q99 AND symb_decoder(16#0d#)) OR
 					(reg_q99 AND symb_decoder(16#0a#));
reg_q100_init <= '0' ;
	p_reg_q100: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q100 <= reg_q100_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q100 <= reg_q100_init;
        else
          reg_q100 <= reg_q100_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q804_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q803 AND symb_decoder(16#0a#)) OR
 					(reg_q803 AND symb_decoder(16#0d#));
reg_q804_init <= '0' ;
	p_reg_q804: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q804 <= reg_q804_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q804 <= reg_q804_init;
        else
          reg_q804 <= reg_q804_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q591_in <= (reg_q590 AND symb_decoder(16#0a#)) OR
 					(reg_q590 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#));
reg_q591_init <= '0' ;
	p_reg_q591: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q591 <= reg_q591_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q591 <= reg_q591_init;
        else
          reg_q591 <= reg_q591_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1310_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q1309 AND symb_decoder(16#0d#)) OR
 					(reg_q1309 AND symb_decoder(16#0a#));
reg_q1310_init <= '0' ;
	p_reg_q1310: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1310 <= reg_q1310_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1310 <= reg_q1310_init;
        else
          reg_q1310 <= reg_q1310_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1205_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q1204 AND symb_decoder(16#0a#)) OR
 					(reg_q1204 AND symb_decoder(16#0d#));
reg_q1205_init <= '0' ;
	p_reg_q1205: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1205 <= reg_q1205_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1205 <= reg_q1205_init;
        else
          reg_q1205 <= reg_q1205_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q517_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q516 AND symb_decoder(16#0a#)) OR
 					(reg_q516 AND symb_decoder(16#0d#));
reg_q517_init <= '0' ;
	p_reg_q517: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q517 <= reg_q517_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q517 <= reg_q517_init;
        else
          reg_q517 <= reg_q517_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q1 AND symb_decoder(16#0d#)) OR
 					(reg_q1 AND symb_decoder(16#0a#));
reg_q2_init <= '0' ;
	p_reg_q2: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2 <= reg_q2_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2 <= reg_q2_init;
        else
          reg_q2 <= reg_q2_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2222_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q2221 AND symb_decoder(16#0d#)) OR
 					(reg_q2221 AND symb_decoder(16#0a#));
reg_q2222_init <= '0' ;
	p_reg_q2222: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2222 <= reg_q2222_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2222 <= reg_q2222_init;
        else
          reg_q2222 <= reg_q2222_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1062_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q1061 AND symb_decoder(16#0d#)) OR
 					(reg_q1061 AND symb_decoder(16#0a#));
reg_q1062_init <= '0' ;
	p_reg_q1062: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1062 <= reg_q1062_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1062 <= reg_q1062_init;
        else
          reg_q1062 <= reg_q1062_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q971_in <= (reg_q2757 AND symb_decoder(16#0d#)) OR
 					(reg_q2757 AND symb_decoder(16#0a#)) OR
 					(reg_q970 AND symb_decoder(16#0d#)) OR
 					(reg_q970 AND symb_decoder(16#0a#));
reg_q971_init <= '0' ;
	p_reg_q971: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q971 <= reg_q971_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q971 <= reg_q971_init;
        else
          reg_q971 <= reg_q971_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q111_in <= (reg_q107 AND symb_decoder(16#0a#)) OR
 					(reg_q113 AND symb_decoder(16#0a#));
reg_q111_init <= '0' ;
	p_reg_q111: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q111 <= reg_q111_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q111 <= reg_q111_init;
        else
          reg_q111 <= reg_q111_in;
        end if;
      end if;
    end if;
  end process;

	
FINAL <= reg_q585 OR reg_q2550 OR reg_q691 OR reg_q513 OR reg_q658 OR reg_q1201 OR reg_q754 OR reg_q1915 OR reg_q767 OR reg_q1814 OR reg_q342 OR reg_q2445 OR reg_q2241 OR reg_q1058 OR reg_q602 OR reg_q960 OR reg_q1520 OR reg_q1216 OR reg_q1949 OR reg_q2675 OR reg_q855 OR reg_q1020 OR reg_q97 OR reg_q1973 OR reg_q2397 OR reg_q768 OR reg_q2214 OR reg_q1680 OR reg_q1306 OR reg_q2054 OR reg_q2631 OR reg_q2755 OR reg_q2227 OR reg_q940 OR reg_q492 OR reg_q1572 OR reg_q1753 OR reg_q2324 OR reg_q1477 OR reg_q1624 OR reg_q467 OR reg_q2754 OR reg_q538 OR reg_q60 OR reg_q2517 OR reg_q391 OR reg_q2050 OR reg_q183 OR reg_q111 OR reg_q959 OR reg_q1932 OR reg_q130 OR reg_q1898 OR reg_q1391 OR reg_q1093 OR reg_q284 OR reg_q798 OR reg_q2580 OR reg_q1142;

	end architecture;
	