-- pattern_match.vhd: a simple pattern matching unit with some optimizations

library ieee;
use ieee.std_logic_1164.all;


architecture backdoor_subset_4 of pattern_match is

  -- state q889
  signal reg_q889        : std_logic;
  signal reg_q889_in     : std_logic;
  signal reg_q889_init   : std_logic;
		

  -- state q896
  signal reg_q896        : std_logic;
  signal reg_q896_in     : std_logic;
  signal reg_q896_init   : std_logic;
		

  -- state q178
  signal reg_q178        : std_logic;
  signal reg_q178_in     : std_logic;
  signal reg_q178_init   : std_logic;
		

  -- state q1812
  signal reg_q1812        : std_logic;
  signal reg_q1812_in     : std_logic;
  signal reg_q1812_init   : std_logic;
		

  -- state q1814
  signal reg_q1814        : std_logic;
  signal reg_q1814_in     : std_logic;
  signal reg_q1814_init   : std_logic;
		

  -- state q1013
  signal reg_q1013        : std_logic;
  signal reg_q1013_in     : std_logic;
  signal reg_q1013_init   : std_logic;
		

  -- state q2695
  signal reg_q2695        : std_logic;
  signal reg_q2695_in     : std_logic;
  signal reg_q2695_init   : std_logic;
		

  -- state q779
  signal reg_q779        : std_logic;
  signal reg_q779_in     : std_logic;
  signal reg_q779_init   : std_logic;
		

  -- state q2124
  signal reg_q2124        : std_logic;
  signal reg_q2124_in     : std_logic;
  signal reg_q2124_init   : std_logic;
		

  -- state q665
  signal reg_q665        : std_logic;
  signal reg_q665_in     : std_logic;
  signal reg_q665_init   : std_logic;
		

  -- state q816
  signal reg_q816        : std_logic;
  signal reg_q816_in     : std_logic;
  signal reg_q816_init   : std_logic;
		

  -- state q1297
  signal reg_q1297        : std_logic;
  signal reg_q1297_in     : std_logic;
  signal reg_q1297_init   : std_logic;
		

  -- state q2618
  signal reg_q2618        : std_logic;
  signal reg_q2618_in     : std_logic;
  signal reg_q2618_init   : std_logic;
		

  -- state q850
  signal reg_q850        : std_logic;
  signal reg_q850_in     : std_logic;
  signal reg_q850_init   : std_logic;
		

  -- state q1224
  signal reg_q1224        : std_logic;
  signal reg_q1224_in     : std_logic;
  signal reg_q1224_init   : std_logic;
		

  -- state q813
  signal reg_q813        : std_logic;
  signal reg_q813_in     : std_logic;
  signal reg_q813_init   : std_logic;
		

  -- state q2000
  signal reg_q2000        : std_logic;
  signal reg_q2000_in     : std_logic;
  signal reg_q2000_init   : std_logic;
		

  -- state q225
  signal reg_q225        : std_logic;
  signal reg_q225_in     : std_logic;
  signal reg_q225_init   : std_logic;
		

  -- state q899
  signal reg_q899        : std_logic;
  signal reg_q899_in     : std_logic;
  signal reg_q899_init   : std_logic;
		

  -- state q1826
  signal reg_q1826        : std_logic;
  signal reg_q1826_in     : std_logic;
  signal reg_q1826_init   : std_logic;
		

  -- state q1452
  signal reg_q1452        : std_logic;
  signal reg_q1452_in     : std_logic;
  signal reg_q1452_init   : std_logic;
		

  -- state q958
  signal reg_q958        : std_logic;
  signal reg_q958_in     : std_logic;
  signal reg_q958_init   : std_logic;
		

  -- state q2211
  signal reg_q2211        : std_logic;
  signal reg_q2211_in     : std_logic;
  signal reg_q2211_init   : std_logic;
		

  -- state q0
  signal reg_q0        : std_logic;
  signal reg_q0_in     : std_logic;
  signal reg_q0_init   : std_logic;
		

  -- state q303
  signal reg_q303        : std_logic;
  signal reg_q303_in     : std_logic;
  signal reg_q303_init   : std_logic;
		

  -- state q247
  signal reg_q247        : std_logic;
  signal reg_q247_in     : std_logic;
  signal reg_q247_init   : std_logic;
		

  -- state q249
  signal reg_q249        : std_logic;
  signal reg_q249_in     : std_logic;
  signal reg_q249_init   : std_logic;
		

  -- state q2615
  signal reg_q2615        : std_logic;
  signal reg_q2615_in     : std_logic;
  signal reg_q2615_init   : std_logic;
		

  -- state q2518
  signal reg_q2518        : std_logic;
  signal reg_q2518_in     : std_logic;
  signal reg_q2518_init   : std_logic;
		

  -- state q791
  signal reg_q791        : std_logic;
  signal reg_q791_in     : std_logic;
  signal reg_q791_init   : std_logic;
		

  -- state q828
  signal reg_q828        : std_logic;
  signal reg_q828_in     : std_logic;
  signal reg_q828_init   : std_logic;
		

  -- state q848
  signal reg_q848        : std_logic;
  signal reg_q848_in     : std_logic;
  signal reg_q848_init   : std_logic;
		

  -- state q119
  signal reg_q119        : std_logic;
  signal reg_q119_in     : std_logic;
  signal reg_q119_init   : std_logic;
		

  -- state q121
  signal reg_q121        : std_logic;
  signal reg_q121_in     : std_logic;
  signal reg_q121_init   : std_logic;
		

  -- state q1207
  signal reg_q1207        : std_logic;
  signal reg_q1207_in     : std_logic;
  signal reg_q1207_init   : std_logic;
		

  -- state q1209
  signal reg_q1209        : std_logic;
  signal reg_q1209_in     : std_logic;
  signal reg_q1209_init   : std_logic;
		

  -- state q74
  signal reg_q74        : std_logic;
  signal reg_q74_in     : std_logic;
  signal reg_q74_init   : std_logic;
		

  -- state q76
  signal reg_q76        : std_logic;
  signal reg_q76_in     : std_logic;
  signal reg_q76_init   : std_logic;
		

  -- state q1189
  signal reg_q1189        : std_logic;
  signal reg_q1189_in     : std_logic;
  signal reg_q1189_init   : std_logic;
		

  -- state q1191
  signal reg_q1191        : std_logic;
  signal reg_q1191_in     : std_logic;
  signal reg_q1191_init   : std_logic;
		

  -- state q262
  signal reg_q262        : std_logic;
  signal reg_q262_in     : std_logic;
  signal reg_q262_init   : std_logic;
		

  -- state q1884
  signal reg_q1884        : std_logic;
  signal reg_q1884_in     : std_logic;
  signal reg_q1884_init   : std_logic;
		

  -- state q2383
  signal reg_q2383        : std_logic;
  signal reg_q2383_in     : std_logic;
  signal reg_q2383_init   : std_logic;
		

  -- state q414
  signal reg_q414        : std_logic;
  signal reg_q414_in     : std_logic;
  signal reg_q414_init   : std_logic;
		

  -- state q2252
  signal reg_q2252        : std_logic;
  signal reg_q2252_in     : std_logic;
  signal reg_q2252_init   : std_logic;
		

  -- state q913
  signal reg_q913        : std_logic;
  signal reg_q913_in     : std_logic;
  signal reg_q913_init   : std_logic;
		

  -- state q915
  signal reg_q915        : std_logic;
  signal reg_q915_in     : std_logic;
  signal reg_q915_init   : std_logic;
		

  -- state q2192
  signal reg_q2192        : std_logic;
  signal reg_q2192_in     : std_logic;
  signal reg_q2192_init   : std_logic;
		

  -- state q2194
  signal reg_q2194        : std_logic;
  signal reg_q2194_in     : std_logic;
  signal reg_q2194_init   : std_logic;
		

  -- state q680
  signal reg_q680        : std_logic;
  signal reg_q680_in     : std_logic;
  signal reg_q680_init   : std_logic;
		

  -- state q452
  signal reg_q452        : std_logic;
  signal reg_q452_in     : std_logic;
  signal reg_q452_init   : std_logic;
		

  -- state q556
  signal reg_q556        : std_logic;
  signal reg_q556_in     : std_logic;
  signal reg_q556_init   : std_logic;
		

  -- state q1111
  signal reg_q1111        : std_logic;
  signal reg_q1111_in     : std_logic;
  signal reg_q1111_init   : std_logic;
		

  -- state q1644
  signal reg_q1644        : std_logic;
  signal reg_q1644_in     : std_logic;
  signal reg_q1644_init   : std_logic;
		

  -- state q2249
  signal reg_q2249        : std_logic;
  signal reg_q2249_in     : std_logic;
  signal reg_q2249_init   : std_logic;
		

  -- state q799
  signal reg_q799        : std_logic;
  signal reg_q799_in     : std_logic;
  signal reg_q799_init   : std_logic;
		

  -- state q801
  signal reg_q801        : std_logic;
  signal reg_q801_in     : std_logic;
  signal reg_q801_init   : std_logic;
		

  -- state q1195
  signal reg_q1195        : std_logic;
  signal reg_q1195_in     : std_logic;
  signal reg_q1195_init   : std_logic;
		

  -- state q2373
  signal reg_q2373        : std_logic;
  signal reg_q2373_in     : std_logic;
  signal reg_q2373_init   : std_logic;
		

  -- state q91
  signal reg_q91        : std_logic;
  signal reg_q91_in     : std_logic;
  signal reg_q91_init   : std_logic;
		

  -- state q125
  signal reg_q125        : std_logic;
  signal reg_q125_in     : std_logic;
  signal reg_q125_init   : std_logic;
		

  -- state q127
  signal reg_q127        : std_logic;
  signal reg_q127_in     : std_logic;
  signal reg_q127_init   : std_logic;
		

  -- state q714
  signal reg_q714        : std_logic;
  signal reg_q714_in     : std_logic;
  signal reg_q714_init   : std_logic;
		

  -- state q1544
  signal reg_q1544        : std_logic;
  signal reg_q1544_in     : std_logic;
  signal reg_q1544_init   : std_logic;
		

  -- state q1928
  signal reg_q1928        : std_logic;
  signal reg_q1928_in     : std_logic;
  signal reg_q1928_init   : std_logic;
		

  -- state q1930
  signal reg_q1930        : std_logic;
  signal reg_q1930_in     : std_logic;
  signal reg_q1930_init   : std_logic;
		

  -- state q2533
  signal reg_q2533        : std_logic;
  signal reg_q2533_in     : std_logic;
  signal reg_q2533_init   : std_logic;
		

  -- state q1742
  signal reg_q1742        : std_logic;
  signal reg_q1742_in     : std_logic;
  signal reg_q1742_init   : std_logic;
		

  -- state q1668
  signal reg_q1668        : std_logic;
  signal reg_q1668_in     : std_logic;
  signal reg_q1668_init   : std_logic;
		

  -- state q1670
  signal reg_q1670        : std_logic;
  signal reg_q1670_in     : std_logic;
  signal reg_q1670_init   : std_logic;
		

  -- state q1050
  signal reg_q1050        : std_logic;
  signal reg_q1050_in     : std_logic;
  signal reg_q1050_init   : std_logic;
		

  -- state q780
  signal reg_q780        : std_logic;
  signal reg_q780_in     : std_logic;
  signal reg_q780_init   : std_logic;
		

  -- state q2156
  signal reg_q2156        : std_logic;
  signal reg_q2156_in     : std_logic;
  signal reg_q2156_init   : std_logic;
		

  -- state q2158
  signal reg_q2158        : std_logic;
  signal reg_q2158_in     : std_logic;
  signal reg_q2158_init   : std_logic;
		

  -- state q1521
  signal reg_q1521        : std_logic;
  signal reg_q1521_in     : std_logic;
  signal reg_q1521_init   : std_logic;
		

  -- state q1377
  signal reg_q1377        : std_logic;
  signal reg_q1377_in     : std_logic;
  signal reg_q1377_init   : std_logic;
		

  -- state q1379
  signal reg_q1379        : std_logic;
  signal reg_q1379_in     : std_logic;
  signal reg_q1379_init   : std_logic;
		

  -- state q688
  signal reg_q688        : std_logic;
  signal reg_q688_in     : std_logic;
  signal reg_q688_init   : std_logic;
		

  -- state q690
  signal reg_q690        : std_logic;
  signal reg_q690_in     : std_logic;
  signal reg_q690_init   : std_logic;
		

  -- state q644
  signal reg_q644        : std_logic;
  signal reg_q644_in     : std_logic;
  signal reg_q644_init   : std_logic;
		

  -- state q646
  signal reg_q646        : std_logic;
  signal reg_q646_in     : std_logic;
  signal reg_q646_init   : std_logic;
		

  -- state q1955
  signal reg_q1955        : std_logic;
  signal reg_q1955_in     : std_logic;
  signal reg_q1955_init   : std_logic;
		

  -- state q1848
  signal reg_q1848        : std_logic;
  signal reg_q1848_in     : std_logic;
  signal reg_q1848_init   : std_logic;
		

  -- state q52
  signal reg_q52        : std_logic;
  signal reg_q52_in     : std_logic;
  signal reg_q52_init   : std_logic;
		

  -- state q54
  signal reg_q54        : std_logic;
  signal reg_q54_in     : std_logic;
  signal reg_q54_init   : std_logic;
		

  -- state q630
  signal reg_q630        : std_logic;
  signal reg_q630_in     : std_logic;
  signal reg_q630_init   : std_logic;
		

  -- state q632
  signal reg_q632        : std_logic;
  signal reg_q632_in     : std_logic;
  signal reg_q632_init   : std_logic;
		

  -- state q703
  signal reg_q703        : std_logic;
  signal reg_q703_in     : std_logic;
  signal reg_q703_init   : std_logic;
		

  -- state q1574
  signal reg_q1574        : std_logic;
  signal reg_q1574_in     : std_logic;
  signal reg_q1574_init   : std_logic;
		

  -- state q1576
  signal reg_q1576        : std_logic;
  signal reg_q1576_in     : std_logic;
  signal reg_q1576_init   : std_logic;
		

  -- state q2172
  signal reg_q2172        : std_logic;
  signal reg_q2172_in     : std_logic;
  signal reg_q2172_init   : std_logic;
		

  -- state q2208
  signal reg_q2208        : std_logic;
  signal reg_q2208_in     : std_logic;
  signal reg_q2208_init   : std_logic;
		

  -- state q1997
  signal reg_q1997        : std_logic;
  signal reg_q1997_in     : std_logic;
  signal reg_q1997_init   : std_logic;
		

  -- state q933
  signal reg_q933        : std_logic;
  signal reg_q933_in     : std_logic;
  signal reg_q933_init   : std_logic;
		

  -- state q955
  signal reg_q955        : std_logic;
  signal reg_q955_in     : std_logic;
  signal reg_q955_init   : std_logic;
		

  -- state q2091
  signal reg_q2091        : std_logic;
  signal reg_q2091_in     : std_logic;
  signal reg_q2091_init   : std_logic;
		

  -- state q2636
  signal reg_q2636        : std_logic;
  signal reg_q2636_in     : std_logic;
  signal reg_q2636_init   : std_logic;
		

  -- state q2638
  signal reg_q2638        : std_logic;
  signal reg_q2638_in     : std_logic;
  signal reg_q2638_init   : std_logic;
		

  -- state q606
  signal reg_q606        : std_logic;
  signal reg_q606_in     : std_logic;
  signal reg_q606_init   : std_logic;
		

  -- state q608
  signal reg_q608        : std_logic;
  signal reg_q608_in     : std_logic;
  signal reg_q608_init   : std_logic;
		

  -- state q1355
  signal reg_q1355        : std_logic;
  signal reg_q1355_in     : std_logic;
  signal reg_q1355_init   : std_logic;
		

  -- state q618
  signal reg_q618        : std_logic;
  signal reg_q618_in     : std_logic;
  signal reg_q618_init   : std_logic;
		

  -- state q1359
  signal reg_q1359        : std_logic;
  signal reg_q1359_in     : std_logic;
  signal reg_q1359_init   : std_logic;
		

  -- state q2052
  signal reg_q2052        : std_logic;
  signal reg_q2052_in     : std_logic;
  signal reg_q2052_init   : std_logic;
		

  -- state q363
  signal reg_q363        : std_logic;
  signal reg_q363_in     : std_logic;
  signal reg_q363_init   : std_logic;
		

  -- state q365
  signal reg_q365        : std_logic;
  signal reg_q365_in     : std_logic;
  signal reg_q365_init   : std_logic;
		

  -- state q1137
  signal reg_q1137        : std_logic;
  signal reg_q1137_in     : std_logic;
  signal reg_q1137_init   : std_logic;
		

  -- state q1139
  signal reg_q1139        : std_logic;
  signal reg_q1139_in     : std_logic;
  signal reg_q1139_init   : std_logic;
		

  -- state q696
  signal reg_q696        : std_logic;
  signal reg_q696_in     : std_logic;
  signal reg_q696_init   : std_logic;
		

  -- state q698
  signal reg_q698        : std_logic;
  signal reg_q698_in     : std_logic;
  signal reg_q698_init   : std_logic;
		

  -- state q472
  signal reg_q472        : std_logic;
  signal reg_q472_in     : std_logic;
  signal reg_q472_init   : std_logic;
		

  -- state q474
  signal reg_q474        : std_logic;
  signal reg_q474_in     : std_logic;
  signal reg_q474_init   : std_logic;
		

  -- state q1816
  signal reg_q1816        : std_logic;
  signal reg_q1816_in     : std_logic;
  signal reg_q1816_init   : std_logic;
		

  -- state q1818
  signal reg_q1818        : std_logic;
  signal reg_q1818_in     : std_logic;
  signal reg_q1818_init   : std_logic;
		

  -- state q1975
  signal reg_q1975        : std_logic;
  signal reg_q1975_in     : std_logic;
  signal reg_q1975_init   : std_logic;
		

  -- state q46
  signal reg_q46        : std_logic;
  signal reg_q46_in     : std_logic;
  signal reg_q46_init   : std_logic;
		

  -- state q2461
  signal reg_q2461        : std_logic;
  signal reg_q2461_in     : std_logic;
  signal reg_q2461_init   : std_logic;
		

  -- state q2463
  signal reg_q2463        : std_logic;
  signal reg_q2463_in     : std_logic;
  signal reg_q2463_init   : std_logic;
		

  -- state q700
  signal reg_q700        : std_logic;
  signal reg_q700_in     : std_logic;
  signal reg_q700_init   : std_logic;
		

  -- state q58
  signal reg_q58        : std_logic;
  signal reg_q58_in     : std_logic;
  signal reg_q58_init   : std_logic;
		

  -- state q2030
  signal reg_q2030        : std_logic;
  signal reg_q2030_in     : std_logic;
  signal reg_q2030_init   : std_logic;
		

  -- state q2032
  signal reg_q2032        : std_logic;
  signal reg_q2032_in     : std_logic;
  signal reg_q2032_init   : std_logic;
		

  -- state q1926
  signal reg_q1926        : std_logic;
  signal reg_q1926_in     : std_logic;
  signal reg_q1926_init   : std_logic;
		

  -- state q1246
  signal reg_q1246        : std_logic;
  signal reg_q1246_in     : std_logic;
  signal reg_q1246_init   : std_logic;
		

  -- state q1248
  signal reg_q1248        : std_logic;
  signal reg_q1248_in     : std_logic;
  signal reg_q1248_init   : std_logic;
		

  -- state q616
  signal reg_q616        : std_logic;
  signal reg_q616_in     : std_logic;
  signal reg_q616_init   : std_logic;
		

  -- state q2411
  signal reg_q2411        : std_logic;
  signal reg_q2411_in     : std_logic;
  signal reg_q2411_init   : std_logic;
		

  -- state q1770
  signal reg_q1770        : std_logic;
  signal reg_q1770_in     : std_logic;
  signal reg_q1770_init   : std_logic;
		

  -- state q1772
  signal reg_q1772        : std_logic;
  signal reg_q1772_in     : std_logic;
  signal reg_q1772_init   : std_logic;
		

  -- state q520
  signal reg_q520        : std_logic;
  signal reg_q520_in     : std_logic;
  signal reg_q520_init   : std_logic;
		

  -- state q522
  signal reg_q522        : std_logic;
  signal reg_q522_in     : std_logic;
  signal reg_q522_init   : std_logic;
		

  -- state q2103
  signal reg_q2103        : std_logic;
  signal reg_q2103_in     : std_logic;
  signal reg_q2103_init   : std_logic;
		

  -- state q2105
  signal reg_q2105        : std_logic;
  signal reg_q2105_in     : std_logic;
  signal reg_q2105_init   : std_logic;
		

  -- state q2300
  signal reg_q2300        : std_logic;
  signal reg_q2300_in     : std_logic;
  signal reg_q2300_init   : std_logic;
		

  -- state q2302
  signal reg_q2302        : std_logic;
  signal reg_q2302_in     : std_logic;
  signal reg_q2302_init   : std_logic;
		

  -- state q2130
  signal reg_q2130        : std_logic;
  signal reg_q2130_in     : std_logic;
  signal reg_q2130_init   : std_logic;
		

  -- state q22
  signal reg_q22        : std_logic;
  signal reg_q22_in     : std_logic;
  signal reg_q22_init   : std_logic;
		

  -- state q2579
  signal reg_q2579        : std_logic;
  signal reg_q2579_in     : std_logic;
  signal reg_q2579_init   : std_logic;
		

  -- state q671
  signal reg_q671        : std_logic;
  signal reg_q671_in     : std_logic;
  signal reg_q671_init   : std_logic;
		

  -- state q673
  signal reg_q673        : std_logic;
  signal reg_q673_in     : std_logic;
  signal reg_q673_init   : std_logic;
		

  -- state q2
  signal reg_q2        : std_logic;
  signal reg_q2_in     : std_logic;
  signal reg_q2_init   : std_logic;
		

  -- state q2323
  signal reg_q2323        : std_logic;
  signal reg_q2323_in     : std_logic;
  signal reg_q2323_init   : std_logic;
		

  -- state q2128
  signal reg_q2128        : std_logic;
  signal reg_q2128_in     : std_logic;
  signal reg_q2128_init   : std_logic;
		

  -- state q2254
  signal reg_q2254        : std_logic;
  signal reg_q2254_in     : std_logic;
  signal reg_q2254_init   : std_logic;
		

  -- state q2256
  signal reg_q2256        : std_logic;
  signal reg_q2256_in     : std_logic;
  signal reg_q2256_init   : std_logic;
		

  -- state q351
  signal reg_q351        : std_logic;
  signal reg_q351_in     : std_logic;
  signal reg_q351_init   : std_logic;
		

  -- state q353
  signal reg_q353        : std_logic;
  signal reg_q353_in     : std_logic;
  signal reg_q353_init   : std_logic;
		

  -- state q2601
  signal reg_q2601        : std_logic;
  signal reg_q2601_in     : std_logic;
  signal reg_q2601_init   : std_logic;
		

  -- state q1393
  signal reg_q1393        : std_logic;
  signal reg_q1393_in     : std_logic;
  signal reg_q1393_init   : std_logic;
		

  -- state q1395
  signal reg_q1395        : std_logic;
  signal reg_q1395_in     : std_logic;
  signal reg_q1395_init   : std_logic;
		

  -- state q876
  signal reg_q876        : std_logic;
  signal reg_q876_in     : std_logic;
  signal reg_q876_init   : std_logic;
		

  -- state q878
  signal reg_q878        : std_logic;
  signal reg_q878_in     : std_logic;
  signal reg_q878_init   : std_logic;
		

  -- state q1535
  signal reg_q1535        : std_logic;
  signal reg_q1535_in     : std_logic;
  signal reg_q1535_init   : std_logic;
		

  -- state q1537
  signal reg_q1537        : std_logic;
  signal reg_q1537_in     : std_logic;
  signal reg_q1537_init   : std_logic;
		

  -- state q844
  signal reg_q844        : std_logic;
  signal reg_q844_in     : std_logic;
  signal reg_q844_init   : std_logic;
		

  -- state q257
  signal reg_q257        : std_logic;
  signal reg_q257_in     : std_logic;
  signal reg_q257_init   : std_logic;
		

  -- state q1313
  signal reg_q1313        : std_logic;
  signal reg_q1313_in     : std_logic;
  signal reg_q1313_init   : std_logic;
		

  -- state q1315
  signal reg_q1315        : std_logic;
  signal reg_q1315_in     : std_logic;
  signal reg_q1315_init   : std_logic;
		

  -- state q880
  signal reg_q880        : std_logic;
  signal reg_q880_in     : std_logic;
  signal reg_q880_init   : std_logic;
		

  -- state q882
  signal reg_q882        : std_logic;
  signal reg_q882_in     : std_logic;
  signal reg_q882_init   : std_logic;
		

  -- state q807
  signal reg_q807        : std_logic;
  signal reg_q807_in     : std_logic;
  signal reg_q807_init   : std_logic;
		

  -- state q809
  signal reg_q809        : std_logic;
  signal reg_q809_in     : std_logic;
  signal reg_q809_init   : std_logic;
		

  -- state q379
  signal reg_q379        : std_logic;
  signal reg_q379_in     : std_logic;
  signal reg_q379_init   : std_logic;
		

  -- state q381
  signal reg_q381        : std_logic;
  signal reg_q381_in     : std_logic;
  signal reg_q381_init   : std_logic;
		

  -- state q832
  signal reg_q832        : std_logic;
  signal reg_q832_in     : std_logic;
  signal reg_q832_init   : std_logic;
		

  -- state q945
  signal reg_q945        : std_logic;
  signal reg_q945_in     : std_logic;
  signal reg_q945_init   : std_logic;
		

  -- state q947
  signal reg_q947        : std_logic;
  signal reg_q947_in     : std_logic;
  signal reg_q947_init   : std_logic;
		

  -- state q2395
  signal reg_q2395        : std_logic;
  signal reg_q2395_in     : std_logic;
  signal reg_q2395_init   : std_logic;
		

  -- state q2397
  signal reg_q2397        : std_logic;
  signal reg_q2397_in     : std_logic;
  signal reg_q2397_init   : std_logic;
		

  -- state q1345
  signal reg_q1345        : std_logic;
  signal reg_q1345_in     : std_logic;
  signal reg_q1345_init   : std_logic;
		

  -- state q566
  signal reg_q566        : std_logic;
  signal reg_q566_in     : std_logic;
  signal reg_q566_init   : std_logic;
		

  -- state q568
  signal reg_q568        : std_logic;
  signal reg_q568_in     : std_logic;
  signal reg_q568_init   : std_logic;
		

  -- state q2514
  signal reg_q2514        : std_logic;
  signal reg_q2514_in     : std_logic;
  signal reg_q2514_init   : std_logic;
		

  -- state q2516
  signal reg_q2516        : std_logic;
  signal reg_q2516_in     : std_logic;
  signal reg_q2516_init   : std_logic;
		

  -- state q2530
  signal reg_q2530        : std_logic;
  signal reg_q2530_in     : std_logic;
  signal reg_q2530_init   : std_logic;
		

  -- state q56
  signal reg_q56        : std_logic;
  signal reg_q56_in     : std_logic;
  signal reg_q56_init   : std_logic;
		

  -- state q530
  signal reg_q530        : std_logic;
  signal reg_q530_in     : std_logic;
  signal reg_q530_init   : std_logic;
		

  -- state q1603
  signal reg_q1603        : std_logic;
  signal reg_q1603_in     : std_logic;
  signal reg_q1603_init   : std_logic;
		

  -- state q907
  signal reg_q907        : std_logic;
  signal reg_q907_in     : std_logic;
  signal reg_q907_init   : std_logic;
		

  -- state q909
  signal reg_q909        : std_logic;
  signal reg_q909_in     : std_logic;
  signal reg_q909_init   : std_logic;
		

  -- state q610
  signal reg_q610        : std_logic;
  signal reg_q610_in     : std_logic;
  signal reg_q610_init   : std_logic;
		

  -- state q612
  signal reg_q612        : std_logic;
  signal reg_q612_in     : std_logic;
  signal reg_q612_init   : std_logic;
		

  -- state q1462
  signal reg_q1462        : std_logic;
  signal reg_q1462_in     : std_logic;
  signal reg_q1462_init   : std_logic;
		

  -- state q123
  signal reg_q123        : std_logic;
  signal reg_q123_in     : std_logic;
  signal reg_q123_init   : std_logic;
		

  -- state q2213
  signal reg_q2213        : std_logic;
  signal reg_q2213_in     : std_logic;
  signal reg_q2213_init   : std_logic;
		

  -- state q426
  signal reg_q426        : std_logic;
  signal reg_q426_in     : std_logic;
  signal reg_q426_init   : std_logic;
		

  -- state q2405
  signal reg_q2405        : std_logic;
  signal reg_q2405_in     : std_logic;
  signal reg_q2405_init   : std_logic;
		

  -- state q2407
  signal reg_q2407        : std_logic;
  signal reg_q2407_in     : std_logic;
  signal reg_q2407_init   : std_logic;
		

  -- state q1470
  signal reg_q1470        : std_logic;
  signal reg_q1470_in     : std_logic;
  signal reg_q1470_init   : std_logic;
		

  -- state q2028
  signal reg_q2028        : std_logic;
  signal reg_q2028_in     : std_logic;
  signal reg_q2028_init   : std_logic;
		

  -- state q1217
  signal reg_q1217        : std_logic;
  signal reg_q1217_in     : std_logic;
  signal reg_q1217_init   : std_logic;
		

  -- state q1219
  signal reg_q1219        : std_logic;
  signal reg_q1219_in     : std_logic;
  signal reg_q1219_init   : std_logic;
		

  -- state q241
  signal reg_q241        : std_logic;
  signal reg_q241_in     : std_logic;
  signal reg_q241_init   : std_logic;
		

  -- state q1088
  signal reg_q1088        : std_logic;
  signal reg_q1088_in     : std_logic;
  signal reg_q1088_init   : std_logic;
		

  -- state q1090
  signal reg_q1090        : std_logic;
  signal reg_q1090_in     : std_logic;
  signal reg_q1090_init   : std_logic;
		

  -- state q1991
  signal reg_q1991        : std_logic;
  signal reg_q1991_in     : std_logic;
  signal reg_q1991_init   : std_logic;
		

  -- state q1993
  signal reg_q1993        : std_logic;
  signal reg_q1993_in     : std_logic;
  signal reg_q1993_init   : std_logic;
		

  -- state q1145
  signal reg_q1145        : std_logic;
  signal reg_q1145_in     : std_logic;
  signal reg_q1145_init   : std_logic;
		

  -- state q1147
  signal reg_q1147        : std_logic;
  signal reg_q1147_in     : std_logic;
  signal reg_q1147_init   : std_logic;
		

  -- state q1967
  signal reg_q1967        : std_logic;
  signal reg_q1967_in     : std_logic;
  signal reg_q1967_init   : std_logic;
		

  -- state q1969
  signal reg_q1969        : std_logic;
  signal reg_q1969_in     : std_logic;
  signal reg_q1969_init   : std_logic;
		

  -- state q1106
  signal reg_q1106        : std_logic;
  signal reg_q1106_in     : std_logic;
  signal reg_q1106_init   : std_logic;
		

  -- state q1205
  signal reg_q1205        : std_logic;
  signal reg_q1205_in     : std_logic;
  signal reg_q1205_init   : std_logic;
		

  -- state q524
  signal reg_q524        : std_logic;
  signal reg_q524_in     : std_logic;
  signal reg_q524_init   : std_logic;
		

  -- state q526
  signal reg_q526        : std_logic;
  signal reg_q526_in     : std_logic;
  signal reg_q526_init   : std_logic;
		

  -- state q1468
  signal reg_q1468        : std_logic;
  signal reg_q1468_in     : std_logic;
  signal reg_q1468_init   : std_logic;
		

  -- state q1672
  signal reg_q1672        : std_logic;
  signal reg_q1672_in     : std_logic;
  signal reg_q1672_init   : std_logic;
		

  -- state q1674
  signal reg_q1674        : std_logic;
  signal reg_q1674_in     : std_logic;
  signal reg_q1674_init   : std_logic;
		

  -- state q2375
  signal reg_q2375        : std_logic;
  signal reg_q2375_in     : std_logic;
  signal reg_q2375_init   : std_logic;
		

  -- state q2377
  signal reg_q2377        : std_logic;
  signal reg_q2377_in     : std_logic;
  signal reg_q2377_init   : std_logic;
		

  -- state q173
  signal reg_q173        : std_logic;
  signal reg_q173_in     : std_logic;
  signal reg_q173_init   : std_logic;
		

  -- state q175
  signal reg_q175        : std_logic;
  signal reg_q175_in     : std_logic;
  signal reg_q175_init   : std_logic;
		

  -- state q309
  signal reg_q309        : std_logic;
  signal reg_q309_in     : std_logic;
  signal reg_q309_init   : std_logic;
		

  -- state q311
  signal reg_q311        : std_logic;
  signal reg_q311_in     : std_logic;
  signal reg_q311_init   : std_logic;
		

  -- state q1421
  signal reg_q1421        : std_logic;
  signal reg_q1421_in     : std_logic;
  signal reg_q1421_init   : std_logic;
		

  -- state q1423
  signal reg_q1423        : std_logic;
  signal reg_q1423_in     : std_logic;
  signal reg_q1423_init   : std_logic;
		

  -- state q803
  signal reg_q803        : std_logic;
  signal reg_q803_in     : std_logic;
  signal reg_q803_init   : std_logic;
		

  -- state q805
  signal reg_q805        : std_logic;
  signal reg_q805_in     : std_logic;
  signal reg_q805_init   : std_logic;
		

  -- state q1335
  signal reg_q1335        : std_logic;
  signal reg_q1335_in     : std_logic;
  signal reg_q1335_init   : std_logic;
		

  -- state q2229
  signal reg_q2229        : std_logic;
  signal reg_q2229_in     : std_logic;
  signal reg_q2229_init   : std_logic;
		

  -- state q2093
  signal reg_q2093        : std_logic;
  signal reg_q2093_in     : std_logic;
  signal reg_q2093_init   : std_logic;
		

  -- state q1983
  signal reg_q1983        : std_logic;
  signal reg_q1983_in     : std_logic;
  signal reg_q1983_init   : std_logic;
		

  -- state q1985
  signal reg_q1985        : std_logic;
  signal reg_q1985_in     : std_logic;
  signal reg_q1985_init   : std_logic;
		

  -- state q1425
  signal reg_q1425        : std_logic;
  signal reg_q1425_in     : std_logic;
  signal reg_q1425_init   : std_logic;
		

  -- state q129
  signal reg_q129        : std_logic;
  signal reg_q129_in     : std_logic;
  signal reg_q129_init   : std_logic;
		

  -- state q1866
  signal reg_q1866        : std_logic;
  signal reg_q1866_in     : std_logic;
  signal reg_q1866_init   : std_logic;
		

  -- state q1868
  signal reg_q1868        : std_logic;
  signal reg_q1868_in     : std_logic;
  signal reg_q1868_init   : std_logic;
		

  -- state q2066
  signal reg_q2066        : std_logic;
  signal reg_q2066_in     : std_logic;
  signal reg_q2066_init   : std_logic;
		

  -- state q1341
  signal reg_q1341        : std_logic;
  signal reg_q1341_in     : std_logic;
  signal reg_q1341_init   : std_logic;
		

  -- state q2215
  signal reg_q2215        : std_logic;
  signal reg_q2215_in     : std_logic;
  signal reg_q2215_init   : std_logic;
		

  -- state q622
  signal reg_q622        : std_logic;
  signal reg_q622_in     : std_logic;
  signal reg_q622_init   : std_logic;
		

  -- state q624
  signal reg_q624        : std_logic;
  signal reg_q624_in     : std_logic;
  signal reg_q624_init   : std_logic;
		

  -- state q1840
  signal reg_q1840        : std_logic;
  signal reg_q1840_in     : std_logic;
  signal reg_q1840_init   : std_logic;
		

  -- state q1842
  signal reg_q1842        : std_logic;
  signal reg_q1842_in     : std_logic;
  signal reg_q1842_init   : std_logic;
		

  -- state q86
  signal reg_q86        : std_logic;
  signal reg_q86_in     : std_logic;
  signal reg_q86_init   : std_logic;
		

  -- state q1522
  signal reg_q1522        : std_logic;
  signal reg_q1522_in     : std_logic;
  signal reg_q1522_init   : std_logic;
		

  -- state q1523
  signal reg_q1523        : std_logic;
  signal reg_q1523_in     : std_logic;
  signal reg_q1523_init   : std_logic;
		

  -- state q1403
  signal reg_q1403        : std_logic;
  signal reg_q1403_in     : std_logic;
  signal reg_q1403_init   : std_logic;
		

  -- state q1405
  signal reg_q1405        : std_logic;
  signal reg_q1405_in     : std_logic;
  signal reg_q1405_init   : std_logic;
		

  -- state q2054
  signal reg_q2054        : std_logic;
  signal reg_q2054_in     : std_logic;
  signal reg_q2054_init   : std_logic;
		

  -- state q1541
  signal reg_q1541        : std_logic;
  signal reg_q1541_in     : std_logic;
  signal reg_q1541_init   : std_logic;
		

  -- state q2684
  signal reg_q2684        : std_logic;
  signal reg_q2684_in     : std_logic;
  signal reg_q2684_init   : std_logic;
		

  -- state q2686
  signal reg_q2686        : std_logic;
  signal reg_q2686_in     : std_logic;
  signal reg_q2686_init   : std_logic;
		

  -- state q1784
  signal reg_q1784        : std_logic;
  signal reg_q1784_in     : std_logic;
  signal reg_q1784_init   : std_logic;
		

  -- state q1786
  signal reg_q1786        : std_logic;
  signal reg_q1786_in     : std_logic;
  signal reg_q1786_init   : std_logic;
		

  -- state q2499
  signal reg_q2499        : std_logic;
  signal reg_q2499_in     : std_logic;
  signal reg_q2499_init   : std_logic;
		

  -- state q1906
  signal reg_q1906        : std_logic;
  signal reg_q1906_in     : std_logic;
  signal reg_q1906_init   : std_logic;
		

  -- state q1908
  signal reg_q1908        : std_logic;
  signal reg_q1908_in     : std_logic;
  signal reg_q1908_init   : std_logic;
		

  -- state q744
  signal reg_q744        : std_logic;
  signal reg_q744_in     : std_logic;
  signal reg_q744_init   : std_logic;
		

  -- state q746
  signal reg_q746        : std_logic;
  signal reg_q746_in     : std_logic;
  signal reg_q746_init   : std_logic;
		

  -- state q1131
  signal reg_q1131        : std_logic;
  signal reg_q1131_in     : std_logic;
  signal reg_q1131_init   : std_logic;
		

  -- state q1133
  signal reg_q1133        : std_logic;
  signal reg_q1133_in     : std_logic;
  signal reg_q1133_init   : std_logic;
		

  -- state q1454
  signal reg_q1454        : std_logic;
  signal reg_q1454_in     : std_logic;
  signal reg_q1454_init   : std_logic;
		

  -- state q1000
  signal reg_q1000        : std_logic;
  signal reg_q1000_in     : std_logic;
  signal reg_q1000_init   : std_logic;
		

  -- state q1002
  signal reg_q1002        : std_logic;
  signal reg_q1002_in     : std_logic;
  signal reg_q1002_init   : std_logic;
		

  -- state q1918
  signal reg_q1918        : std_logic;
  signal reg_q1918_in     : std_logic;
  signal reg_q1918_init   : std_logic;
		

  -- state q2280
  signal reg_q2280        : std_logic;
  signal reg_q2280_in     : std_logic;
  signal reg_q2280_init   : std_logic;
		

  -- state q2282
  signal reg_q2282        : std_logic;
  signal reg_q2282_in     : std_logic;
  signal reg_q2282_init   : std_logic;
		

  -- state q239
  signal reg_q239        : std_logic;
  signal reg_q239_in     : std_logic;
  signal reg_q239_init   : std_logic;
		

  -- state q2620
  signal reg_q2620        : std_logic;
  signal reg_q2620_in     : std_logic;
  signal reg_q2620_init   : std_logic;
		

  -- state q2622
  signal reg_q2622        : std_logic;
  signal reg_q2622_in     : std_logic;
  signal reg_q2622_init   : std_logic;
		

  -- state q2569
  signal reg_q2569        : std_logic;
  signal reg_q2569_in     : std_logic;
  signal reg_q2569_init   : std_logic;
		

  -- state q2571
  signal reg_q2571        : std_logic;
  signal reg_q2571_in     : std_logic;
  signal reg_q2571_init   : std_logic;
		

  -- state q2072
  signal reg_q2072        : std_logic;
  signal reg_q2072_in     : std_logic;
  signal reg_q2072_init   : std_logic;
		

  -- state q2074
  signal reg_q2074        : std_logic;
  signal reg_q2074_in     : std_logic;
  signal reg_q2074_init   : std_logic;
		

  -- state q1060
  signal reg_q1060        : std_logic;
  signal reg_q1060_in     : std_logic;
  signal reg_q1060_init   : std_logic;
		

  -- state q1062
  signal reg_q1062        : std_logic;
  signal reg_q1062_in     : std_logic;
  signal reg_q1062_init   : std_logic;
		

  -- state q133
  signal reg_q133        : std_logic;
  signal reg_q133_in     : std_logic;
  signal reg_q133_init   : std_logic;
		

  -- state q135
  signal reg_q135        : std_logic;
  signal reg_q135_in     : std_logic;
  signal reg_q135_init   : std_logic;
		

  -- state q341
  signal reg_q341        : std_logic;
  signal reg_q341_in     : std_logic;
  signal reg_q341_init   : std_logic;
		

  -- state q343
  signal reg_q343        : std_logic;
  signal reg_q343_in     : std_logic;
  signal reg_q343_init   : std_logic;
		

  -- state q797
  signal reg_q797        : std_logic;
  signal reg_q797_in     : std_logic;
  signal reg_q797_init   : std_logic;
		

  -- state q1301
  signal reg_q1301        : std_logic;
  signal reg_q1301_in     : std_logic;
  signal reg_q1301_init   : std_logic;
		

  -- state q1303
  signal reg_q1303        : std_logic;
  signal reg_q1303_in     : std_logic;
  signal reg_q1303_init   : std_logic;
		

  -- state q80
  signal reg_q80        : std_logic;
  signal reg_q80_in     : std_logic;
  signal reg_q80_init   : std_logic;
		

  -- state q82
  signal reg_q82        : std_logic;
  signal reg_q82_in     : std_logic;
  signal reg_q82_init   : std_logic;
		

  -- state q233
  signal reg_q233        : std_logic;
  signal reg_q233_in     : std_logic;
  signal reg_q233_init   : std_logic;
		

  -- state q840
  signal reg_q840        : std_logic;
  signal reg_q840_in     : std_logic;
  signal reg_q840_init   : std_logic;
		

  -- state q14
  signal reg_q14        : std_logic;
  signal reg_q14_in     : std_logic;
  signal reg_q14_init   : std_logic;
		

  -- state q16
  signal reg_q16        : std_logic;
  signal reg_q16_in     : std_logic;
  signal reg_q16_init   : std_logic;
		

  -- state q1333
  signal reg_q1333        : std_logic;
  signal reg_q1333_in     : std_logic;
  signal reg_q1333_init   : std_logic;
		

  -- state q2367
  signal reg_q2367        : std_logic;
  signal reg_q2367_in     : std_logic;
  signal reg_q2367_init   : std_logic;
		

  -- state q2369
  signal reg_q2369        : std_logic;
  signal reg_q2369_in     : std_logic;
  signal reg_q2369_init   : std_logic;
		

  -- state q1068
  signal reg_q1068        : std_logic;
  signal reg_q1068_in     : std_logic;
  signal reg_q1068_init   : std_logic;
		

  -- state q1070
  signal reg_q1070        : std_logic;
  signal reg_q1070_in     : std_logic;
  signal reg_q1070_init   : std_logic;
		

  -- state q732
  signal reg_q732        : std_logic;
  signal reg_q732_in     : std_logic;
  signal reg_q732_init   : std_logic;
		

  -- state q734
  signal reg_q734        : std_logic;
  signal reg_q734_in     : std_logic;
  signal reg_q734_init   : std_logic;
		

  -- state q1762
  signal reg_q1762        : std_logic;
  signal reg_q1762_in     : std_logic;
  signal reg_q1762_init   : std_logic;
		

  -- state q1764
  signal reg_q1764        : std_logic;
  signal reg_q1764_in     : std_logic;
  signal reg_q1764_init   : std_logic;
		

  -- state q1250
  signal reg_q1250        : std_logic;
  signal reg_q1250_in     : std_logic;
  signal reg_q1250_init   : std_logic;
		

  -- state q1252
  signal reg_q1252        : std_logic;
  signal reg_q1252_in     : std_logic;
  signal reg_q1252_init   : std_logic;
		

  -- state q1666
  signal reg_q1666        : std_logic;
  signal reg_q1666_in     : std_logic;
  signal reg_q1666_init   : std_logic;
		

  -- state q1127
  signal reg_q1127        : std_logic;
  signal reg_q1127_in     : std_logic;
  signal reg_q1127_init   : std_logic;
		

  -- state q1129
  signal reg_q1129        : std_logic;
  signal reg_q1129_in     : std_logic;
  signal reg_q1129_init   : std_logic;
		

  -- state q558
  signal reg_q558        : std_logic;
  signal reg_q558_in     : std_logic;
  signal reg_q558_init   : std_logic;
		

  -- state q560
  signal reg_q560        : std_logic;
  signal reg_q560_in     : std_logic;
  signal reg_q560_init   : std_logic;
		

  -- state q2415
  signal reg_q2415        : std_logic;
  signal reg_q2415_in     : std_logic;
  signal reg_q2415_init   : std_logic;
		

  -- state q2417
  signal reg_q2417        : std_logic;
  signal reg_q2417_in     : std_logic;
  signal reg_q2417_init   : std_logic;
		

  -- state q781
  signal reg_q781        : std_logic;
  signal reg_q781_in     : std_logic;
  signal reg_q781_init   : std_logic;
		

  -- state q397
  signal reg_q397        : std_logic;
  signal reg_q397_in     : std_logic;
  signal reg_q397_init   : std_logic;
		

  -- state q742
  signal reg_q742        : std_logic;
  signal reg_q742_in     : std_logic;
  signal reg_q742_init   : std_logic;
		

  -- state q2241
  signal reg_q2241        : std_logic;
  signal reg_q2241_in     : std_logic;
  signal reg_q2241_init   : std_logic;
		

  -- state q2243
  signal reg_q2243        : std_logic;
  signal reg_q2243_in     : std_logic;
  signal reg_q2243_init   : std_logic;
		

  -- state q251
  signal reg_q251        : std_logic;
  signal reg_q251_in     : std_logic;
  signal reg_q251_init   : std_logic;
		

  -- state q253
  signal reg_q253        : std_logic;
  signal reg_q253_in     : std_logic;
  signal reg_q253_init   : std_logic;
		

  -- state q1712
  signal reg_q1712        : std_logic;
  signal reg_q1712_in     : std_logic;
  signal reg_q1712_init   : std_logic;
		

  -- state q1714
  signal reg_q1714        : std_logic;
  signal reg_q1714_in     : std_logic;
  signal reg_q1714_init   : std_logic;
		

  -- state q371
  signal reg_q371        : std_logic;
  signal reg_q371_in     : std_logic;
  signal reg_q371_init   : std_logic;
		

  -- state q1756
  signal reg_q1756        : std_logic;
  signal reg_q1756_in     : std_logic;
  signal reg_q1756_init   : std_logic;
		

  -- state q1758
  signal reg_q1758        : std_logic;
  signal reg_q1758_in     : std_logic;
  signal reg_q1758_init   : std_logic;
		

  -- state q2468
  signal reg_q2468        : std_logic;
  signal reg_q2468_in     : std_logic;
  signal reg_q2468_init   : std_logic;
		

  -- state q2470
  signal reg_q2470        : std_logic;
  signal reg_q2470_in     : std_logic;
  signal reg_q2470_init   : std_logic;
		

  -- state q1696
  signal reg_q1696        : std_logic;
  signal reg_q1696_in     : std_logic;
  signal reg_q1696_init   : std_logic;
		

  -- state q1698
  signal reg_q1698        : std_logic;
  signal reg_q1698_in     : std_logic;
  signal reg_q1698_init   : std_logic;
		

  -- state q704
  signal reg_q704        : std_logic;
  signal reg_q704_in     : std_logic;
  signal reg_q704_init   : std_logic;
		

  -- state q901
  signal reg_q901        : std_logic;
  signal reg_q901_in     : std_logic;
  signal reg_q901_init   : std_logic;
		

  -- state q2624
  signal reg_q2624        : std_logic;
  signal reg_q2624_in     : std_logic;
  signal reg_q2624_init   : std_logic;
		

  -- state q962
  signal reg_q962        : std_logic;
  signal reg_q962_in     : std_logic;
  signal reg_q962_init   : std_logic;
		

  -- state q964
  signal reg_q964        : std_logic;
  signal reg_q964_in     : std_logic;
  signal reg_q964_init   : std_logic;
		

  -- state q424
  signal reg_q424        : std_logic;
  signal reg_q424_in     : std_logic;
  signal reg_q424_init   : std_logic;
		

  -- state q1822
  signal reg_q1822        : std_logic;
  signal reg_q1822_in     : std_logic;
  signal reg_q1822_init   : std_logic;
		

  -- state q1824
  signal reg_q1824        : std_logic;
  signal reg_q1824_in     : std_logic;
  signal reg_q1824_init   : std_logic;
		

  -- state q1317
  signal reg_q1317        : std_logic;
  signal reg_q1317_in     : std_logic;
  signal reg_q1317_init   : std_logic;
		

  -- state q1319
  signal reg_q1319        : std_logic;
  signal reg_q1319_in     : std_logic;
  signal reg_q1319_init   : std_logic;
		

  -- state q2577
  signal reg_q2577        : std_logic;
  signal reg_q2577_in     : std_logic;
  signal reg_q2577_init   : std_logic;
		

  -- state q620
  signal reg_q620        : std_logic;
  signal reg_q620_in     : std_logic;
  signal reg_q620_init   : std_logic;
		

  -- state q692
  signal reg_q692        : std_logic;
  signal reg_q692_in     : std_logic;
  signal reg_q692_init   : std_logic;
		

  -- state q367
  signal reg_q367        : std_logic;
  signal reg_q367_in     : std_logic;
  signal reg_q367_init   : std_logic;
		

  -- state q369
  signal reg_q369        : std_logic;
  signal reg_q369_in     : std_logic;
  signal reg_q369_init   : std_logic;
		

  -- state q2535
  signal reg_q2535        : std_logic;
  signal reg_q2535_in     : std_logic;
  signal reg_q2535_init   : std_logic;
		

  -- state q1221
  signal reg_q1221        : std_logic;
  signal reg_q1221_in     : std_logic;
  signal reg_q1221_init   : std_logic;
		

  -- state q1108
  signal reg_q1108        : std_logic;
  signal reg_q1108_in     : std_logic;
  signal reg_q1108_init   : std_logic;
		

  -- state q686
  signal reg_q686        : std_logic;
  signal reg_q686_in     : std_logic;
  signal reg_q686_init   : std_logic;
		

  -- state q1580
  signal reg_q1580        : std_logic;
  signal reg_q1580_in     : std_logic;
  signal reg_q1580_init   : std_logic;
		

  -- state q866
  signal reg_q866        : std_logic;
  signal reg_q866_in     : std_logic;
  signal reg_q866_init   : std_logic;
		

  -- state q868
  signal reg_q868        : std_logic;
  signal reg_q868_in     : std_logic;
  signal reg_q868_init   : std_logic;
		

  -- state q1371
  signal reg_q1371        : std_logic;
  signal reg_q1371_in     : std_logic;
  signal reg_q1371_init   : std_logic;
		

  -- state q1373
  signal reg_q1373        : std_logic;
  signal reg_q1373_in     : std_logic;
  signal reg_q1373_init   : std_logic;
		

  -- state q1558
  signal reg_q1558        : std_logic;
  signal reg_q1558_in     : std_logic;
  signal reg_q1558_init   : std_logic;
		

  -- state q1045
  signal reg_q1045        : std_logic;
  signal reg_q1045_in     : std_logic;
  signal reg_q1045_init   : std_logic;
		

  -- state q1047
  signal reg_q1047        : std_logic;
  signal reg_q1047_in     : std_logic;
  signal reg_q1047_init   : std_logic;
		

  -- state q2599
  signal reg_q2599        : std_logic;
  signal reg_q2599_in     : std_logic;
  signal reg_q2599_init   : std_logic;
		

  -- state q2016
  signal reg_q2016        : std_logic;
  signal reg_q2016_in     : std_logic;
  signal reg_q2016_init   : std_logic;
		

  -- state q2018
  signal reg_q2018        : std_logic;
  signal reg_q2018_in     : std_logic;
  signal reg_q2018_init   : std_logic;
		

  -- state q1989
  signal reg_q1989        : std_logic;
  signal reg_q1989_in     : std_logic;
  signal reg_q1989_init   : std_logic;
		

  -- state q2543
  signal reg_q2543        : std_logic;
  signal reg_q2543_in     : std_logic;
  signal reg_q2543_init   : std_logic;
		

  -- state q2545
  signal reg_q2545        : std_logic;
  signal reg_q2545_in     : std_logic;
  signal reg_q2545_init   : std_logic;
		

  -- state q1728
  signal reg_q1728        : std_logic;
  signal reg_q1728_in     : std_logic;
  signal reg_q1728_init   : std_logic;
		

  -- state q1730
  signal reg_q1730        : std_logic;
  signal reg_q1730_in     : std_logic;
  signal reg_q1730_init   : std_logic;
		

  -- state q438
  signal reg_q438        : std_logic;
  signal reg_q438_in     : std_logic;
  signal reg_q438_init   : std_logic;
		

  -- state q440
  signal reg_q440        : std_logic;
  signal reg_q440_in     : std_logic;
  signal reg_q440_init   : std_logic;
		

  -- state q772
  signal reg_q772        : std_logic;
  signal reg_q772_in     : std_logic;
  signal reg_q772_init   : std_logic;
		

  -- state q774
  signal reg_q774        : std_logic;
  signal reg_q774_in     : std_logic;
  signal reg_q774_init   : std_logic;
		

  -- state q2630
  signal reg_q2630        : std_logic;
  signal reg_q2630_in     : std_logic;
  signal reg_q2630_init   : std_logic;
		

  -- state q2632
  signal reg_q2632        : std_logic;
  signal reg_q2632_in     : std_logic;
  signal reg_q2632_init   : std_logic;
		

  -- state q528
  signal reg_q528        : std_logic;
  signal reg_q528_in     : std_logic;
  signal reg_q528_init   : std_logic;
		

  -- state q1963
  signal reg_q1963        : std_logic;
  signal reg_q1963_in     : std_logic;
  signal reg_q1963_init   : std_logic;
		

  -- state q1965
  signal reg_q1965        : std_logic;
  signal reg_q1965_in     : std_logic;
  signal reg_q1965_init   : std_logic;
		

  -- state q1264
  signal reg_q1264        : std_logic;
  signal reg_q1264_in     : std_logic;
  signal reg_q1264_init   : std_logic;
		

  -- state q1266
  signal reg_q1266        : std_logic;
  signal reg_q1266_in     : std_logic;
  signal reg_q1266_init   : std_logic;
		

  -- state q255
  signal reg_q255        : std_logic;
  signal reg_q255_in     : std_logic;
  signal reg_q255_init   : std_logic;
		

  -- state q596
  signal reg_q596        : std_logic;
  signal reg_q596_in     : std_logic;
  signal reg_q596_init   : std_logic;
		

  -- state q245
  signal reg_q245        : std_logic;
  signal reg_q245_in     : std_logic;
  signal reg_q245_init   : std_logic;
		

  -- state q2160
  signal reg_q2160        : std_logic;
  signal reg_q2160_in     : std_logic;
  signal reg_q2160_init   : std_logic;
		

  -- state q2573
  signal reg_q2573        : std_logic;
  signal reg_q2573_in     : std_logic;
  signal reg_q2573_init   : std_logic;
		

  -- state q1648
  signal reg_q1648        : std_logic;
  signal reg_q1648_in     : std_logic;
  signal reg_q1648_init   : std_logic;
		

  -- state q1650
  signal reg_q1650        : std_logic;
  signal reg_q1650_in     : std_logic;
  signal reg_q1650_init   : std_logic;
		

  -- state q2480
  signal reg_q2480        : std_logic;
  signal reg_q2480_in     : std_logic;
  signal reg_q2480_init   : std_logic;
		

  -- state q2482
  signal reg_q2482        : std_logic;
  signal reg_q2482_in     : std_logic;
  signal reg_q2482_init   : std_logic;
		

  -- state q107
  signal reg_q107        : std_logic;
  signal reg_q107_in     : std_logic;
  signal reg_q107_init   : std_logic;
		

  -- state q109
  signal reg_q109        : std_logic;
  signal reg_q109_in     : std_logic;
  signal reg_q109_init   : std_logic;
		

  -- state q1213
  signal reg_q1213        : std_logic;
  signal reg_q1213_in     : std_logic;
  signal reg_q1213_init   : std_logic;
		

  -- state q1215
  signal reg_q1215        : std_logic;
  signal reg_q1215_in     : std_logic;
  signal reg_q1215_init   : std_logic;
		

  -- state q2355
  signal reg_q2355        : std_logic;
  signal reg_q2355_in     : std_logic;
  signal reg_q2355_init   : std_logic;
		

  -- state q2357
  signal reg_q2357        : std_logic;
  signal reg_q2357_in     : std_logic;
  signal reg_q2357_init   : std_logic;
		

  -- state q1609
  signal reg_q1609        : std_logic;
  signal reg_q1609_in     : std_logic;
  signal reg_q1609_init   : std_logic;
		

  -- state q1611
  signal reg_q1611        : std_logic;
  signal reg_q1611_in     : std_logic;
  signal reg_q1611_init   : std_logic;
		

  -- state q2092
  signal reg_q2092        : std_logic;
  signal reg_q2092_in     : std_logic;
  signal reg_q2092_init   : std_logic;
		

  -- state q1613
  signal reg_q1613        : std_logic;
  signal reg_q1613_in     : std_logic;
  signal reg_q1613_init   : std_logic;
		

  -- state q2152
  signal reg_q2152        : std_logic;
  signal reg_q2152_in     : std_logic;
  signal reg_q2152_init   : std_logic;
		

  -- state q2154
  signal reg_q2154        : std_logic;
  signal reg_q2154_in     : std_logic;
  signal reg_q2154_init   : std_logic;
		

  -- state q1460
  signal reg_q1460        : std_logic;
  signal reg_q1460_in     : std_logic;
  signal reg_q1460_init   : std_logic;
		

  -- state q1339
  signal reg_q1339        : std_logic;
  signal reg_q1339_in     : std_logic;
  signal reg_q1339_init   : std_logic;
		

  -- state q2528
  signal reg_q2528        : std_logic;
  signal reg_q2528_in     : std_logic;
  signal reg_q2528_init   : std_logic;
		

  -- state q694
  signal reg_q694        : std_logic;
  signal reg_q694_in     : std_logic;
  signal reg_q694_init   : std_logic;
		

  -- state q1578
  signal reg_q1578        : std_logic;
  signal reg_q1578_in     : std_logic;
  signal reg_q1578_init   : std_logic;
		

  -- state q2520
  signal reg_q2520        : std_logic;
  signal reg_q2520_in     : std_logic;
  signal reg_q2520_init   : std_logic;
		

  -- state q2042
  signal reg_q2042        : std_logic;
  signal reg_q2042_in     : std_logic;
  signal reg_q2042_init   : std_logic;
		

  -- state q2044
  signal reg_q2044        : std_logic;
  signal reg_q2044_in     : std_logic;
  signal reg_q2044_init   : std_logic;
		

  -- state q2524
  signal reg_q2524        : std_logic;
  signal reg_q2524_in     : std_logic;
  signal reg_q2524_init   : std_logic;
		

  -- state q2526
  signal reg_q2526        : std_logic;
  signal reg_q2526_in     : std_logic;
  signal reg_q2526_init   : std_logic;
		

  -- state q1272
  signal reg_q1272        : std_logic;
  signal reg_q1272_in     : std_logic;
  signal reg_q1272_init   : std_logic;
		

  -- state q1274
  signal reg_q1274        : std_logic;
  signal reg_q1274_in     : std_logic;
  signal reg_q1274_init   : std_logic;
		

  -- state q111
  signal reg_q111        : std_logic;
  signal reg_q111_in     : std_logic;
  signal reg_q111_init   : std_logic;
		

  -- state q941
  signal reg_q941        : std_logic;
  signal reg_q941_in     : std_logic;
  signal reg_q941_init   : std_logic;
		

  -- state q943
  signal reg_q943        : std_logic;
  signal reg_q943_in     : std_logic;
  signal reg_q943_init   : std_logic;
		

  -- state q709
  signal reg_q709        : std_logic;
  signal reg_q709_in     : std_logic;
  signal reg_q709_init   : std_logic;
		

  -- state q711
  signal reg_q711        : std_logic;
  signal reg_q711_in     : std_logic;
  signal reg_q711_init   : std_logic;
		

  -- state q1226
  signal reg_q1226        : std_logic;
  signal reg_q1226_in     : std_logic;
  signal reg_q1226_init   : std_logic;
		

  -- state q1228
  signal reg_q1228        : std_logic;
  signal reg_q1228_in     : std_logic;
  signal reg_q1228_init   : std_logic;
		

  -- state q101
  signal reg_q101        : std_logic;
  signal reg_q101_in     : std_logic;
  signal reg_q101_init   : std_logic;
		

  -- state q103
  signal reg_q103        : std_logic;
  signal reg_q103_in     : std_logic;
  signal reg_q103_init   : std_logic;
		

  -- state q237
  signal reg_q237        : std_logic;
  signal reg_q237_in     : std_logic;
  signal reg_q237_init   : std_logic;
		

  -- state q226
  signal reg_q226        : std_logic;
  signal reg_q226_in     : std_logic;
  signal reg_q226_init   : std_logic;
		

  -- state q937
  signal reg_q937        : std_logic;
  signal reg_q937_in     : std_logic;
  signal reg_q937_init   : std_logic;
		

  -- state q939
  signal reg_q939        : std_logic;
  signal reg_q939_in     : std_logic;
  signal reg_q939_init   : std_logic;
		

  -- state q321
  signal reg_q321        : std_logic;
  signal reg_q321_in     : std_logic;
  signal reg_q321_init   : std_logic;
		

  -- state q323
  signal reg_q323        : std_logic;
  signal reg_q323_in     : std_logic;
  signal reg_q323_init   : std_logic;
		

  -- state q2253
  signal reg_q2253        : std_logic;
  signal reg_q2253_in     : std_logic;
  signal reg_q2253_init   : std_logic;
		

  -- state q2178
  signal reg_q2178        : std_logic;
  signal reg_q2178_in     : std_logic;
  signal reg_q2178_init   : std_logic;
		

  -- state q2180
  signal reg_q2180        : std_logic;
  signal reg_q2180_in     : std_logic;
  signal reg_q2180_init   : std_logic;
		

  -- state q2565
  signal reg_q2565        : std_logic;
  signal reg_q2565_in     : std_logic;
  signal reg_q2565_init   : std_logic;
		

  -- state q1443
  signal reg_q1443        : std_logic;
  signal reg_q1443_in     : std_logic;
  signal reg_q1443_init   : std_logic;
		

  -- state q1445
  signal reg_q1445        : std_logic;
  signal reg_q1445_in     : std_logic;
  signal reg_q1445_init   : std_logic;
		

  -- state q2148
  signal reg_q2148        : std_logic;
  signal reg_q2148_in     : std_logic;
  signal reg_q2148_init   : std_logic;
		

  -- state q590
  signal reg_q590        : std_logic;
  signal reg_q590_in     : std_logic;
  signal reg_q590_init   : std_logic;
		

  -- state q592
  signal reg_q592        : std_logic;
  signal reg_q592_in     : std_logic;
  signal reg_q592_init   : std_logic;
		

  -- state q949
  signal reg_q949        : std_logic;
  signal reg_q949_in     : std_logic;
  signal reg_q949_init   : std_logic;
		

  -- state q951
  signal reg_q951        : std_logic;
  signal reg_q951_in     : std_logic;
  signal reg_q951_init   : std_logic;
		

  -- state q1660
  signal reg_q1660        : std_logic;
  signal reg_q1660_in     : std_logic;
  signal reg_q1660_init   : std_logic;
		

  -- state q1113
  signal reg_q1113        : std_logic;
  signal reg_q1113_in     : std_logic;
  signal reg_q1113_init   : std_logic;
		

  -- state q974
  signal reg_q974        : std_logic;
  signal reg_q974_in     : std_logic;
  signal reg_q974_init   : std_logic;
		

  -- state q976
  signal reg_q976        : std_logic;
  signal reg_q976_in     : std_logic;
  signal reg_q976_init   : std_logic;
		

  -- state q84
  signal reg_q84        : std_logic;
  signal reg_q84_in     : std_logic;
  signal reg_q84_init   : std_logic;
		

  -- state q1902
  signal reg_q1902        : std_logic;
  signal reg_q1902_in     : std_logic;
  signal reg_q1902_init   : std_logic;
		

  -- state q1904
  signal reg_q1904        : std_logic;
  signal reg_q1904_in     : std_logic;
  signal reg_q1904_init   : std_logic;
		

  -- state q2613
  signal reg_q2613        : std_logic;
  signal reg_q2613_in     : std_logic;
  signal reg_q2613_init   : std_logic;
		

  -- state q532
  signal reg_q532        : std_logic;
  signal reg_q532_in     : std_logic;
  signal reg_q532_init   : std_logic;
		

  -- state q534
  signal reg_q534        : std_logic;
  signal reg_q534_in     : std_logic;
  signal reg_q534_init   : std_logic;
		

  -- state q1916
  signal reg_q1916        : std_logic;
  signal reg_q1916_in     : std_logic;
  signal reg_q1916_init   : std_logic;
		

  -- state q1498
  signal reg_q1498        : std_logic;
  signal reg_q1498_in     : std_logic;
  signal reg_q1498_init   : std_logic;
		

  -- state q1500
  signal reg_q1500        : std_logic;
  signal reg_q1500_in     : std_logic;
  signal reg_q1500_init   : std_logic;
		

  -- state q684
  signal reg_q684        : std_logic;
  signal reg_q684_in     : std_logic;
  signal reg_q684_init   : std_logic;
		

  -- state q2506
  signal reg_q2506        : std_logic;
  signal reg_q2506_in     : std_logic;
  signal reg_q2506_init   : std_logic;
		

  -- state q2508
  signal reg_q2508        : std_logic;
  signal reg_q2508_in     : std_logic;
  signal reg_q2508_init   : std_logic;
		

  -- state q1894
  signal reg_q1894        : std_logic;
  signal reg_q1894_in     : std_logic;
  signal reg_q1894_init   : std_logic;
		

  -- state q1896
  signal reg_q1896        : std_logic;
  signal reg_q1896_in     : std_logic;
  signal reg_q1896_init   : std_logic;
		

  -- state q304
  signal reg_q304        : std_logic;
  signal reg_q304_in     : std_logic;
  signal reg_q304_init   : std_logic;
		

  -- state q462
  signal reg_q462        : std_logic;
  signal reg_q462_in     : std_logic;
  signal reg_q462_init   : std_logic;
		

  -- state q464
  signal reg_q464        : std_logic;
  signal reg_q464_in     : std_logic;
  signal reg_q464_init   : std_logic;
		

  -- state q2646
  signal reg_q2646        : std_logic;
  signal reg_q2646_in     : std_logic;
  signal reg_q2646_init   : std_logic;
		

  -- state q2648
  signal reg_q2648        : std_logic;
  signal reg_q2648_in     : std_logic;
  signal reg_q2648_init   : std_logic;
		

  -- state q1149
  signal reg_q1149        : std_logic;
  signal reg_q1149_in     : std_logic;
  signal reg_q1149_init   : std_logic;
		

  -- state q2658
  signal reg_q2658        : std_logic;
  signal reg_q2658_in     : std_logic;
  signal reg_q2658_init   : std_logic;
		

  -- state q2660
  signal reg_q2660        : std_logic;
  signal reg_q2660_in     : std_logic;
  signal reg_q2660_init   : std_logic;
		

  -- state q1076
  signal reg_q1076        : std_logic;
  signal reg_q1076_in     : std_logic;
  signal reg_q1076_init   : std_logic;
		

  -- state q1078
  signal reg_q1078        : std_logic;
  signal reg_q1078_in     : std_logic;
  signal reg_q1078_init   : std_logic;
		

  -- state q658
  signal reg_q658        : std_logic;
  signal reg_q658_in     : std_logic;
  signal reg_q658_init   : std_logic;
		

  -- state q660
  signal reg_q660        : std_logic;
  signal reg_q660_in     : std_logic;
  signal reg_q660_init   : std_logic;
		

  -- state q418
  signal reg_q418        : std_logic;
  signal reg_q418_in     : std_logic;
  signal reg_q418_init   : std_logic;
		

  -- state q420
  signal reg_q420        : std_logic;
  signal reg_q420_in     : std_logic;
  signal reg_q420_init   : std_logic;
		

  -- state q1086
  signal reg_q1086        : std_logic;
  signal reg_q1086_in     : std_logic;
  signal reg_q1086_init   : std_logic;
		

  -- state q726
  signal reg_q726        : std_logic;
  signal reg_q726_in     : std_logic;
  signal reg_q726_init   : std_logic;
		

  -- state q728
  signal reg_q728        : std_logic;
  signal reg_q728_in     : std_logic;
  signal reg_q728_init   : std_logic;
		

  -- state q795
  signal reg_q795        : std_logic;
  signal reg_q795_in     : std_logic;
  signal reg_q795_init   : std_logic;
		

  -- state q978
  signal reg_q978        : std_logic;
  signal reg_q978_in     : std_logic;
  signal reg_q978_init   : std_logic;
		

  -- state q1778
  signal reg_q1778        : std_logic;
  signal reg_q1778_in     : std_logic;
  signal reg_q1778_init   : std_logic;
		

  -- state q1780
  signal reg_q1780        : std_logic;
  signal reg_q1780_in     : std_logic;
  signal reg_q1780_init   : std_logic;
		

  -- state q47
  signal reg_q47        : std_logic;
  signal reg_q47_in     : std_logic;
  signal reg_q47_init   : std_logic;
		

  -- state q48
  signal reg_q48        : std_logic;
  signal reg_q48_in     : std_logic;
  signal reg_q48_init   : std_logic;
		

  -- state q707
  signal reg_q707        : std_logic;
  signal reg_q707_in     : std_logic;
  signal reg_q707_init   : std_logic;
		

  -- state q1199
  signal reg_q1199        : std_logic;
  signal reg_q1199_in     : std_logic;
  signal reg_q1199_init   : std_logic;
		

  -- state q1201
  signal reg_q1201        : std_logic;
  signal reg_q1201_in     : std_logic;
  signal reg_q1201_init   : std_logic;
		

  -- state q2304
  signal reg_q2304        : std_logic;
  signal reg_q2304_in     : std_logic;
  signal reg_q2304_init   : std_logic;
		

  -- state q2306
  signal reg_q2306        : std_logic;
  signal reg_q2306_in     : std_logic;
  signal reg_q2306_init   : std_logic;
		

  -- state q448
  signal reg_q448        : std_logic;
  signal reg_q448_in     : std_logic;
  signal reg_q448_init   : std_logic;
		

  -- state q1453
  signal reg_q1453        : std_logic;
  signal reg_q1453_in     : std_logic;
  signal reg_q1453_init   : std_logic;
		

  -- state q1363
  signal reg_q1363        : std_logic;
  signal reg_q1363_in     : std_logic;
  signal reg_q1363_init   : std_logic;
		

  -- state q1365
  signal reg_q1365        : std_logic;
  signal reg_q1365_in     : std_logic;
  signal reg_q1365_init   : std_logic;
		

  -- state q1631
  signal reg_q1631        : std_logic;
  signal reg_q1631_in     : std_logic;
  signal reg_q1631_init   : std_logic;
		

  -- state q1633
  signal reg_q1633        : std_logic;
  signal reg_q1633_in     : std_logic;
  signal reg_q1633_init   : std_logic;
		

  -- state q1790
  signal reg_q1790        : std_logic;
  signal reg_q1790_in     : std_logic;
  signal reg_q1790_init   : std_logic;
		

  -- state q1792
  signal reg_q1792        : std_logic;
  signal reg_q1792_in     : std_logic;
  signal reg_q1792_init   : std_logic;
		

  -- state q836
  signal reg_q836        : std_logic;
  signal reg_q836_in     : std_logic;
  signal reg_q836_init   : std_logic;
		

  -- state q1539
  signal reg_q1539        : std_logic;
  signal reg_q1539_in     : std_logic;
  signal reg_q1539_init   : std_logic;
		

  -- state q510
  signal reg_q510        : std_logic;
  signal reg_q510_in     : std_logic;
  signal reg_q510_init   : std_logic;
		

  -- state q512
  signal reg_q512        : std_logic;
  signal reg_q512_in     : std_logic;
  signal reg_q512_init   : std_logic;
		

  -- state q1284
  signal reg_q1284        : std_logic;
  signal reg_q1284_in     : std_logic;
  signal reg_q1284_init   : std_logic;
		

  -- state q1286
  signal reg_q1286        : std_logic;
  signal reg_q1286_in     : std_logic;
  signal reg_q1286_init   : std_logic;
		

  -- state q1256
  signal reg_q1256        : std_logic;
  signal reg_q1256_in     : std_logic;
  signal reg_q1256_init   : std_logic;
		

  -- state q1258
  signal reg_q1258        : std_logic;
  signal reg_q1258_in     : std_logic;
  signal reg_q1258_init   : std_logic;
		

  -- state q113
  signal reg_q113        : std_logic;
  signal reg_q113_in     : std_logic;
  signal reg_q113_init   : std_logic;
		

  -- state q1987
  signal reg_q1987        : std_logic;
  signal reg_q1987_in     : std_logic;
  signal reg_q1987_init   : std_logic;
		

  -- state q298
  signal reg_q298        : std_logic;
  signal reg_q298_in     : std_logic;
  signal reg_q298_init   : std_logic;
		

  -- state q300
  signal reg_q300        : std_logic;
  signal reg_q300_in     : std_logic;
  signal reg_q300_init   : std_logic;
		

  -- state q1025
  signal reg_q1025        : std_logic;
  signal reg_q1025_in     : std_logic;
  signal reg_q1025_init   : std_logic;
		

  -- state q1027
  signal reg_q1027        : std_logic;
  signal reg_q1027_in     : std_logic;
  signal reg_q1027_init   : std_logic;
		

  -- state q179
  signal reg_q179        : std_logic;
  signal reg_q179_in     : std_logic;
  signal reg_q179_init   : std_logic;
		

  -- state q1621
  signal reg_q1621        : std_logic;
  signal reg_q1621_in     : std_logic;
  signal reg_q1621_init   : std_logic;
		

  -- state q1623
  signal reg_q1623        : std_logic;
  signal reg_q1623_in     : std_logic;
  signal reg_q1623_init   : std_logic;
		

  -- state q766
  signal reg_q766        : std_logic;
  signal reg_q766_in     : std_logic;
  signal reg_q766_init   : std_logic;
		

  -- state q768
  signal reg_q768        : std_logic;
  signal reg_q768_in     : std_logic;
  signal reg_q768_init   : std_logic;
		

  -- state q1752
  signal reg_q1752        : std_logic;
  signal reg_q1752_in     : std_logic;
  signal reg_q1752_init   : std_logic;
		

  -- state q1754
  signal reg_q1754        : std_logic;
  signal reg_q1754_in     : std_logic;
  signal reg_q1754_init   : std_logic;
		

  -- state q1072
  signal reg_q1072        : std_logic;
  signal reg_q1072_in     : std_logic;
  signal reg_q1072_init   : std_logic;
		

  -- state q2324
  signal reg_q2324        : std_logic;
  signal reg_q2324_in     : std_logic;
  signal reg_q2324_init   : std_logic;
		

  -- state q1850
  signal reg_q1850        : std_logic;
  signal reg_q1850_in     : std_logic;
  signal reg_q1850_init   : std_logic;
		

  -- state q1852
  signal reg_q1852        : std_logic;
  signal reg_q1852_in     : std_logic;
  signal reg_q1852_init   : std_logic;
		

  -- state q137
  signal reg_q137        : std_logic;
  signal reg_q137_in     : std_logic;
  signal reg_q137_init   : std_logic;
		

  -- state q139
  signal reg_q139        : std_logic;
  signal reg_q139_in     : std_logic;
  signal reg_q139_init   : std_logic;
		

  -- state q2278
  signal reg_q2278        : std_logic;
  signal reg_q2278_in     : std_logic;
  signal reg_q2278_init   : std_logic;
		

  -- state q286
  signal reg_q286        : std_logic;
  signal reg_q286_in     : std_logic;
  signal reg_q286_init   : std_logic;
		

  -- state q288
  signal reg_q288        : std_logic;
  signal reg_q288_in     : std_logic;
  signal reg_q288_init   : std_logic;
		

  -- state q614
  signal reg_q614        : std_logic;
  signal reg_q614_in     : std_logic;
  signal reg_q614_init   : std_logic;
		

  -- state q887
  signal reg_q887        : std_logic;
  signal reg_q887_in     : std_logic;
  signal reg_q887_init   : std_logic;
		

  -- state q231
  signal reg_q231        : std_logic;
  signal reg_q231_in     : std_logic;
  signal reg_q231_init   : std_logic;
		

  -- state q2429
  signal reg_q2429        : std_logic;
  signal reg_q2429_in     : std_logic;
  signal reg_q2429_init   : std_logic;
		

  -- state q2431
  signal reg_q2431        : std_logic;
  signal reg_q2431_in     : std_logic;
  signal reg_q2431_init   : std_logic;
		

  -- state q1545
  signal reg_q1545        : std_logic;
  signal reg_q1545_in     : std_logic;
  signal reg_q1545_init   : std_logic;
		

  -- state q1546
  signal reg_q1546        : std_logic;
  signal reg_q1546_in     : std_logic;
  signal reg_q1546_init   : std_logic;
		

  -- state q1806
  signal reg_q1806        : std_logic;
  signal reg_q1806_in     : std_logic;
  signal reg_q1806_init   : std_logic;
		

  -- state q1808
  signal reg_q1808        : std_logic;
  signal reg_q1808_in     : std_logic;
  signal reg_q1808_init   : std_logic;
		

  -- state q2202
  signal reg_q2202        : std_logic;
  signal reg_q2202_in     : std_logic;
  signal reg_q2202_init   : std_logic;
		

  -- state q2204
  signal reg_q2204        : std_logic;
  signal reg_q2204_in     : std_logic;
  signal reg_q2204_init   : std_logic;
		

  -- state q1554
  signal reg_q1554        : std_logic;
  signal reg_q1554_in     : std_logic;
  signal reg_q1554_init   : std_logic;
		

  -- state q1556
  signal reg_q1556        : std_logic;
  signal reg_q1556_in     : std_logic;
  signal reg_q1556_init   : std_logic;
		

  -- state q1882
  signal reg_q1882        : std_logic;
  signal reg_q1882_in     : std_logic;
  signal reg_q1882_init   : std_logic;
		

  -- state q1165
  signal reg_q1165        : std_logic;
  signal reg_q1165_in     : std_logic;
  signal reg_q1165_init   : std_logic;
		

  -- state q1167
  signal reg_q1167        : std_logic;
  signal reg_q1167_in     : std_logic;
  signal reg_q1167_init   : std_logic;
		

  -- state q1846
  signal reg_q1846        : std_logic;
  signal reg_q1846_in     : std_logic;
  signal reg_q1846_init   : std_logic;
		

  -- state q884
  signal reg_q884        : std_logic;
  signal reg_q884_in     : std_logic;
  signal reg_q884_init   : std_logic;
		

  -- state q2537
  signal reg_q2537        : std_logic;
  signal reg_q2537_in     : std_logic;
  signal reg_q2537_init   : std_logic;
		

  -- state q149
  signal reg_q149        : std_logic;
  signal reg_q149_in     : std_logic;
  signal reg_q149_init   : std_logic;
		

  -- state q151
  signal reg_q151        : std_logic;
  signal reg_q151_in     : std_logic;
  signal reg_q151_init   : std_logic;
		

  -- state q1173
  signal reg_q1173        : std_logic;
  signal reg_q1173_in     : std_logic;
  signal reg_q1173_init   : std_logic;
		

  -- state q1175
  signal reg_q1175        : std_logic;
  signal reg_q1175_in     : std_logic;
  signal reg_q1175_init   : std_logic;
		

  -- state q2351
  signal reg_q2351        : std_logic;
  signal reg_q2351_in     : std_logic;
  signal reg_q2351_init   : std_logic;
		

  -- state q2553
  signal reg_q2553        : std_logic;
  signal reg_q2553_in     : std_logic;
  signal reg_q2553_init   : std_logic;
		

  -- state q2555
  signal reg_q2555        : std_logic;
  signal reg_q2555_in     : std_logic;
  signal reg_q2555_init   : std_logic;
		

  -- state q20
  signal reg_q20        : std_logic;
  signal reg_q20_in     : std_logic;
  signal reg_q20_init   : std_logic;
		

  -- state q2245
  signal reg_q2245        : std_logic;
  signal reg_q2245_in     : std_logic;
  signal reg_q2245_init   : std_logic;
		

  -- state q1041
  signal reg_q1041        : std_logic;
  signal reg_q1041_in     : std_logic;
  signal reg_q1041_init   : std_logic;
		

  -- state q1043
  signal reg_q1043        : std_logic;
  signal reg_q1043_in     : std_logic;
  signal reg_q1043_init   : std_logic;
		

  -- state q1981
  signal reg_q1981        : std_logic;
  signal reg_q1981_in     : std_logic;
  signal reg_q1981_init   : std_logic;
		

  -- state q2276
  signal reg_q2276        : std_logic;
  signal reg_q2276_in     : std_logic;
  signal reg_q2276_init   : std_logic;
		

  -- state q1288
  signal reg_q1288        : std_logic;
  signal reg_q1288_in     : std_logic;
  signal reg_q1288_init   : std_logic;
		

  -- state q602
  signal reg_q602        : std_logic;
  signal reg_q602_in     : std_logic;
  signal reg_q602_init   : std_logic;
		

  -- state q604
  signal reg_q604        : std_logic;
  signal reg_q604_in     : std_logic;
  signal reg_q604_init   : std_logic;
		

  -- state q2034
  signal reg_q2034        : std_logic;
  signal reg_q2034_in     : std_logic;
  signal reg_q2034_init   : std_logic;
		

  -- state q1006
  signal reg_q1006        : std_logic;
  signal reg_q1006_in     : std_logic;
  signal reg_q1006_init   : std_logic;
		

  -- state q1008
  signal reg_q1008        : std_logic;
  signal reg_q1008_in     : std_logic;
  signal reg_q1008_init   : std_logic;
		

  -- state q266
  signal reg_q266        : std_logic;
  signal reg_q266_in     : std_logic;
  signal reg_q266_init   : std_logic;
		

  -- state q268
  signal reg_q268        : std_logic;
  signal reg_q268_in     : std_logic;
  signal reg_q268_init   : std_logic;
		

  -- state q2333
  signal reg_q2333        : std_logic;
  signal reg_q2333_in     : std_logic;
  signal reg_q2333_init   : std_logic;
		

  -- state q2335
  signal reg_q2335        : std_logic;
  signal reg_q2335_in     : std_logic;
  signal reg_q2335_init   : std_logic;
		

  -- state q1211
  signal reg_q1211        : std_logic;
  signal reg_q1211_in     : std_logic;
  signal reg_q1211_init   : std_logic;
		

  -- state q1197
  signal reg_q1197        : std_logic;
  signal reg_q1197_in     : std_logic;
  signal reg_q1197_init   : std_logic;
		

  -- state q1242
  signal reg_q1242        : std_logic;
  signal reg_q1242_in     : std_logic;
  signal reg_q1242_init   : std_logic;
		

  -- state q1244
  signal reg_q1244        : std_logic;
  signal reg_q1244_in     : std_logic;
  signal reg_q1244_init   : std_logic;
		

  -- state q198
  signal reg_q198        : std_logic;
  signal reg_q198_in     : std_logic;
  signal reg_q198_init   : std_logic;
		

  -- state q200
  signal reg_q200        : std_logic;
  signal reg_q200_in     : std_logic;
  signal reg_q200_init   : std_logic;
		

  -- state q2487
  signal reg_q2487        : std_logic;
  signal reg_q2487_in     : std_logic;
  signal reg_q2487_init   : std_logic;
		

  -- state q2489
  signal reg_q2489        : std_logic;
  signal reg_q2489_in     : std_logic;
  signal reg_q2489_init   : std_logic;
		

  -- state q2268
  signal reg_q2268        : std_logic;
  signal reg_q2268_in     : std_logic;
  signal reg_q2268_init   : std_logic;
		

  -- state q2270
  signal reg_q2270        : std_logic;
  signal reg_q2270_in     : std_logic;
  signal reg_q2270_init   : std_logic;
		

  -- state q243
  signal reg_q243        : std_logic;
  signal reg_q243_in     : std_logic;
  signal reg_q243_init   : std_logic;
		

  -- state q1056
  signal reg_q1056        : std_logic;
  signal reg_q1056_in     : std_logic;
  signal reg_q1056_init   : std_logic;
		

  -- state q1058
  signal reg_q1058        : std_logic;
  signal reg_q1058_in     : std_logic;
  signal reg_q1058_init   : std_logic;
		

  -- state q1115
  signal reg_q1115        : std_logic;
  signal reg_q1115_in     : std_logic;
  signal reg_q1115_init   : std_logic;
		

  -- state q1117
  signal reg_q1117        : std_logic;
  signal reg_q1117_in     : std_logic;
  signal reg_q1117_init   : std_logic;
		

  -- state q1135
  signal reg_q1135        : std_logic;
  signal reg_q1135_in     : std_logic;
  signal reg_q1135_init   : std_logic;
		

  -- state q864
  signal reg_q864        : std_logic;
  signal reg_q864_in     : std_logic;
  signal reg_q864_init   : std_logic;
		

  -- state q2048
  signal reg_q2048        : std_logic;
  signal reg_q2048_in     : std_logic;
  signal reg_q2048_init   : std_logic;
		

  -- state q2050
  signal reg_q2050        : std_logic;
  signal reg_q2050_in     : std_logic;
  signal reg_q2050_init   : std_logic;
		

  -- state q2113
  signal reg_q2113        : std_logic;
  signal reg_q2113_in     : std_logic;
  signal reg_q2113_init   : std_logic;
		

  -- state q2115
  signal reg_q2115        : std_logic;
  signal reg_q2115_in     : std_logic;
  signal reg_q2115_init   : std_logic;
		

  -- state q2095
  signal reg_q2095        : std_logic;
  signal reg_q2095_in     : std_logic;
  signal reg_q2095_init   : std_logic;
		

  -- state q2097
  signal reg_q2097        : std_logic;
  signal reg_q2097_in     : std_logic;
  signal reg_q2097_init   : std_logic;
		

  -- state q145
  signal reg_q145        : std_logic;
  signal reg_q145_in     : std_logic;
  signal reg_q145_init   : std_logic;
		

  -- state q147
  signal reg_q147        : std_logic;
  signal reg_q147_in     : std_logic;
  signal reg_q147_init   : std_logic;
		

  -- state q900
  signal reg_q900        : std_logic;
  signal reg_q900_in     : std_logic;
  signal reg_q900_init   : std_logic;
		

  -- state q2233
  signal reg_q2233        : std_logic;
  signal reg_q2233_in     : std_logic;
  signal reg_q2233_init   : std_logic;
		

  -- state q2235
  signal reg_q2235        : std_logic;
  signal reg_q2235_in     : std_logic;
  signal reg_q2235_init   : std_logic;
		

  -- state q1104
  signal reg_q1104        : std_logic;
  signal reg_q1104_in     : std_logic;
  signal reg_q1104_init   : std_logic;
		

  -- state q1482
  signal reg_q1482        : std_logic;
  signal reg_q1482_in     : std_logic;
  signal reg_q1482_init   : std_logic;
		

  -- state q715
  signal reg_q715        : std_logic;
  signal reg_q715_in     : std_logic;
  signal reg_q715_init   : std_logic;
		

  -- state q716
  signal reg_q716        : std_logic;
  signal reg_q716_in     : std_logic;
  signal reg_q716_init   : std_logic;
		

  -- state q514
  signal reg_q514        : std_logic;
  signal reg_q514_in     : std_logic;
  signal reg_q514_init   : std_logic;
		

  -- state q516
  signal reg_q516        : std_logic;
  signal reg_q516_in     : std_logic;
  signal reg_q516_init   : std_logic;
		

  -- state q24
  signal reg_q24        : std_logic;
  signal reg_q24_in     : std_logic;
  signal reg_q24_init   : std_logic;
		

  -- state q26
  signal reg_q26        : std_logic;
  signal reg_q26_in     : std_logic;
  signal reg_q26_init   : std_logic;
		

  -- state q454
  signal reg_q454        : std_logic;
  signal reg_q454_in     : std_logic;
  signal reg_q454_init   : std_logic;
		

  -- state q752
  signal reg_q752        : std_logic;
  signal reg_q752_in     : std_logic;
  signal reg_q752_init   : std_logic;
		

  -- state q754
  signal reg_q754        : std_logic;
  signal reg_q754_in     : std_logic;
  signal reg_q754_init   : std_logic;
		

  -- state q1720
  signal reg_q1720        : std_logic;
  signal reg_q1720_in     : std_logic;
  signal reg_q1720_init   : std_logic;
		

  -- state q1886
  signal reg_q1886        : std_logic;
  signal reg_q1886_in     : std_logic;
  signal reg_q1886_init   : std_logic;
		

  -- state q2164
  signal reg_q2164        : std_logic;
  signal reg_q2164_in     : std_logic;
  signal reg_q2164_init   : std_logic;
		

  -- state q2166
  signal reg_q2166        : std_logic;
  signal reg_q2166_in     : std_logic;
  signal reg_q2166_init   : std_logic;
		

  -- state q1435
  signal reg_q1435        : std_logic;
  signal reg_q1435_in     : std_logic;
  signal reg_q1435_init   : std_logic;
		

  -- state q1437
  signal reg_q1437        : std_logic;
  signal reg_q1437_in     : std_logic;
  signal reg_q1437_init   : std_logic;
		

  -- state q1810
  signal reg_q1810        : std_logic;
  signal reg_q1810_in     : std_logic;
  signal reg_q1810_init   : std_logic;
		

  -- state q1254
  signal reg_q1254        : std_logic;
  signal reg_q1254_in     : std_logic;
  signal reg_q1254_init   : std_logic;
		

  -- state q1652
  signal reg_q1652        : std_logic;
  signal reg_q1652_in     : std_logic;
  signal reg_q1652_init   : std_logic;
		

  -- state q1654
  signal reg_q1654        : std_logic;
  signal reg_q1654_in     : std_logic;
  signal reg_q1654_init   : std_logic;
		

  -- state q1327
  signal reg_q1327        : std_logic;
  signal reg_q1327_in     : std_logic;
  signal reg_q1327_init   : std_logic;
		

  -- state q1329
  signal reg_q1329        : std_logic;
  signal reg_q1329_in     : std_logic;
  signal reg_q1329_init   : std_logic;
		

  -- state q2070
  signal reg_q2070        : std_logic;
  signal reg_q2070_in     : std_logic;
  signal reg_q2070_init   : std_logic;
		

  -- state q1125
  signal reg_q1125        : std_logic;
  signal reg_q1125_in     : std_logic;
  signal reg_q1125_init   : std_logic;
		

  -- state q2409
  signal reg_q2409        : std_logic;
  signal reg_q2409_in     : std_logic;
  signal reg_q2409_init   : std_logic;
		

  -- state q986
  signal reg_q986        : std_logic;
  signal reg_q986_in     : std_logic;
  signal reg_q986_init   : std_logic;
		

  -- state q1794
  signal reg_q1794        : std_logic;
  signal reg_q1794_in     : std_logic;
  signal reg_q1794_init   : std_logic;
		

  -- state q1796
  signal reg_q1796        : std_logic;
  signal reg_q1796_in     : std_logic;
  signal reg_q1796_init   : std_logic;
		

  -- state q385
  signal reg_q385        : std_logic;
  signal reg_q385_in     : std_logic;
  signal reg_q385_init   : std_logic;
		

  -- state q387
  signal reg_q387        : std_logic;
  signal reg_q387_in     : std_logic;
  signal reg_q387_init   : std_logic;
		

  -- state q1490
  signal reg_q1490        : std_logic;
  signal reg_q1490_in     : std_logic;
  signal reg_q1490_init   : std_logic;
		

  -- state q1922
  signal reg_q1922        : std_logic;
  signal reg_q1922_in     : std_logic;
  signal reg_q1922_init   : std_logic;
		

  -- state q1924
  signal reg_q1924        : std_logic;
  signal reg_q1924_in     : std_logic;
  signal reg_q1924_init   : std_logic;
		

  -- state q862
  signal reg_q862        : std_logic;
  signal reg_q862_in     : std_logic;
  signal reg_q862_init   : std_logic;
		

  -- state q2258
  signal reg_q2258        : std_logic;
  signal reg_q2258_in     : std_logic;
  signal reg_q2258_init   : std_logic;
		

  -- state q1433
  signal reg_q1433        : std_logic;
  signal reg_q1433_in     : std_logic;
  signal reg_q1433_init   : std_logic;
		

  -- state q1920
  signal reg_q1920        : std_logic;
  signal reg_q1920_in     : std_logic;
  signal reg_q1920_init   : std_logic;
		

  -- state q2341
  signal reg_q2341        : std_logic;
  signal reg_q2341_in     : std_logic;
  signal reg_q2341_init   : std_logic;
		

  -- state q2343
  signal reg_q2343        : std_logic;
  signal reg_q2343_in     : std_logic;
  signal reg_q2343_init   : std_logic;
		

  -- state q1309
  signal reg_q1309        : std_logic;
  signal reg_q1309_in     : std_logic;
  signal reg_q1309_init   : std_logic;
		

  -- state q1311
  signal reg_q1311        : std_logic;
  signal reg_q1311_in     : std_logic;
  signal reg_q1311_init   : std_logic;
		

  -- state q2286
  signal reg_q2286        : std_logic;
  signal reg_q2286_in     : std_logic;
  signal reg_q2286_init   : std_logic;
		

  -- state q325
  signal reg_q325        : std_logic;
  signal reg_q325_in     : std_logic;
  signal reg_q325_init   : std_logic;
		

  -- state q327
  signal reg_q327        : std_logic;
  signal reg_q327_in     : std_logic;
  signal reg_q327_init   : std_logic;
		

  -- state q2247
  signal reg_q2247        : std_logic;
  signal reg_q2247_in     : std_logic;
  signal reg_q2247_init   : std_logic;
		

  -- state q1193
  signal reg_q1193        : std_logic;
  signal reg_q1193_in     : std_logic;
  signal reg_q1193_init   : std_logic;
		

  -- state q450
  signal reg_q450        : std_logic;
  signal reg_q450_in     : std_logic;
  signal reg_q450_init   : std_logic;
		

  -- state q911
  signal reg_q911        : std_logic;
  signal reg_q911_in     : std_logic;
  signal reg_q911_init   : std_logic;
		

  -- state q980
  signal reg_q980        : std_logic;
  signal reg_q980_in     : std_logic;
  signal reg_q980_init   : std_logic;
		

  -- state q1268
  signal reg_q1268        : std_logic;
  signal reg_q1268_in     : std_logic;
  signal reg_q1268_init   : std_logic;
		

  -- state q1270
  signal reg_q1270        : std_logic;
  signal reg_q1270_in     : std_logic;
  signal reg_q1270_init   : std_logic;
		

  -- state q305
  signal reg_q305        : std_logic;
  signal reg_q305_in     : std_logic;
  signal reg_q305_init   : std_logic;
		

  -- state q988
  signal reg_q988        : std_logic;
  signal reg_q988_in     : std_logic;
  signal reg_q988_init   : std_logic;
		

  -- state q990
  signal reg_q990        : std_logic;
  signal reg_q990_in     : std_logic;
  signal reg_q990_init   : std_logic;
		

  -- state q1750
  signal reg_q1750        : std_logic;
  signal reg_q1750_in     : std_logic;
  signal reg_q1750_init   : std_logic;
		

  -- state q1419
  signal reg_q1419        : std_logic;
  signal reg_q1419_in     : std_logic;
  signal reg_q1419_init   : std_logic;
		

  -- state q1854
  signal reg_q1854        : std_logic;
  signal reg_q1854_in     : std_logic;
  signal reg_q1854_init   : std_logic;
		

  -- state q88
  signal reg_q88        : std_logic;
  signal reg_q88_in     : std_logic;
  signal reg_q88_init   : std_logic;
		

  -- state q1800
  signal reg_q1800        : std_logic;
  signal reg_q1800_in     : std_logic;
  signal reg_q1800_init   : std_logic;
		

  -- state q1802
  signal reg_q1802        : std_logic;
  signal reg_q1802_in     : std_logic;
  signal reg_q1802_init   : std_logic;
		

  -- state q2002
  signal reg_q2002        : std_logic;
  signal reg_q2002_in     : std_logic;
  signal reg_q2002_init   : std_logic;
		

  -- state q2296
  signal reg_q2296        : std_logic;
  signal reg_q2296_in     : std_logic;
  signal reg_q2296_init   : std_logic;
		

  -- state q2298
  signal reg_q2298        : std_logic;
  signal reg_q2298_in     : std_logic;
  signal reg_q2298_init   : std_logic;
		

  -- state q966
  signal reg_q966        : std_logic;
  signal reg_q966_in     : std_logic;
  signal reg_q966_init   : std_logic;
		

  -- state q2652
  signal reg_q2652        : std_logic;
  signal reg_q2652_in     : std_logic;
  signal reg_q2652_init   : std_logic;
		

  -- state q2654
  signal reg_q2654        : std_logic;
  signal reg_q2654_in     : std_logic;
  signal reg_q2654_init   : std_logic;
		

  -- state q1938
  signal reg_q1938        : std_logic;
  signal reg_q1938_in     : std_logic;
  signal reg_q1938_init   : std_logic;
		

  -- state q1102
  signal reg_q1102        : std_logic;
  signal reg_q1102_in     : std_logic;
  signal reg_q1102_init   : std_logic;
		

  -- state q1766
  signal reg_q1766        : std_logic;
  signal reg_q1766_in     : std_logic;
  signal reg_q1766_init   : std_logic;
		

  -- state q1407
  signal reg_q1407        : std_logic;
  signal reg_q1407_in     : std_logic;
  signal reg_q1407_init   : std_logic;
		

  -- state q1409
  signal reg_q1409        : std_logic;
  signal reg_q1409_in     : std_logic;
  signal reg_q1409_init   : std_logic;
		

  -- state q235
  signal reg_q235        : std_logic;
  signal reg_q235_in     : std_logic;
  signal reg_q235_init   : std_logic;
		

  -- state q1381
  signal reg_q1381        : std_logic;
  signal reg_q1381_in     : std_logic;
  signal reg_q1381_init   : std_logic;
		

  -- state q1383
  signal reg_q1383        : std_logic;
  signal reg_q1383_in     : std_logic;
  signal reg_q1383_init   : std_logic;
		

  -- state q2642
  signal reg_q2642        : std_logic;
  signal reg_q2642_in     : std_logic;
  signal reg_q2642_init   : std_logic;
		

  -- state q2644
  signal reg_q2644        : std_logic;
  signal reg_q2644_in     : std_logic;
  signal reg_q2644_init   : std_logic;
		

  -- state q740
  signal reg_q740        : std_logic;
  signal reg_q740_in     : std_logic;
  signal reg_q740_init   : std_logic;
		

  -- state q1369
  signal reg_q1369        : std_logic;
  signal reg_q1369_in     : std_logic;
  signal reg_q1369_init   : std_logic;
		

  -- state q2399
  signal reg_q2399        : std_logic;
  signal reg_q2399_in     : std_logic;
  signal reg_q2399_init   : std_logic;
		

  -- state q2401
  signal reg_q2401        : std_logic;
  signal reg_q2401_in     : std_logic;
  signal reg_q2401_init   : std_logic;
		

  -- state q92
  signal reg_q92        : std_logic;
  signal reg_q92_in     : std_logic;
  signal reg_q92_init   : std_logic;
		

  -- state q960
  signal reg_q960        : std_logic;
  signal reg_q960_in     : std_logic;
  signal reg_q960_init   : std_logic;
		

  -- state q204
  signal reg_q204        : std_logic;
  signal reg_q204_in     : std_logic;
  signal reg_q204_init   : std_logic;
		

  -- state q206
  signal reg_q206        : std_logic;
  signal reg_q206_in     : std_logic;
  signal reg_q206_init   : std_logic;
		

  -- state q1566
  signal reg_q1566        : std_logic;
  signal reg_q1566_in     : std_logic;
  signal reg_q1566_init   : std_logic;
		

  -- state q1568
  signal reg_q1568        : std_logic;
  signal reg_q1568_in     : std_logic;
  signal reg_q1568_init   : std_logic;
		

  -- state q2502
  signal reg_q2502        : std_logic;
  signal reg_q2502_in     : std_logic;
  signal reg_q2502_init   : std_logic;
		

  -- state q2262
  signal reg_q2262        : std_logic;
  signal reg_q2262_in     : std_logic;
  signal reg_q2262_init   : std_logic;
		

  -- state q2264
  signal reg_q2264        : std_logic;
  signal reg_q2264_in     : std_logic;
  signal reg_q2264_init   : std_logic;
		

  -- state q430
  signal reg_q430        : std_logic;
  signal reg_q430_in     : std_logic;
  signal reg_q430_init   : std_logic;
		

  -- state q432
  signal reg_q432        : std_logic;
  signal reg_q432_in     : std_logic;
  signal reg_q432_init   : std_logic;
		

  -- state q2427
  signal reg_q2427        : std_logic;
  signal reg_q2427_in     : std_logic;
  signal reg_q2427_init   : std_logic;
		

  -- state q2371
  signal reg_q2371        : std_logic;
  signal reg_q2371_in     : std_logic;
  signal reg_q2371_init   : std_logic;
		

  -- state q1645
  signal reg_q1645        : std_logic;
  signal reg_q1645_in     : std_logic;
  signal reg_q1645_init   : std_logic;
		

  -- state q1646
  signal reg_q1646        : std_logic;
  signal reg_q1646_in     : std_logic;
  signal reg_q1646_init   : std_logic;
		

  -- state q2290
  signal reg_q2290        : std_logic;
  signal reg_q2290_in     : std_logic;
  signal reg_q2290_init   : std_logic;
		

  -- state q2292
  signal reg_q2292        : std_logic;
  signal reg_q2292_in     : std_logic;
  signal reg_q2292_init   : std_logic;
		

  -- state q2046
  signal reg_q2046        : std_logic;
  signal reg_q2046_in     : std_logic;
  signal reg_q2046_init   : std_logic;
		

  -- state q2064
  signal reg_q2064        : std_logic;
  signal reg_q2064_in     : std_logic;
  signal reg_q2064_init   : std_logic;
		

  -- state q1427
  signal reg_q1427        : std_logic;
  signal reg_q1427_in     : std_logic;
  signal reg_q1427_init   : std_logic;
		

  -- state q1429
  signal reg_q1429        : std_logic;
  signal reg_q1429_in     : std_logic;
  signal reg_q1429_init   : std_logic;
		

  -- state q2038
  signal reg_q2038        : std_logic;
  signal reg_q2038_in     : std_logic;
  signal reg_q2038_init   : std_logic;
		

  -- state q2040
  signal reg_q2040        : std_logic;
  signal reg_q2040_in     : std_logic;
  signal reg_q2040_init   : std_logic;
		

  -- state q2379
  signal reg_q2379        : std_logic;
  signal reg_q2379_in     : std_logic;
  signal reg_q2379_init   : std_logic;
		

  -- state q99
  signal reg_q99        : std_logic;
  signal reg_q99_in     : std_logic;
  signal reg_q99_init   : std_logic;
		

  -- state q1880
  signal reg_q1880        : std_logic;
  signal reg_q1880_in     : std_logic;
  signal reg_q1880_init   : std_logic;
		

  -- state q1171
  signal reg_q1171        : std_logic;
  signal reg_q1171_in     : std_logic;
  signal reg_q1171_init   : std_logic;
		

  -- state q870
  signal reg_q870        : std_logic;
  signal reg_q870_in     : std_logic;
  signal reg_q870_init   : std_logic;
		

  -- state q872
  signal reg_q872        : std_logic;
  signal reg_q872_in     : std_logic;
  signal reg_q872_init   : std_logic;
		

  -- state q1064
  signal reg_q1064        : std_logic;
  signal reg_q1064_in     : std_logic;
  signal reg_q1064_init   : std_logic;
		

  -- state q2353
  signal reg_q2353        : std_logic;
  signal reg_q2353_in     : std_logic;
  signal reg_q2353_init   : std_logic;
		

  -- state q1718
  signal reg_q1718        : std_logic;
  signal reg_q1718_in     : std_logic;
  signal reg_q1718_init   : std_logic;
		

  -- state q1828
  signal reg_q1828        : std_logic;
  signal reg_q1828_in     : std_logic;
  signal reg_q1828_init   : std_logic;
		

  -- state q70
  signal reg_q70        : std_logic;
  signal reg_q70_in     : std_logic;
  signal reg_q70_init   : std_logic;
		

  -- state q72
  signal reg_q72        : std_logic;
  signal reg_q72_in     : std_logic;
  signal reg_q72_init   : std_logic;
		

  -- state q2119
  signal reg_q2119        : std_logic;
  signal reg_q2119_in     : std_logic;
  signal reg_q2119_init   : std_logic;
		

  -- state q2121
  signal reg_q2121        : std_logic;
  signal reg_q2121_in     : std_logic;
  signal reg_q2121_init   : std_logic;
		

  -- state q1343
  signal reg_q1343        : std_logic;
  signal reg_q1343_in     : std_logic;
  signal reg_q1343_init   : std_logic;
		

  -- state q1112
  signal reg_q1112        : std_logic;
  signal reg_q1112_in     : std_logic;
  signal reg_q1112_init   : std_logic;
		

  -- state q2227
  signal reg_q2227        : std_logic;
  signal reg_q2227_in     : std_logic;
  signal reg_q2227_init   : std_logic;
		

  -- state q1037
  signal reg_q1037        : std_logic;
  signal reg_q1037_in     : std_logic;
  signal reg_q1037_init   : std_logic;
		

  -- state q1039
  signal reg_q1039        : std_logic;
  signal reg_q1039_in     : std_logic;
  signal reg_q1039_init   : std_logic;
		

  -- state q1161
  signal reg_q1161        : std_logic;
  signal reg_q1161_in     : std_logic;
  signal reg_q1161_init   : std_logic;
		

  -- state q1163
  signal reg_q1163        : std_logic;
  signal reg_q1163_in     : std_logic;
  signal reg_q1163_init   : std_logic;
		

  -- state q1399
  signal reg_q1399        : std_logic;
  signal reg_q1399_in     : std_logic;
  signal reg_q1399_init   : std_logic;
		

  -- state q1401
  signal reg_q1401        : std_logic;
  signal reg_q1401_in     : std_logic;
  signal reg_q1401_init   : std_logic;
		

  -- state q1582
  signal reg_q1582        : std_logic;
  signal reg_q1582_in     : std_logic;
  signal reg_q1582_init   : std_logic;
		

  -- state q1584
  signal reg_q1584        : std_logic;
  signal reg_q1584_in     : std_logic;
  signal reg_q1584_init   : std_logic;
		

  -- state q12
  signal reg_q12        : std_logic;
  signal reg_q12_in     : std_logic;
  signal reg_q12_init   : std_logic;
		

  -- state q143
  signal reg_q143        : std_logic;
  signal reg_q143_in     : std_logic;
  signal reg_q143_init   : std_logic;
		

  -- state q1504
  signal reg_q1504        : std_logic;
  signal reg_q1504_in     : std_logic;
  signal reg_q1504_init   : std_logic;
		

  -- state q1506
  signal reg_q1506        : std_logic;
  signal reg_q1506_in     : std_logic;
  signal reg_q1506_init   : std_logic;
		

  -- state q208
  signal reg_q208        : std_logic;
  signal reg_q208_in     : std_logic;
  signal reg_q208_init   : std_logic;
		

  -- state q210
  signal reg_q210        : std_logic;
  signal reg_q210_in     : std_logic;
  signal reg_q210_init   : std_logic;
		

  -- state q2170
  signal reg_q2170        : std_logic;
  signal reg_q2170_in     : std_logic;
  signal reg_q2170_init   : std_logic;
		

  -- state q1844
  signal reg_q1844        : std_logic;
  signal reg_q1844_in     : std_logic;
  signal reg_q1844_init   : std_logic;
		

  -- state q357
  signal reg_q357        : std_logic;
  signal reg_q357_in     : std_logic;
  signal reg_q357_init   : std_logic;
		

  -- state q359
  signal reg_q359        : std_logic;
  signal reg_q359_in     : std_logic;
  signal reg_q359_init   : std_logic;
		

  -- state q669
  signal reg_q669        : std_logic;
  signal reg_q669_in     : std_logic;
  signal reg_q669_init   : std_logic;
		

  -- state q1942
  signal reg_q1942        : std_logic;
  signal reg_q1942_in     : std_logic;
  signal reg_q1942_init   : std_logic;
		

  -- state q1944
  signal reg_q1944        : std_logic;
  signal reg_q1944_in     : std_logic;
  signal reg_q1944_init   : std_logic;
		

  -- state q1029
  signal reg_q1029        : std_logic;
  signal reg_q1029_in     : std_logic;
  signal reg_q1029_init   : std_logic;
		

  -- state q1031
  signal reg_q1031        : std_logic;
  signal reg_q1031_in     : std_logic;
  signal reg_q1031_init   : std_logic;
		

  -- state q1361
  signal reg_q1361        : std_logic;
  signal reg_q1361_in     : std_logic;
  signal reg_q1361_init   : std_logic;
		

  -- state q383
  signal reg_q383        : std_logic;
  signal reg_q383_in     : std_logic;
  signal reg_q383_init   : std_logic;
		

  -- state q642
  signal reg_q642        : std_logic;
  signal reg_q642_in     : std_logic;
  signal reg_q642_init   : std_logic;
		

  -- state q1604
  signal reg_q1604        : std_logic;
  signal reg_q1604_in     : std_logic;
  signal reg_q1604_init   : std_logic;
		

  -- state q1664
  signal reg_q1664        : std_logic;
  signal reg_q1664_in     : std_logic;
  signal reg_q1664_init   : std_logic;
		

  -- state q1932
  signal reg_q1932        : std_logic;
  signal reg_q1932_in     : std_logic;
  signal reg_q1932_init   : std_logic;
		

  -- state q2497
  signal reg_q2497        : std_logic;
  signal reg_q2497_in     : std_logic;
  signal reg_q2497_init   : std_logic;
		

  -- state q626
  signal reg_q626        : std_logic;
  signal reg_q626_in     : std_logic;
  signal reg_q626_init   : std_logic;
		

  -- state q2109
  signal reg_q2109        : std_logic;
  signal reg_q2109_in     : std_logic;
  signal reg_q2109_init   : std_logic;
		

  -- state q2111
  signal reg_q2111        : std_logic;
  signal reg_q2111_in     : std_logic;
  signal reg_q2111_init   : std_logic;
		

  -- state q2585
  signal reg_q2585        : std_logic;
  signal reg_q2585_in     : std_logic;
  signal reg_q2585_init   : std_logic;
		

  -- state q2587
  signal reg_q2587        : std_logic;
  signal reg_q2587_in     : std_logic;
  signal reg_q2587_init   : std_logic;
		

  -- state q307
  signal reg_q307        : std_logic;
  signal reg_q307_in     : std_logic;
  signal reg_q307_init   : std_logic;
		

  -- state q1533
  signal reg_q1533        : std_logic;
  signal reg_q1533_in     : std_logic;
  signal reg_q1533_init   : std_logic;
		

  -- state q2575
  signal reg_q2575        : std_logic;
  signal reg_q2575_in     : std_logic;
  signal reg_q2575_init   : std_logic;
		

  -- state q518
  signal reg_q518        : std_logic;
  signal reg_q518_in     : std_logic;
  signal reg_q518_init   : std_logic;
		

  -- state q789
  signal reg_q789        : std_logic;
  signal reg_q789_in     : std_logic;
  signal reg_q789_init   : std_logic;
		

  -- state q1734
  signal reg_q1734        : std_logic;
  signal reg_q1734_in     : std_logic;
  signal reg_q1734_init   : std_logic;
		

  -- state q1736
  signal reg_q1736        : std_logic;
  signal reg_q1736_in     : std_logic;
  signal reg_q1736_init   : std_logic;
		

  -- state q2221
  signal reg_q2221        : std_logic;
  signal reg_q2221_in     : std_logic;
  signal reg_q2221_init   : std_logic;
		

  -- state q2223
  signal reg_q2223        : std_logic;
  signal reg_q2223_in     : std_logic;
  signal reg_q2223_init   : std_logic;
		

  -- state q598
  signal reg_q598        : std_logic;
  signal reg_q598_in     : std_logic;
  signal reg_q598_init   : std_logic;
		

  -- state q600
  signal reg_q600        : std_logic;
  signal reg_q600_in     : std_logic;
  signal reg_q600_init   : std_logic;
		

  -- state q1832
  signal reg_q1832        : std_logic;
  signal reg_q1832_in     : std_logic;
  signal reg_q1832_init   : std_logic;
		

  -- state q1834
  signal reg_q1834        : std_logic;
  signal reg_q1834_in     : std_logic;
  signal reg_q1834_init   : std_logic;
		

  -- state q64
  signal reg_q64        : std_logic;
  signal reg_q64_in     : std_logic;
  signal reg_q64_init   : std_logic;
		

  -- state q66
  signal reg_q66        : std_logic;
  signal reg_q66_in     : std_logic;
  signal reg_q66_init   : std_logic;
		

  -- state q1015
  signal reg_q1015        : std_logic;
  signal reg_q1015_in     : std_logic;
  signal reg_q1015_init   : std_logic;
		

  -- state q2413
  signal reg_q2413        : std_logic;
  signal reg_q2413_in     : std_logic;
  signal reg_q2413_init   : std_logic;
		

  -- state q2385
  signal reg_q2385        : std_logic;
  signal reg_q2385_in     : std_logic;
  signal reg_q2385_init   : std_logic;
		

  -- state q2387
  signal reg_q2387        : std_logic;
  signal reg_q2387_in     : std_logic;
  signal reg_q2387_init   : std_logic;
		

  -- state q131
  signal reg_q131        : std_logic;
  signal reg_q131_in     : std_logic;
  signal reg_q131_init   : std_logic;
		

  -- state q2217
  signal reg_q2217        : std_logic;
  signal reg_q2217_in     : std_logic;
  signal reg_q2217_init   : std_logic;
		

  -- state q38
  signal reg_q38        : std_logic;
  signal reg_q38_in     : std_logic;
  signal reg_q38_init   : std_logic;
		

  -- state q40
  signal reg_q40        : std_logic;
  signal reg_q40_in     : std_logic;
  signal reg_q40_init   : std_logic;
		

  -- state q155
  signal reg_q155        : std_logic;
  signal reg_q155_in     : std_logic;
  signal reg_q155_init   : std_logic;
		

  -- state q157
  signal reg_q157        : std_logic;
  signal reg_q157_in     : std_logic;
  signal reg_q157_init   : std_logic;
		

  -- state q373
  signal reg_q373        : std_logic;
  signal reg_q373_in     : std_logic;
  signal reg_q373_init   : std_logic;
		

  -- state q36
  signal reg_q36        : std_logic;
  signal reg_q36_in     : std_logic;
  signal reg_q36_init   : std_logic;
		

  -- state q1550
  signal reg_q1550        : std_logic;
  signal reg_q1550_in     : std_logic;
  signal reg_q1550_init   : std_logic;
		

  -- state q1552
  signal reg_q1552        : std_logic;
  signal reg_q1552_in     : std_logic;
  signal reg_q1552_init   : std_logic;
		

  -- state q834
  signal reg_q834        : std_logic;
  signal reg_q834_in     : std_logic;
  signal reg_q834_init   : std_logic;
		

  -- state q923
  signal reg_q923        : std_logic;
  signal reg_q923_in     : std_logic;
  signal reg_q923_init   : std_logic;
		

  -- state q925
  signal reg_q925        : std_logic;
  signal reg_q925_in     : std_logic;
  signal reg_q925_init   : std_logic;
		

  -- state q1820
  signal reg_q1820        : std_logic;
  signal reg_q1820_in     : std_logic;
  signal reg_q1820_init   : std_logic;
		

  -- state q1143
  signal reg_q1143        : std_logic;
  signal reg_q1143_in     : std_logic;
  signal reg_q1143_init   : std_logic;
		

  -- state q1480
  signal reg_q1480        : std_logic;
  signal reg_q1480_in     : std_logic;
  signal reg_q1480_init   : std_logic;
		

  -- state q638
  signal reg_q638        : std_logic;
  signal reg_q638_in     : std_logic;
  signal reg_q638_init   : std_logic;
		

  -- state q640
  signal reg_q640        : std_logic;
  signal reg_q640_in     : std_logic;
  signal reg_q640_init   : std_logic;
		

  -- state q1179
  signal reg_q1179        : std_logic;
  signal reg_q1179_in     : std_logic;
  signal reg_q1179_init   : std_logic;
		

  -- state q1181
  signal reg_q1181        : std_logic;
  signal reg_q1181_in     : std_logic;
  signal reg_q1181_init   : std_logic;
		

  -- state q1375
  signal reg_q1375        : std_logic;
  signal reg_q1375_in     : std_logic;
  signal reg_q1375_init   : std_logic;
		

  -- state q2308
  signal reg_q2308        : std_logic;
  signal reg_q2308_in     : std_logic;
  signal reg_q2308_init   : std_logic;
		

  -- state q750
  signal reg_q750        : std_logic;
  signal reg_q750_in     : std_logic;
  signal reg_q750_init   : std_logic;
		

  -- state q1084
  signal reg_q1084        : std_logic;
  signal reg_q1084_in     : std_logic;
  signal reg_q1084_init   : std_logic;
		

  -- state q333
  signal reg_q333        : std_logic;
  signal reg_q333_in     : std_logic;
  signal reg_q333_init   : std_logic;
		

  -- state q335
  signal reg_q335        : std_logic;
  signal reg_q335_in     : std_logic;
  signal reg_q335_init   : std_logic;
		

  -- state q2288
  signal reg_q2288        : std_logic;
  signal reg_q2288_in     : std_logic;
  signal reg_q2288_init   : std_logic;
		

  -- state q6
  signal reg_q6        : std_logic;
  signal reg_q6_in     : std_logic;
  signal reg_q6_init   : std_logic;
		

  -- state q8
  signal reg_q8        : std_logic;
  signal reg_q8_in     : std_logic;
  signal reg_q8_init   : std_logic;
		

  -- state q1560
  signal reg_q1560        : std_logic;
  signal reg_q1560_in     : std_logic;
  signal reg_q1560_init   : std_logic;
		

  -- state q2266
  signal reg_q2266        : std_logic;
  signal reg_q2266_in     : std_logic;
  signal reg_q2266_init   : std_logic;
		

  -- state q1141
  signal reg_q1141        : std_logic;
  signal reg_q1141_in     : std_logic;
  signal reg_q1141_init   : std_logic;
		

  -- state q329
  signal reg_q329        : std_logic;
  signal reg_q329_in     : std_logic;
  signal reg_q329_init   : std_logic;
		

  -- state q331
  signal reg_q331        : std_logic;
  signal reg_q331_in     : std_logic;
  signal reg_q331_init   : std_logic;
		

  -- state q1488
  signal reg_q1488        : std_logic;
  signal reg_q1488_in     : std_logic;
  signal reg_q1488_init   : std_logic;
		

  -- state q1337
  signal reg_q1337        : std_logic;
  signal reg_q1337_in     : std_logic;
  signal reg_q1337_init   : std_logic;
		

  -- state q2274
  signal reg_q2274        : std_logic;
  signal reg_q2274_in     : std_logic;
  signal reg_q2274_init   : std_logic;
		

  -- state q1706
  signal reg_q1706        : std_logic;
  signal reg_q1706_in     : std_logic;
  signal reg_q1706_init   : std_logic;
		

  -- state q1708
  signal reg_q1708        : std_logic;
  signal reg_q1708_in     : std_logic;
  signal reg_q1708_init   : std_logic;
		

  -- state q1946
  signal reg_q1946        : std_logic;
  signal reg_q1946_in     : std_logic;
  signal reg_q1946_init   : std_logic;
		

  -- state q2435
  signal reg_q2435        : std_logic;
  signal reg_q2435_in     : std_logic;
  signal reg_q2435_init   : std_logic;
		

  -- state q2437
  signal reg_q2437        : std_logic;
  signal reg_q2437_in     : std_logic;
  signal reg_q2437_init   : std_logic;
		

  -- state q1464
  signal reg_q1464        : std_logic;
  signal reg_q1464_in     : std_logic;
  signal reg_q1464_init   : std_logic;
		

  -- state q1082
  signal reg_q1082        : std_logic;
  signal reg_q1082_in     : std_logic;
  signal reg_q1082_init   : std_logic;
		

  -- state q770
  signal reg_q770        : std_logic;
  signal reg_q770_in     : std_logic;
  signal reg_q770_init   : std_logic;
		

  -- state q1439
  signal reg_q1439        : std_logic;
  signal reg_q1439_in     : std_logic;
  signal reg_q1439_init   : std_logic;
		

  -- state q1744
  signal reg_q1744        : std_logic;
  signal reg_q1744_in     : std_logic;
  signal reg_q1744_init   : std_logic;
		

  -- state q1598
  signal reg_q1598        : std_logic;
  signal reg_q1598_in     : std_logic;
  signal reg_q1598_init   : std_logic;
		

  -- state q1600
  signal reg_q1600        : std_logic;
  signal reg_q1600_in     : std_logic;
  signal reg_q1600_init   : std_logic;
		

  -- state q1323
  signal reg_q1323        : std_logic;
  signal reg_q1323_in     : std_logic;
  signal reg_q1323_init   : std_logic;
		

  -- state q1325
  signal reg_q1325        : std_logic;
  signal reg_q1325_in     : std_logic;
  signal reg_q1325_init   : std_logic;
		

  -- state q1298
  signal reg_q1298        : std_logic;
  signal reg_q1298_in     : std_logic;
  signal reg_q1298_init   : std_logic;
		

  -- state q2138
  signal reg_q2138        : std_logic;
  signal reg_q2138_in     : std_logic;
  signal reg_q2138_init   : std_logic;
		

  -- state q2140
  signal reg_q2140        : std_logic;
  signal reg_q2140_in     : std_logic;
  signal reg_q2140_init   : std_logic;
		

  -- state q161
  signal reg_q161        : std_logic;
  signal reg_q161_in     : std_logic;
  signal reg_q161_init   : std_logic;
		

  -- state q163
  signal reg_q163        : std_logic;
  signal reg_q163_in     : std_logic;
  signal reg_q163_init   : std_logic;
		

  -- state q2294
  signal reg_q2294        : std_logic;
  signal reg_q2294_in     : std_logic;
  signal reg_q2294_init   : std_logic;
		

  -- state q1367
  signal reg_q1367        : std_logic;
  signal reg_q1367_in     : std_logic;
  signal reg_q1367_init   : std_logic;
		

  -- state q1748
  signal reg_q1748        : std_logic;
  signal reg_q1748_in     : std_logic;
  signal reg_q1748_init   : std_logic;
		

  -- state q2284
  signal reg_q2284        : std_logic;
  signal reg_q2284_in     : std_logic;
  signal reg_q2284_init   : std_logic;
		

  -- state q68
  signal reg_q68        : std_logic;
  signal reg_q68_in     : std_logic;
  signal reg_q68_init   : std_logic;
		

  -- state q2329
  signal reg_q2329        : std_logic;
  signal reg_q2329_in     : std_logic;
  signal reg_q2329_init   : std_logic;
		

  -- state q2331
  signal reg_q2331        : std_logic;
  signal reg_q2331_in     : std_logic;
  signal reg_q2331_init   : std_logic;
		

  -- state q984
  signal reg_q984        : std_logic;
  signal reg_q984_in     : std_logic;
  signal reg_q984_init   : std_logic;
		

  -- state q60
  signal reg_q60        : std_logic;
  signal reg_q60_in     : std_logic;
  signal reg_q60_init   : std_logic;
		

  -- state q1692
  signal reg_q1692        : std_logic;
  signal reg_q1692_in     : std_logic;
  signal reg_q1692_init   : std_logic;
		

  -- state q62
  signal reg_q62        : std_logic;
  signal reg_q62_in     : std_logic;
  signal reg_q62_init   : std_logic;
		

  -- state q395
  signal reg_q395        : std_logic;
  signal reg_q395_in     : std_logic;
  signal reg_q395_init   : std_logic;
		

  -- state q1688
  signal reg_q1688        : std_logic;
  signal reg_q1688_in     : std_logic;
  signal reg_q1688_init   : std_logic;
		

  -- state q1690
  signal reg_q1690        : std_logic;
  signal reg_q1690_in     : std_logic;
  signal reg_q1690_init   : std_logic;
		

  -- state q2134
  signal reg_q2134        : std_logic;
  signal reg_q2134_in     : std_logic;
  signal reg_q2134_init   : std_logic;
		

  -- state q2136
  signal reg_q2136        : std_logic;
  signal reg_q2136_in     : std_logic;
  signal reg_q2136_init   : std_logic;
		

  -- state q1910
  signal reg_q1910        : std_logic;
  signal reg_q1910_in     : std_logic;
  signal reg_q1910_init   : std_logic;
		

  -- state q1492
  signal reg_q1492        : std_logic;
  signal reg_q1492_in     : std_logic;
  signal reg_q1492_init   : std_logic;
		

  -- state q2117
  signal reg_q2117        : std_logic;
  signal reg_q2117_in     : std_logic;
  signal reg_q2117_init   : std_logic;
		

  -- state q2650
  signal reg_q2650        : std_logic;
  signal reg_q2650_in     : std_logic;
  signal reg_q2650_init   : std_logic;
		

  -- state q675
  signal reg_q675        : std_logic;
  signal reg_q675_in     : std_logic;
  signal reg_q675_init   : std_logic;
		

  -- state q1531
  signal reg_q1531        : std_logic;
  signal reg_q1531_in     : std_logic;
  signal reg_q1531_init   : std_logic;
		

  -- state q1900
  signal reg_q1900        : std_logic;
  signal reg_q1900_in     : std_logic;
  signal reg_q1900_init   : std_logic;
		

  -- state q1411
  signal reg_q1411        : std_logic;
  signal reg_q1411_in     : std_logic;
  signal reg_q1411_init   : std_logic;
		

  -- state q1413
  signal reg_q1413        : std_logic;
  signal reg_q1413_in     : std_logic;
  signal reg_q1413_init   : std_logic;
		

  -- state q105
  signal reg_q105        : std_logic;
  signal reg_q105_in     : std_logic;
  signal reg_q105_init   : std_logic;
		

  -- state q159
  signal reg_q159        : std_logic;
  signal reg_q159_in     : std_logic;
  signal reg_q159_init   : std_logic;
		

  -- state q2107
  signal reg_q2107        : std_logic;
  signal reg_q2107_in     : std_logic;
  signal reg_q2107_init   : std_logic;
		

  -- state q1936
  signal reg_q1936        : std_logic;
  signal reg_q1936_in     : std_logic;
  signal reg_q1936_init   : std_logic;
		

  -- state q1676
  signal reg_q1676        : std_logic;
  signal reg_q1676_in     : std_logic;
  signal reg_q1676_init   : std_logic;
		

  -- state q1678
  signal reg_q1678        : std_logic;
  signal reg_q1678_in     : std_logic;
  signal reg_q1678_init   : std_logic;
		

  -- state q1502
  signal reg_q1502        : std_logic;
  signal reg_q1502_in     : std_logic;
  signal reg_q1502_init   : std_logic;
		

  -- state q1768
  signal reg_q1768        : std_logic;
  signal reg_q1768_in     : std_logic;
  signal reg_q1768_init   : std_logic;
		

  -- state q202
  signal reg_q202        : std_logic;
  signal reg_q202_in     : std_logic;
  signal reg_q202_init   : std_logic;
		

  -- state q2510
  signal reg_q2510        : std_logic;
  signal reg_q2510_in     : std_logic;
  signal reg_q2510_init   : std_logic;
		

  -- state q2512
  signal reg_q2512        : std_logic;
  signal reg_q2512_in     : std_logic;
  signal reg_q2512_init   : std_logic;
		

  -- state q1527
  signal reg_q1527        : std_logic;
  signal reg_q1527_in     : std_logic;
  signal reg_q1527_init   : std_logic;
		

  -- state q1529
  signal reg_q1529        : std_logic;
  signal reg_q1529_in     : std_logic;
  signal reg_q1529_init   : std_logic;
		

  -- state q1496
  signal reg_q1496        : std_logic;
  signal reg_q1496_in     : std_logic;
  signal reg_q1496_init   : std_logic;
		

  -- state q2312
  signal reg_q2312        : std_logic;
  signal reg_q2312_in     : std_logic;
  signal reg_q2312_init   : std_logic;
		

  -- state q2314
  signal reg_q2314        : std_logic;
  signal reg_q2314_in     : std_logic;
  signal reg_q2314_init   : std_logic;
		

  -- state q1456
  signal reg_q1456        : std_logic;
  signal reg_q1456_in     : std_logic;
  signal reg_q1456_init   : std_logic;
		

  -- state q2692
  signal reg_q2692        : std_logic;
  signal reg_q2692_in     : std_logic;
  signal reg_q2692_init   : std_logic;
		

  -- state q2693
  signal reg_q2693        : std_logic;
  signal reg_q2693_in     : std_logic;
  signal reg_q2693_init   : std_logic;
		

  -- state q18
  signal reg_q18        : std_logic;
  signal reg_q18_in     : std_logic;
  signal reg_q18_init   : std_logic;
		

  -- state q959
  signal reg_q959        : std_logic;
  signal reg_q959_in     : std_logic;
  signal reg_q959_init   : std_logic;
		

  -- state q377
  signal reg_q377        : std_logic;
  signal reg_q377_in     : std_logic;
  signal reg_q377_init   : std_logic;
		

  -- state q2597
  signal reg_q2597        : std_logic;
  signal reg_q2597_in     : std_logic;
  signal reg_q2597_init   : std_logic;
		

  -- state q903
  signal reg_q903        : std_logic;
  signal reg_q903_in     : std_logic;
  signal reg_q903_init   : std_logic;
		

  -- state q905
  signal reg_q905        : std_logic;
  signal reg_q905_in     : std_logic;
  signal reg_q905_init   : std_logic;
		

  -- state q1415
  signal reg_q1415        : std_logic;
  signal reg_q1415_in     : std_logic;
  signal reg_q1415_init   : std_logic;
		

  -- state q1417
  signal reg_q1417        : std_logic;
  signal reg_q1417_in     : std_logic;
  signal reg_q1417_init   : std_logic;
		

  -- state q2337
  signal reg_q2337        : std_logic;
  signal reg_q2337_in     : std_logic;
  signal reg_q2337_init   : std_logic;
		

  -- state q1151
  signal reg_q1151        : std_logic;
  signal reg_q1151_in     : std_logic;
  signal reg_q1151_init   : std_logic;
		

  -- state q1153
  signal reg_q1153        : std_logic;
  signal reg_q1153_in     : std_logic;
  signal reg_q1153_init   : std_logic;
		

  -- state q2662
  signal reg_q2662        : std_logic;
  signal reg_q2662_in     : std_logic;
  signal reg_q2662_init   : std_logic;
		

  -- state q2339
  signal reg_q2339        : std_logic;
  signal reg_q2339_in     : std_logic;
  signal reg_q2339_init   : std_logic;
		

  -- state q705
  signal reg_q705        : std_logic;
  signal reg_q705_in     : std_logic;
  signal reg_q705_init   : std_logic;
		

  -- state q2345
  signal reg_q2345        : std_logic;
  signal reg_q2345_in     : std_logic;
  signal reg_q2345_init   : std_logic;
		

  -- state q1548
  signal reg_q1548        : std_logic;
  signal reg_q1548_in     : std_logic;
  signal reg_q1548_init   : std_logic;
		

  -- state q337
  signal reg_q337        : std_logic;
  signal reg_q337_in     : std_logic;
  signal reg_q337_init   : std_logic;
		

  -- state q476
  signal reg_q476        : std_logic;
  signal reg_q476_in     : std_logic;
  signal reg_q476_init   : std_logic;
		

  -- state q1478
  signal reg_q1478        : std_logic;
  signal reg_q1478_in     : std_logic;
  signal reg_q1478_init   : std_logic;
		

  -- state q2272
  signal reg_q2272        : std_logic;
  signal reg_q2272_in     : std_logic;
  signal reg_q2272_init   : std_logic;
		

  -- state q1656
  signal reg_q1656        : std_logic;
  signal reg_q1656_in     : std_logic;
  signal reg_q1656_init   : std_logic;
		

  -- state q1658
  signal reg_q1658        : std_logic;
  signal reg_q1658_in     : std_logic;
  signal reg_q1658_init   : std_logic;
		

  -- state q842
  signal reg_q842        : std_logic;
  signal reg_q842_in     : std_logic;
  signal reg_q842_init   : std_logic;
		

  -- state q1321
  signal reg_q1321        : std_logic;
  signal reg_q1321_in     : std_logic;
  signal reg_q1321_init   : std_logic;
		

  -- state q1004
  signal reg_q1004        : std_logic;
  signal reg_q1004_in     : std_logic;
  signal reg_q1004_init   : std_logic;
		

  -- state q594
  signal reg_q594        : std_logic;
  signal reg_q594_in     : std_logic;
  signal reg_q594_init   : std_logic;
		

  -- state q1051
  signal reg_q1051        : std_logic;
  signal reg_q1051_in     : std_logic;
  signal reg_q1051_init   : std_logic;
		

  -- state q2196
  signal reg_q2196        : std_logic;
  signal reg_q2196_in     : std_logic;
  signal reg_q2196_init   : std_logic;
		

  -- state q2198
  signal reg_q2198        : std_logic;
  signal reg_q2198_in     : std_logic;
  signal reg_q2198_init   : std_logic;
		

  -- state q2231
  signal reg_q2231        : std_logic;
  signal reg_q2231_in     : std_logic;
  signal reg_q2231_init   : std_logic;
		

  -- state q2455
  signal reg_q2455        : std_logic;
  signal reg_q2455_in     : std_logic;
  signal reg_q2455_init   : std_logic;
		

  -- state q2457
  signal reg_q2457        : std_logic;
  signal reg_q2457_in     : std_logic;
  signal reg_q2457_init   : std_logic;
		

  -- state q748
  signal reg_q748        : std_logic;
  signal reg_q748_in     : std_logic;
  signal reg_q748_init   : std_logic;
		

  -- state q2557
  signal reg_q2557        : std_logic;
  signal reg_q2557_in     : std_logic;
  signal reg_q2557_init   : std_logic;
		

  -- state q2559
  signal reg_q2559        : std_logic;
  signal reg_q2559_in     : std_logic;
  signal reg_q2559_init   : std_logic;
		

  -- state q2668
  signal reg_q2668        : std_logic;
  signal reg_q2668_in     : std_logic;
  signal reg_q2668_init   : std_logic;
		

  -- state q2670
  signal reg_q2670        : std_logic;
  signal reg_q2670_in     : std_logic;
  signal reg_q2670_init   : std_logic;
		

  -- state q2310
  signal reg_q2310        : std_logic;
  signal reg_q2310_in     : std_logic;
  signal reg_q2310_init   : std_logic;
		

  -- state q2150
  signal reg_q2150        : std_logic;
  signal reg_q2150_in     : std_logic;
  signal reg_q2150_init   : std_logic;
		

  -- state q466
  signal reg_q466        : std_logic;
  signal reg_q466_in     : std_logic;
  signal reg_q466_init   : std_logic;
		

  -- state q468
  signal reg_q468        : std_logic;
  signal reg_q468_in     : std_logic;
  signal reg_q468_init   : std_logic;
		

  -- state q852
  signal reg_q852        : std_logic;
  signal reg_q852_in     : std_logic;
  signal reg_q852_init   : std_logic;
		

  -- state q854
  signal reg_q854        : std_logic;
  signal reg_q854_in     : std_logic;
  signal reg_q854_init   : std_logic;
		

  -- state q415
  signal reg_q415        : std_logic;
  signal reg_q415_in     : std_logic;
  signal reg_q415_init   : std_logic;
		

  -- state q416
  signal reg_q416        : std_logic;
  signal reg_q416_in     : std_logic;
  signal reg_q416_init   : std_logic;
		

  -- state q1914
  signal reg_q1914        : std_logic;
  signal reg_q1914_in     : std_logic;
  signal reg_q1914_init   : std_logic;
		

  -- state q2439
  signal reg_q2439        : std_logic;
  signal reg_q2439_in     : std_logic;
  signal reg_q2439_init   : std_logic;
		

  -- state q1307
  signal reg_q1307        : std_logic;
  signal reg_q1307_in     : std_logic;
  signal reg_q1307_init   : std_logic;
		

  -- state q628
  signal reg_q628        : std_logic;
  signal reg_q628_in     : std_logic;
  signal reg_q628_init   : std_logic;
		

  -- state q2132
  signal reg_q2132        : std_logic;
  signal reg_q2132_in     : std_logic;
  signal reg_q2132_init   : std_logic;
		

  -- state q2459
  signal reg_q2459        : std_logic;
  signal reg_q2459_in     : std_logic;
  signal reg_q2459_init   : std_logic;
		

  -- state q1726
  signal reg_q1726        : std_logic;
  signal reg_q1726_in     : std_logic;
  signal reg_q1726_init   : std_logic;
		

  -- state q538
  signal reg_q538        : std_logic;
  signal reg_q538_in     : std_logic;
  signal reg_q538_init   : std_logic;
		

  -- state q540
  signal reg_q540        : std_logic;
  signal reg_q540_in     : std_logic;
  signal reg_q540_init   : std_logic;
		

  -- state q2583
  signal reg_q2583        : std_logic;
  signal reg_q2583_in     : std_logic;
  signal reg_q2583_init   : std_logic;
		

  -- state q588
  signal reg_q588        : std_logic;
  signal reg_q588_in     : std_logic;
  signal reg_q588_init   : std_logic;
		

  -- state q1684
  signal reg_q1684        : std_logic;
  signal reg_q1684_in     : std_logic;
  signal reg_q1684_init   : std_logic;
		

  -- state q1686
  signal reg_q1686        : std_logic;
  signal reg_q1686_in     : std_logic;
  signal reg_q1686_init   : std_logic;
		

  -- state q403
  signal reg_q403        : std_logic;
  signal reg_q403_in     : std_logic;
  signal reg_q403_init   : std_logic;
		

  -- state q405
  signal reg_q405        : std_logic;
  signal reg_q405_in     : std_logic;
  signal reg_q405_init   : std_logic;
		

  -- state q2347
  signal reg_q2347        : std_logic;
  signal reg_q2347_in     : std_logic;
  signal reg_q2347_init   : std_logic;
		

  -- state q446
  signal reg_q446        : std_logic;
  signal reg_q446_in     : std_logic;
  signal reg_q446_init   : std_logic;
		

  -- state q1014
  signal reg_q1014        : std_logic;
  signal reg_q1014_in     : std_logic;
  signal reg_q1014_init   : std_logic;
		

  -- state q570
  signal reg_q570        : std_logic;
  signal reg_q570_in     : std_logic;
  signal reg_q570_init   : std_logic;
		

  -- state q1183
  signal reg_q1183        : std_logic;
  signal reg_q1183_in     : std_logic;
  signal reg_q1183_init   : std_logic;
		

  -- state q1185
  signal reg_q1185        : std_logic;
  signal reg_q1185_in     : std_logic;
  signal reg_q1185_init   : std_logic;
		

  -- state q194
  signal reg_q194        : std_logic;
  signal reg_q194_in     : std_logic;
  signal reg_q194_init   : std_logic;
		

  -- state q196
  signal reg_q196        : std_logic;
  signal reg_q196_in     : std_logic;
  signal reg_q196_init   : std_logic;
		

  -- state q1331
  signal reg_q1331        : std_logic;
  signal reg_q1331_in     : std_logic;
  signal reg_q1331_init   : std_logic;
		

  -- state q294
  signal reg_q294        : std_logic;
  signal reg_q294_in     : std_logic;
  signal reg_q294_init   : std_logic;
		

  -- state q296
  signal reg_q296        : std_logic;
  signal reg_q296_in     : std_logic;
  signal reg_q296_init   : std_logic;
		

  -- state q1615
  signal reg_q1615        : std_logic;
  signal reg_q1615_in     : std_logic;
  signal reg_q1615_init   : std_logic;
		

  -- state q1617
  signal reg_q1617        : std_logic;
  signal reg_q1617_in     : std_logic;
  signal reg_q1617_init   : std_logic;
		

  -- state q1682
  signal reg_q1682        : std_logic;
  signal reg_q1682_in     : std_logic;
  signal reg_q1682_init   : std_logic;
		

  -- state q1892
  signal reg_q1892        : std_logic;
  signal reg_q1892_in     : std_logic;
  signal reg_q1892_init   : std_logic;
		

  -- state q502
  signal reg_q502        : std_logic;
  signal reg_q502_in     : std_logic;
  signal reg_q502_init   : std_logic;
		

  -- state q504
  signal reg_q504        : std_logic;
  signal reg_q504_in     : std_logic;
  signal reg_q504_init   : std_logic;
		

  -- state q1957
  signal reg_q1957        : std_logic;
  signal reg_q1957_in     : std_logic;
  signal reg_q1957_init   : std_logic;
		

  -- state q1959
  signal reg_q1959        : std_logic;
  signal reg_q1959_in     : std_logic;
  signal reg_q1959_init   : std_logic;
		

  -- state q1035
  signal reg_q1035        : std_logic;
  signal reg_q1035_in     : std_logic;
  signal reg_q1035_init   : std_logic;
		

  -- state q2425
  signal reg_q2425        : std_logic;
  signal reg_q2425_in     : std_logic;
  signal reg_q2425_init   : std_logic;
		

  -- state q1017
  signal reg_q1017        : std_logic;
  signal reg_q1017_in     : std_logic;
  signal reg_q1017_init   : std_logic;
		

  -- state q1019
  signal reg_q1019        : std_logic;
  signal reg_q1019_in     : std_logic;
  signal reg_q1019_init   : std_logic;
		

  -- state q361
  signal reg_q361        : std_logic;
  signal reg_q361_in     : std_logic;
  signal reg_q361_init   : std_logic;
		

  -- state q141
  signal reg_q141        : std_logic;
  signal reg_q141_in     : std_logic;
  signal reg_q141_init   : std_logic;
		

  -- state q50
  signal reg_q50        : std_logic;
  signal reg_q50_in     : std_logic;
  signal reg_q50_init   : std_logic;
		

  -- state q2522
  signal reg_q2522        : std_logic;
  signal reg_q2522_in     : std_logic;
  signal reg_q2522_init   : std_logic;
		

  -- state q586
  signal reg_q586        : std_logic;
  signal reg_q586_in     : std_logic;
  signal reg_q586_init   : std_logic;
		

  -- state q724
  signal reg_q724        : std_logic;
  signal reg_q724_in     : std_logic;
  signal reg_q724_init   : std_logic;
		

  -- state q968
  signal reg_q968        : std_logic;
  signal reg_q968_in     : std_logic;
  signal reg_q968_init   : std_logic;
		

  -- state q970
  signal reg_q970        : std_logic;
  signal reg_q970_in     : std_logic;
  signal reg_q970_init   : std_logic;
		

  -- state q1023
  signal reg_q1023        : std_logic;
  signal reg_q1023_in     : std_logic;
  signal reg_q1023_init   : std_logic;
		

  -- state q1159
  signal reg_q1159        : std_logic;
  signal reg_q1159_in     : std_logic;
  signal reg_q1159_init   : std_logic;
		

  -- state q2534
  signal reg_q2534        : std_logic;
  signal reg_q2534_in     : std_logic;
  signal reg_q2534_init   : std_logic;
		

  -- state q1169
  signal reg_q1169        : std_logic;
  signal reg_q1169_in     : std_logic;
  signal reg_q1169_init   : std_logic;
		

  -- state q349
  signal reg_q349        : std_logic;
  signal reg_q349_in     : std_logic;
  signal reg_q349_init   : std_logic;
		

  -- state q2403
  signal reg_q2403        : std_logic;
  signal reg_q2403_in     : std_logic;
  signal reg_q2403_init   : std_logic;
		

  -- state q2182
  signal reg_q2182        : std_logic;
  signal reg_q2182_in     : std_logic;
  signal reg_q2182_init   : std_logic;
		

  -- state q1033
  signal reg_q1033        : std_logic;
  signal reg_q1033_in     : std_logic;
  signal reg_q1033_init   : std_logic;
		

  -- state q2445
  signal reg_q2445        : std_logic;
  signal reg_q2445_in     : std_logic;
  signal reg_q2445_init   : std_logic;
		

  -- state q2447
  signal reg_q2447        : std_logic;
  signal reg_q2447_in     : std_logic;
  signal reg_q2447_init   : std_logic;
		

  -- state q1971
  signal reg_q1971        : std_logic;
  signal reg_q1971_in     : std_logic;
  signal reg_q1971_init   : std_logic;
		

  -- state q1973
  signal reg_q1973        : std_logic;
  signal reg_q1973_in     : std_logic;
  signal reg_q1973_init   : std_logic;
		

  -- state q2640
  signal reg_q2640        : std_logic;
  signal reg_q2640_in     : std_logic;
  signal reg_q2640_init   : std_logic;
		

  -- state q399
  signal reg_q399        : std_logic;
  signal reg_q399_in     : std_logic;
  signal reg_q399_init   : std_logic;
		

  -- state q401
  signal reg_q401        : std_logic;
  signal reg_q401_in     : std_logic;
  signal reg_q401_init   : std_logic;
		

  -- state q1447
  signal reg_q1447        : std_logic;
  signal reg_q1447_in     : std_logic;
  signal reg_q1447_init   : std_logic;
		

  -- state q1449
  signal reg_q1449        : std_logic;
  signal reg_q1449_in     : std_logic;
  signal reg_q1449_init   : std_logic;
		

  -- state q1716
  signal reg_q1716        : std_logic;
  signal reg_q1716_in     : std_logic;
  signal reg_q1716_init   : std_logic;
		

  -- state q580
  signal reg_q580        : std_logic;
  signal reg_q580_in     : std_logic;
  signal reg_q580_init   : std_logic;
		

  -- state q582
  signal reg_q582        : std_logic;
  signal reg_q582_in     : std_logic;
  signal reg_q582_init   : std_logic;
		

  -- state q1710
  signal reg_q1710        : std_logic;
  signal reg_q1710_in     : std_logic;
  signal reg_q1710_init   : std_logic;
		

  -- state q2474
  signal reg_q2474        : std_logic;
  signal reg_q2474_in     : std_logic;
  signal reg_q2474_init   : std_logic;
		

  -- state q2476
  signal reg_q2476        : std_logic;
  signal reg_q2476_in     : std_logic;
  signal reg_q2476_init   : std_logic;
		

  -- state q758
  signal reg_q758        : std_logic;
  signal reg_q758_in     : std_logic;
  signal reg_q758_init   : std_logic;
		

  -- state q760
  signal reg_q760        : std_logic;
  signal reg_q760_in     : std_logic;
  signal reg_q760_init   : std_logic;
		

  -- state q820
  signal reg_q820        : std_logic;
  signal reg_q820_in     : std_logic;
  signal reg_q820_init   : std_logic;
		

  -- state q822
  signal reg_q822        : std_logic;
  signal reg_q822_in     : std_logic;
  signal reg_q822_init   : std_logic;
		

  -- state q2010
  signal reg_q2010        : std_logic;
  signal reg_q2010_in     : std_logic;
  signal reg_q2010_init   : std_logic;
		

  -- state q2012
  signal reg_q2012        : std_logic;
  signal reg_q2012_in     : std_logic;
  signal reg_q2012_init   : std_logic;
		

  -- state q496
  signal reg_q496        : std_logic;
  signal reg_q496_in     : std_logic;
  signal reg_q496_init   : std_logic;
		

  -- state q498
  signal reg_q498        : std_logic;
  signal reg_q498_in     : std_logic;
  signal reg_q498_init   : std_logic;
		

  -- state q972
  signal reg_q972        : std_logic;
  signal reg_q972_in     : std_logic;
  signal reg_q972_init   : std_logic;
		

  -- state q730
  signal reg_q730        : std_logic;
  signal reg_q730_in     : std_logic;
  signal reg_q730_init   : std_logic;
		

  -- state q1260
  signal reg_q1260        : std_logic;
  signal reg_q1260_in     : std_logic;
  signal reg_q1260_init   : std_logic;
		

  -- state q1387
  signal reg_q1387        : std_logic;
  signal reg_q1387_in     : std_logic;
  signal reg_q1387_init   : std_logic;
		

  -- state q1389
  signal reg_q1389        : std_logic;
  signal reg_q1389_in     : std_logic;
  signal reg_q1389_init   : std_logic;
		

  -- state q1979
  signal reg_q1979        : std_logic;
  signal reg_q1979_in     : std_logic;
  signal reg_q1979_init   : std_logic;
		

  -- state q442
  signal reg_q442        : std_logic;
  signal reg_q442_in     : std_logic;
  signal reg_q442_init   : std_logic;
		

  -- state q444
  signal reg_q444        : std_logic;
  signal reg_q444_in     : std_logic;
  signal reg_q444_init   : std_logic;
		

  -- state q1092
  signal reg_q1092        : std_logic;
  signal reg_q1092_in     : std_logic;
  signal reg_q1092_init   : std_logic;
		

  -- state q1594
  signal reg_q1594        : std_logic;
  signal reg_q1594_in     : std_logic;
  signal reg_q1594_init   : std_logic;
		

  -- state q1596
  signal reg_q1596        : std_logic;
  signal reg_q1596_in     : std_logic;
  signal reg_q1596_init   : std_logic;
		

  -- state q2260
  signal reg_q2260        : std_logic;
  signal reg_q2260_in     : std_logic;
  signal reg_q2260_init   : std_logic;
		

  -- state q1956
  signal reg_q1956        : std_logic;
  signal reg_q1956_in     : std_logic;
  signal reg_q1956_init   : std_logic;
		

  -- state q1858
  signal reg_q1858        : std_logic;
  signal reg_q1858_in     : std_logic;
  signal reg_q1858_init   : std_logic;
		

  -- state q1860
  signal reg_q1860        : std_logic;
  signal reg_q1860_in     : std_logic;
  signal reg_q1860_init   : std_logic;
		

  -- state q1397
  signal reg_q1397        : std_logic;
  signal reg_q1397_in     : std_logic;
  signal reg_q1397_init   : std_logic;
		

  -- state q78
  signal reg_q78        : std_logic;
  signal reg_q78_in     : std_logic;
  signal reg_q78_init   : std_logic;
		

  -- state q229
  signal reg_q229        : std_logic;
  signal reg_q229_in     : std_logic;
  signal reg_q229_init   : std_logic;
		

  -- state q666
  signal reg_q666        : std_logic;
  signal reg_q666_in     : std_logic;
  signal reg_q666_init   : std_logic;
		

  -- state q1619
  signal reg_q1619        : std_logic;
  signal reg_q1619_in     : std_logic;
  signal reg_q1619_init   : std_logic;
		

  -- state q10
  signal reg_q10        : std_logic;
  signal reg_q10_in     : std_logic;
  signal reg_q10_init   : std_logic;
		

  -- state q1872
  signal reg_q1872        : std_logic;
  signal reg_q1872_in     : std_logic;
  signal reg_q1872_init   : std_logic;
		

  -- state q1874
  signal reg_q1874        : std_logic;
  signal reg_q1874_in     : std_logic;
  signal reg_q1874_init   : std_logic;
		

  -- state q1299
  signal reg_q1299        : std_logic;
  signal reg_q1299_in     : std_logic;
  signal reg_q1299_init   : std_logic;
		

  -- state q93
  signal reg_q93        : std_logic;
  signal reg_q93_in     : std_logic;
  signal reg_q93_init   : std_logic;
		

  -- state q95
  signal reg_q95        : std_logic;
  signal reg_q95_in     : std_logic;
  signal reg_q95_init   : std_logic;
		

  -- state q391
  signal reg_q391        : std_logic;
  signal reg_q391_in     : std_logic;
  signal reg_q391_init   : std_logic;
		

  -- state q393
  signal reg_q393        : std_logic;
  signal reg_q393_in     : std_logic;
  signal reg_q393_init   : std_logic;
		

  -- state q28
  signal reg_q28        : std_logic;
  signal reg_q28_in     : std_logic;
  signal reg_q28_init   : std_logic;
		

  -- state q1961
  signal reg_q1961        : std_logic;
  signal reg_q1961_in     : std_logic;
  signal reg_q1961_init   : std_logic;
		

  -- state q389
  signal reg_q389        : std_logic;
  signal reg_q389_in     : std_logic;
  signal reg_q389_init   : std_logic;
		

  -- state q756
  signal reg_q756        : std_logic;
  signal reg_q756_in     : std_logic;
  signal reg_q756_init   : std_logic;
		

  -- state q1760
  signal reg_q1760        : std_logic;
  signal reg_q1760_in     : std_logic;
  signal reg_q1760_init   : std_logic;
		

  -- state q838
  signal reg_q838        : std_logic;
  signal reg_q838_in     : std_logic;
  signal reg_q838_init   : std_logic;
		

  -- state q824
  signal reg_q824        : std_logic;
  signal reg_q824_in     : std_logic;
  signal reg_q824_init   : std_logic;
		

  -- state q826
  signal reg_q826        : std_logic;
  signal reg_q826_in     : std_logic;
  signal reg_q826_init   : std_logic;
		

  -- state q2680
  signal reg_q2680        : std_logic;
  signal reg_q2680_in     : std_logic;
  signal reg_q2680_init   : std_logic;
		

  -- state q2682
  signal reg_q2682        : std_logic;
  signal reg_q2682_in     : std_logic;
  signal reg_q2682_init   : std_logic;
		

  -- state q858
  signal reg_q858        : std_logic;
  signal reg_q858_in     : std_logic;
  signal reg_q858_init   : std_logic;
		

  -- state q860
  signal reg_q860        : std_logic;
  signal reg_q860_in     : std_logic;
  signal reg_q860_init   : std_logic;
		

  -- state q874
  signal reg_q874        : std_logic;
  signal reg_q874_in     : std_logic;
  signal reg_q874_init   : std_logic;
		

  -- state q2656
  signal reg_q2656        : std_logic;
  signal reg_q2656_in     : std_logic;
  signal reg_q2656_init   : std_logic;
		

  -- state q656
  signal reg_q656        : std_logic;
  signal reg_q656_in     : std_logic;
  signal reg_q656_init   : std_logic;
		

  -- state q407
  signal reg_q407        : std_logic;
  signal reg_q407_in     : std_logic;
  signal reg_q407_init   : std_logic;
		

  -- state q1466
  signal reg_q1466        : std_logic;
  signal reg_q1466_in     : std_logic;
  signal reg_q1466_init   : std_logic;
		

  -- state q2349
  signal reg_q2349        : std_logic;
  signal reg_q2349_in     : std_logic;
  signal reg_q2349_init   : std_logic;
		

  -- state q1525
  signal reg_q1525        : std_logic;
  signal reg_q1525_in     : std_logic;
  signal reg_q1525_init   : std_logic;
		

  -- state q1351
  signal reg_q1351        : std_logic;
  signal reg_q1351_in     : std_logic;
  signal reg_q1351_init   : std_logic;
		

  -- state q1353
  signal reg_q1353        : std_logic;
  signal reg_q1353_in     : std_logic;
  signal reg_q1353_init   : std_logic;
		

  -- state q1564
  signal reg_q1564        : std_logic;
  signal reg_q1564_in     : std_logic;
  signal reg_q1564_init   : std_logic;
		

  -- state q115
  signal reg_q115        : std_logic;
  signal reg_q115_in     : std_logic;
  signal reg_q115_init   : std_logic;
		

  -- state q117
  signal reg_q117        : std_logic;
  signal reg_q117_in     : std_logic;
  signal reg_q117_init   : std_logic;
		

  -- state q1123
  signal reg_q1123        : std_logic;
  signal reg_q1123_in     : std_logic;
  signal reg_q1123_init   : std_logic;
		

  -- state q550
  signal reg_q550        : std_logic;
  signal reg_q550_in     : std_logic;
  signal reg_q550_init   : std_logic;
		

  -- state q552
  signal reg_q552        : std_logic;
  signal reg_q552_in     : std_logic;
  signal reg_q552_init   : std_logic;
		

  -- state q2026
  signal reg_q2026        : std_logic;
  signal reg_q2026_in     : std_logic;
  signal reg_q2026_init   : std_logic;
		

  -- state q317
  signal reg_q317        : std_logic;
  signal reg_q317_in     : std_logic;
  signal reg_q317_init   : std_logic;
		

  -- state q319
  signal reg_q319        : std_logic;
  signal reg_q319_in     : std_logic;
  signal reg_q319_init   : std_logic;
		

  -- state q1225
  signal reg_q1225        : std_logic;
  signal reg_q1225_in     : std_logic;
  signal reg_q1225_init   : std_logic;
		

  -- state q1782
  signal reg_q1782        : std_logic;
  signal reg_q1782_in     : std_logic;
  signal reg_q1782_init   : std_logic;
		

  -- state q409
  signal reg_q409        : std_logic;
  signal reg_q409_in     : std_logic;
  signal reg_q409_init   : std_logic;
		

  -- state q411
  signal reg_q411        : std_logic;
  signal reg_q411_in     : std_logic;
  signal reg_q411_init   : std_logic;
		

  -- state q2188
  signal reg_q2188        : std_logic;
  signal reg_q2188_in     : std_logic;
  signal reg_q2188_init   : std_logic;
		

  -- state q2190
  signal reg_q2190        : std_logic;
  signal reg_q2190_in     : std_logic;
  signal reg_q2190_init   : std_logic;
		

  -- state q1177
  signal reg_q1177        : std_logic;
  signal reg_q1177_in     : std_logic;
  signal reg_q1177_init   : std_logic;
		

  -- state q2672
  signal reg_q2672        : std_logic;
  signal reg_q2672_in     : std_logic;
  signal reg_q2672_init   : std_logic;
		

  -- state q2674
  signal reg_q2674        : std_logic;
  signal reg_q2674_in     : std_logic;
  signal reg_q2674_init   : std_logic;
		

  -- state q634
  signal reg_q634        : std_logic;
  signal reg_q634_in     : std_logic;
  signal reg_q634_init   : std_logic;
		

  -- state q2125
  signal reg_q2125        : std_logic;
  signal reg_q2125_in     : std_logic;
  signal reg_q2125_init   : std_logic;
		

  -- state q2126
  signal reg_q2126        : std_logic;
  signal reg_q2126_in     : std_logic;
  signal reg_q2126_init   : std_logic;
		

  -- state q1878
  signal reg_q1878        : std_logic;
  signal reg_q1878_in     : std_logic;
  signal reg_q1878_init   : std_logic;
		

  -- state q681
  signal reg_q681        : std_logic;
  signal reg_q681_in     : std_logic;
  signal reg_q681_init   : std_logic;
		

  -- state q1836
  signal reg_q1836        : std_logic;
  signal reg_q1836_in     : std_logic;
  signal reg_q1836_init   : std_logic;
		

  -- state q1838
  signal reg_q1838        : std_logic;
  signal reg_q1838_in     : std_logic;
  signal reg_q1838_init   : std_logic;
		

  -- state q1458
  signal reg_q1458        : std_logic;
  signal reg_q1458_in     : std_logic;
  signal reg_q1458_init   : std_logic;
		

  -- state q787
  signal reg_q787        : std_logic;
  signal reg_q787_in     : std_logic;
  signal reg_q787_init   : std_logic;
		

  -- state q1391
  signal reg_q1391        : std_logic;
  signal reg_q1391_in     : std_logic;
  signal reg_q1391_init   : std_logic;
		

  -- state q1888
  signal reg_q1888        : std_logic;
  signal reg_q1888_in     : std_logic;
  signal reg_q1888_init   : std_logic;
		

  -- state q1876
  signal reg_q1876        : std_logic;
  signal reg_q1876_in     : std_logic;
  signal reg_q1876_init   : std_logic;
		

  -- state q1898
  signal reg_q1898        : std_logic;
  signal reg_q1898_in     : std_logic;
  signal reg_q1898_init   : std_logic;
		

  -- state q2176
  signal reg_q2176        : std_logic;
  signal reg_q2176_in     : std_logic;
  signal reg_q2176_init   : std_logic;
		

  -- state q434
  signal reg_q434        : std_logic;
  signal reg_q434_in     : std_logic;
  signal reg_q434_init   : std_logic;
		

  -- state q436
  signal reg_q436        : std_logic;
  signal reg_q436_in     : std_logic;
  signal reg_q436_init   : std_logic;
		

  -- state q1494
  signal reg_q1494        : std_logic;
  signal reg_q1494_in     : std_logic;
  signal reg_q1494_init   : std_logic;
		

  -- state q2146
  signal reg_q2146        : std_logic;
  signal reg_q2146_in     : std_logic;
  signal reg_q2146_init   : std_logic;
		

  -- state q1788
  signal reg_q1788        : std_logic;
  signal reg_q1788_in     : std_logic;
  signal reg_q1788_init   : std_logic;
		

  -- state q270
  signal reg_q270        : std_logic;
  signal reg_q270_in     : std_logic;
  signal reg_q270_init   : std_logic;
		

  -- state q1347
  signal reg_q1347        : std_logic;
  signal reg_q1347_in     : std_logic;
  signal reg_q1347_init   : std_logic;
		

  -- state q1349
  signal reg_q1349        : std_logic;
  signal reg_q1349_in     : std_logic;
  signal reg_q1349_init   : std_logic;
		

  -- state q1238
  signal reg_q1238        : std_logic;
  signal reg_q1238_in     : std_logic;
  signal reg_q1238_init   : std_logic;
		

  -- state q1240
  signal reg_q1240        : std_logic;
  signal reg_q1240_in     : std_logic;
  signal reg_q1240_init   : std_logic;
		

  -- state q422
  signal reg_q422        : std_logic;
  signal reg_q422_in     : std_logic;
  signal reg_q422_init   : std_logic;
		

  -- state q982
  signal reg_q982        : std_logic;
  signal reg_q982_in     : std_logic;
  signal reg_q982_init   : std_logic;
		

  -- state q1562
  signal reg_q1562        : std_logic;
  signal reg_q1562_in     : std_logic;
  signal reg_q1562_init   : std_logic;
		

  -- state q817
  signal reg_q817        : std_logic;
  signal reg_q817_in     : std_logic;
  signal reg_q817_init   : std_logic;
		

  -- state q818
  signal reg_q818        : std_logic;
  signal reg_q818_in     : std_logic;
  signal reg_q818_init   : std_logic;
		

  -- state q263
  signal reg_q263        : std_logic;
  signal reg_q263_in     : std_logic;
  signal reg_q263_init   : std_logic;
		

  -- state q264
  signal reg_q264        : std_logic;
  signal reg_q264_in     : std_logic;
  signal reg_q264_init   : std_logic;
		

  -- state q470
  signal reg_q470        : std_logic;
  signal reg_q470_in     : std_logic;
  signal reg_q470_init   : std_logic;
		

  -- state q1096
  signal reg_q1096        : std_logic;
  signal reg_q1096_in     : std_logic;
  signal reg_q1096_init   : std_logic;
		

  -- state q2441
  signal reg_q2441        : std_logic;
  signal reg_q2441_in     : std_logic;
  signal reg_q2441_init   : std_logic;
		

  -- state q2443
  signal reg_q2443        : std_logic;
  signal reg_q2443_in     : std_logic;
  signal reg_q2443_init   : std_logic;
		

  -- state q1590
  signal reg_q1590        : std_logic;
  signal reg_q1590_in     : std_logic;
  signal reg_q1590_init   : std_logic;
		

  -- state q1592
  signal reg_q1592        : std_logic;
  signal reg_q1592_in     : std_logic;
  signal reg_q1592_init   : std_logic;
		

  -- state q1774
  signal reg_q1774        : std_logic;
  signal reg_q1774_in     : std_logic;
  signal reg_q1774_init   : std_logic;
		

  -- state q1776
  signal reg_q1776        : std_logic;
  signal reg_q1776_in     : std_logic;
  signal reg_q1776_init   : std_logic;
		

  -- state q1094
  signal reg_q1094        : std_logic;
  signal reg_q1094_in     : std_logic;
  signal reg_q1094_init   : std_logic;
		

  -- state q927
  signal reg_q927        : std_logic;
  signal reg_q927_in     : std_logic;
  signal reg_q927_init   : std_logic;
		

  -- state q785
  signal reg_q785        : std_logic;
  signal reg_q785_in     : std_logic;
  signal reg_q785_init   : std_logic;
		

  -- state q2611
  signal reg_q2611        : std_logic;
  signal reg_q2611_in     : std_logic;
  signal reg_q2611_init   : std_logic;
		

  -- state q2423
  signal reg_q2423        : std_logic;
  signal reg_q2423_in     : std_logic;
  signal reg_q2423_init   : std_logic;
		

  -- state q1230
  signal reg_q1230        : std_logic;
  signal reg_q1230_in     : std_logic;
  signal reg_q1230_init   : std_logic;
		

  -- state q994
  signal reg_q994        : std_logic;
  signal reg_q994_in     : std_logic;
  signal reg_q994_init   : std_logic;
		

  -- state q996
  signal reg_q996        : std_logic;
  signal reg_q996_in     : std_logic;
  signal reg_q996_init   : std_logic;
		

  -- state q2144
  signal reg_q2144        : std_logic;
  signal reg_q2144_in     : std_logic;
  signal reg_q2144_init   : std_logic;
		

  -- state q1234
  signal reg_q1234        : std_logic;
  signal reg_q1234_in     : std_logic;
  signal reg_q1234_init   : std_logic;
		

  -- state q1236
  signal reg_q1236        : std_logic;
  signal reg_q1236_in     : std_logic;
  signal reg_q1236_init   : std_logic;
		

  -- state q2239
  signal reg_q2239        : std_logic;
  signal reg_q2239_in     : std_logic;
  signal reg_q2239_init   : std_logic;
		

  -- state q992
  signal reg_q992        : std_logic;
  signal reg_q992_in     : std_logic;
  signal reg_q992_init   : std_logic;
		

  -- state q186
  signal reg_q186        : std_logic;
  signal reg_q186_in     : std_logic;
  signal reg_q186_init   : std_logic;
		

  -- state q188
  signal reg_q188        : std_logic;
  signal reg_q188_in     : std_logic;
  signal reg_q188_init   : std_logic;
		

  -- state q1862
  signal reg_q1862        : std_logic;
  signal reg_q1862_in     : std_logic;
  signal reg_q1862_init   : std_logic;
		

  -- state q153
  signal reg_q153        : std_logic;
  signal reg_q153_in     : std_logic;
  signal reg_q153_init   : std_logic;
		

  -- state q1738
  signal reg_q1738        : std_logic;
  signal reg_q1738_in     : std_logic;
  signal reg_q1738_init   : std_logic;
		

  -- state q1740
  signal reg_q1740        : std_logic;
  signal reg_q1740_in     : std_logic;
  signal reg_q1740_init   : std_logic;
		

  -- state q282
  signal reg_q282        : std_logic;
  signal reg_q282_in     : std_logic;
  signal reg_q282_init   : std_logic;
		

  -- state q284
  signal reg_q284        : std_logic;
  signal reg_q284_in     : std_logic;
  signal reg_q284_init   : std_logic;
		

  -- state q2688
  signal reg_q2688        : std_logic;
  signal reg_q2688_in     : std_logic;
  signal reg_q2688_init   : std_logic;
		

  -- state q1280
  signal reg_q1280        : std_logic;
  signal reg_q1280_in     : std_logic;
  signal reg_q1280_init   : std_logic;
		

  -- state q1282
  signal reg_q1282        : std_logic;
  signal reg_q1282_in     : std_logic;
  signal reg_q1282_init   : std_logic;
		

  -- state q494
  signal reg_q494        : std_logic;
  signal reg_q494_in     : std_logic;
  signal reg_q494_init   : std_logic;
		

  -- state q1694
  signal reg_q1694        : std_logic;
  signal reg_q1694_in     : std_logic;
  signal reg_q1694_init   : std_logic;
		

  -- state q1431
  signal reg_q1431        : std_logic;
  signal reg_q1431_in     : std_logic;
  signal reg_q1431_init   : std_logic;
		

  -- state q2325
  signal reg_q2325        : std_logic;
  signal reg_q2325_in     : std_logic;
  signal reg_q2325_init   : std_logic;
		

  -- state q2421
  signal reg_q2421        : std_logic;
  signal reg_q2421_in     : std_logic;
  signal reg_q2421_init   : std_logic;
		

  -- state q290
  signal reg_q290        : std_logic;
  signal reg_q290_in     : std_logic;
  signal reg_q290_init   : std_logic;
		

  -- state q1570
  signal reg_q1570        : std_logic;
  signal reg_q1570_in     : std_logic;
  signal reg_q1570_init   : std_logic;
		

  -- state q1662
  signal reg_q1662        : std_logic;
  signal reg_q1662_in     : std_logic;
  signal reg_q1662_init   : std_logic;
		

  -- state q2219
  signal reg_q2219        : std_logic;
  signal reg_q2219_in     : std_logic;
  signal reg_q2219_init   : std_logic;
		

  -- state q2605
  signal reg_q2605        : std_logic;
  signal reg_q2605_in     : std_logic;
  signal reg_q2605_init   : std_logic;
		

  -- state q2607
  signal reg_q2607        : std_logic;
  signal reg_q2607_in     : std_logic;
  signal reg_q2607_init   : std_logic;
		

  -- state q32
  signal reg_q32        : std_logic;
  signal reg_q32_in     : std_logic;
  signal reg_q32_init   : std_logic;
		

  -- state q34
  signal reg_q34        : std_logic;
  signal reg_q34_in     : std_logic;
  signal reg_q34_init   : std_logic;
		

  -- state q339
  signal reg_q339        : std_logic;
  signal reg_q339_in     : std_logic;
  signal reg_q339_init   : std_logic;
		

  -- state q165
  signal reg_q165        : std_logic;
  signal reg_q165_in     : std_logic;
  signal reg_q165_init   : std_logic;
		

  -- state q1508
  signal reg_q1508        : std_logic;
  signal reg_q1508_in     : std_logic;
  signal reg_q1508_init   : std_logic;
		

  -- state q167
  signal reg_q167        : std_logic;
  signal reg_q167_in     : std_logic;
  signal reg_q167_init   : std_logic;
		

  -- state q169
  signal reg_q169        : std_logic;
  signal reg_q169_in     : std_logic;
  signal reg_q169_init   : std_logic;
		

  -- state q536
  signal reg_q536        : std_logic;
  signal reg_q536_in     : std_logic;
  signal reg_q536_init   : std_logic;
		

  -- state q1232
  signal reg_q1232        : std_logic;
  signal reg_q1232_in     : std_logic;
  signal reg_q1232_init   : std_logic;
		

  -- state q184
  signal reg_q184        : std_logic;
  signal reg_q184_in     : std_logic;
  signal reg_q184_init   : std_logic;
		

  -- state q856
  signal reg_q856        : std_logic;
  signal reg_q856_in     : std_logic;
  signal reg_q856_init   : std_logic;
		

  -- state q718
  signal reg_q718        : std_logic;
  signal reg_q718_in     : std_logic;
  signal reg_q718_init   : std_logic;
		

  -- state q1605
  signal reg_q1605        : std_logic;
  signal reg_q1605_in     : std_logic;
  signal reg_q1605_init   : std_logic;
		

  -- state q2678
  signal reg_q2678        : std_logic;
  signal reg_q2678_in     : std_logic;
  signal reg_q2678_init   : std_logic;
		

  -- state q917
  signal reg_q917        : std_logic;
  signal reg_q917_in     : std_logic;
  signal reg_q917_init   : std_logic;
		

  -- state q919
  signal reg_q919        : std_logic;
  signal reg_q919_in     : std_logic;
  signal reg_q919_init   : std_logic;
		

  -- state q2001
  signal reg_q2001        : std_logic;
  signal reg_q2001_in     : std_logic;
  signal reg_q2001_init   : std_logic;
		

  -- state q2036
  signal reg_q2036        : std_logic;
  signal reg_q2036_in     : std_logic;
  signal reg_q2036_init   : std_logic;
		

  -- state q546
  signal reg_q546        : std_logic;
  signal reg_q546_in     : std_logic;
  signal reg_q546_init   : std_logic;
		

  -- state q548
  signal reg_q548        : std_logic;
  signal reg_q548_in     : std_logic;
  signal reg_q548_init   : std_logic;
		

  -- state q2634
  signal reg_q2634        : std_logic;
  signal reg_q2634_in     : std_logic;
  signal reg_q2634_init   : std_logic;
		

  -- state q2162
  signal reg_q2162        : std_logic;
  signal reg_q2162_in     : std_logic;
  signal reg_q2162_init   : std_logic;
		

  -- state q2365
  signal reg_q2365        : std_logic;
  signal reg_q2365_in     : std_logic;
  signal reg_q2365_init   : std_logic;
		

  -- state q762
  signal reg_q762        : std_logic;
  signal reg_q762_in     : std_logic;
  signal reg_q762_init   : std_logic;
		

  -- state q764
  signal reg_q764        : std_logic;
  signal reg_q764_in     : std_logic;
  signal reg_q764_init   : std_logic;
		

  -- state q218
  signal reg_q218        : std_logic;
  signal reg_q218_in     : std_logic;
  signal reg_q218_init   : std_logic;
		

  -- state q220
  signal reg_q220        : std_logic;
  signal reg_q220_in     : std_logic;
  signal reg_q220_init   : std_logic;
		

  -- state q1357
  signal reg_q1357        : std_logic;
  signal reg_q1357_in     : std_logic;
  signal reg_q1357_init   : std_logic;
		

  -- state q1995
  signal reg_q1995        : std_logic;
  signal reg_q1995_in     : std_logic;
  signal reg_q1995_init   : std_logic;
		

  -- state q2024
  signal reg_q2024        : std_logic;
  signal reg_q2024_in     : std_logic;
  signal reg_q2024_init   : std_logic;
		

  -- state q1934
  signal reg_q1934        : std_logic;
  signal reg_q1934_in     : std_logic;
  signal reg_q1934_init   : std_logic;
		

  -- state q375
  signal reg_q375        : std_logic;
  signal reg_q375_in     : std_logic;
  signal reg_q375_init   : std_logic;
		

  -- state q2472
  signal reg_q2472        : std_logic;
  signal reg_q2472_in     : std_logic;
  signal reg_q2472_init   : std_logic;
		

  -- state q2628
  signal reg_q2628        : std_logic;
  signal reg_q2628_in     : std_logic;
  signal reg_q2628_init   : std_logic;
		

  -- state q292
  signal reg_q292        : std_logic;
  signal reg_q292_in     : std_logic;
  signal reg_q292_init   : std_logic;
		

  -- state q1702
  signal reg_q1702        : std_logic;
  signal reg_q1702_in     : std_logic;
  signal reg_q1702_init   : std_logic;
		

  -- state q1704
  signal reg_q1704        : std_logic;
  signal reg_q1704_in     : std_logic;
  signal reg_q1704_init   : std_logic;
		

  -- state q2491
  signal reg_q2491        : std_logic;
  signal reg_q2491_in     : std_logic;
  signal reg_q2491_init   : std_logic;
		

  -- state q2493
  signal reg_q2493        : std_logic;
  signal reg_q2493_in     : std_logic;
  signal reg_q2493_init   : std_logic;
		

  -- state q2451
  signal reg_q2451        : std_logic;
  signal reg_q2451_in     : std_logic;
  signal reg_q2451_init   : std_logic;
		

  -- state q2453
  signal reg_q2453        : std_logic;
  signal reg_q2453_in     : std_logic;
  signal reg_q2453_init   : std_logic;
		

  -- state q1722
  signal reg_q1722        : std_logic;
  signal reg_q1722_in     : std_logic;
  signal reg_q1722_init   : std_logic;
		

  -- state q1724
  signal reg_q1724        : std_logic;
  signal reg_q1724_in     : std_logic;
  signal reg_q1724_init   : std_logic;
		

  -- state q2101
  signal reg_q2101        : std_logic;
  signal reg_q2101_in     : std_logic;
  signal reg_q2101_init   : std_logic;
		

  -- state q1510
  signal reg_q1510        : std_logic;
  signal reg_q1510_in     : std_logic;
  signal reg_q1510_init   : std_logic;
		

  -- state q1512
  signal reg_q1512        : std_logic;
  signal reg_q1512_in     : std_logic;
  signal reg_q1512_init   : std_logic;
		

  -- state q1607
  signal reg_q1607        : std_logic;
  signal reg_q1607_in     : std_logic;
  signal reg_q1607_init   : std_logic;
		

  -- state q720
  signal reg_q720        : std_logic;
  signal reg_q720_in     : std_logic;
  signal reg_q720_init   : std_logic;
		

  -- state q722
  signal reg_q722        : std_logic;
  signal reg_q722_in     : std_logic;
  signal reg_q722_init   : std_logic;
		

  -- state q1572
  signal reg_q1572        : std_logic;
  signal reg_q1572_in     : std_logic;
  signal reg_q1572_init   : std_logic;
		

  -- state q562
  signal reg_q562        : std_logic;
  signal reg_q562_in     : std_logic;
  signal reg_q562_init   : std_logic;
		

  -- state q564
  signal reg_q564        : std_logic;
  signal reg_q564_in     : std_logic;
  signal reg_q564_init   : std_logic;
		

  -- state q1680
  signal reg_q1680        : std_logic;
  signal reg_q1680_in     : std_logic;
  signal reg_q1680_init   : std_logic;
		

  -- state q736
  signal reg_q736        : std_logic;
  signal reg_q736_in     : std_logic;
  signal reg_q736_init   : std_logic;
		

  -- state q738
  signal reg_q738        : std_logic;
  signal reg_q738_in     : std_logic;
  signal reg_q738_init   : std_logic;
		

  -- state q486
  signal reg_q486        : std_logic;
  signal reg_q486_in     : std_logic;
  signal reg_q486_init   : std_logic;
		

  -- state q488
  signal reg_q488        : std_logic;
  signal reg_q488_in     : std_logic;
  signal reg_q488_init   : std_logic;
		

  -- state q2142
  signal reg_q2142        : std_logic;
  signal reg_q2142_in     : std_logic;
  signal reg_q2142_init   : std_logic;
		

  -- state q1276
  signal reg_q1276        : std_logic;
  signal reg_q1276_in     : std_logic;
  signal reg_q1276_init   : std_logic;
		

  -- state q2237
  signal reg_q2237        : std_logic;
  signal reg_q2237_in     : std_logic;
  signal reg_q2237_init   : std_logic;
		

  -- state q1890
  signal reg_q1890        : std_logic;
  signal reg_q1890_in     : std_logic;
  signal reg_q1890_init   : std_logic;
		

  -- state q2014
  signal reg_q2014        : std_logic;
  signal reg_q2014_in     : std_logic;
  signal reg_q2014_init   : std_logic;
		

  -- state q1305
  signal reg_q1305        : std_logic;
  signal reg_q1305_in     : std_logic;
  signal reg_q1305_init   : std_logic;
		

  -- state q2549
  signal reg_q2549        : std_logic;
  signal reg_q2549_in     : std_logic;
  signal reg_q2549_init   : std_logic;
		

  -- state q2551
  signal reg_q2551        : std_logic;
  signal reg_q2551_in     : std_logic;
  signal reg_q2551_init   : std_logic;
		

  -- state q1804
  signal reg_q1804        : std_logic;
  signal reg_q1804_in     : std_logic;
  signal reg_q1804_init   : std_logic;
		

  -- state q1098
  signal reg_q1098        : std_logic;
  signal reg_q1098_in     : std_logic;
  signal reg_q1098_init   : std_logic;
		

  -- state q2200
  signal reg_q2200        : std_logic;
  signal reg_q2200_in     : std_logic;
  signal reg_q2200_init   : std_logic;
		

  -- state q182
  signal reg_q182        : std_logic;
  signal reg_q182_in     : std_logic;
  signal reg_q182_init   : std_logic;
		

  -- state q2567
  signal reg_q2567        : std_logic;
  signal reg_q2567_in     : std_logic;
  signal reg_q2567_init   : std_logic;
		

  -- state q654
  signal reg_q654        : std_logic;
  signal reg_q654_in     : std_logic;
  signal reg_q654_init   : std_logic;
		

  -- state q278
  signal reg_q278        : std_logic;
  signal reg_q278_in     : std_logic;
  signal reg_q278_init   : std_logic;
		

  -- state q280
  signal reg_q280        : std_logic;
  signal reg_q280_in     : std_logic;
  signal reg_q280_init   : std_logic;
		

  -- state q584
  signal reg_q584        : std_logic;
  signal reg_q584_in     : std_logic;
  signal reg_q584_init   : std_logic;
		

  -- state q1625
  signal reg_q1625        : std_logic;
  signal reg_q1625_in     : std_logic;
  signal reg_q1625_init   : std_logic;
		

  -- state q1627
  signal reg_q1627        : std_logic;
  signal reg_q1627_in     : std_logic;
  signal reg_q1627_init   : std_logic;
		

  -- state q1441
  signal reg_q1441        : std_logic;
  signal reg_q1441_in     : std_logic;
  signal reg_q1441_init   : std_logic;
		

  -- state q456
  signal reg_q456        : std_logic;
  signal reg_q456_in     : std_logic;
  signal reg_q456_init   : std_logic;
		

  -- state q458
  signal reg_q458        : std_logic;
  signal reg_q458_in     : std_logic;
  signal reg_q458_init   : std_logic;
		

  -- state q1732
  signal reg_q1732        : std_logic;
  signal reg_q1732_in     : std_logic;
  signal reg_q1732_init   : std_logic;
		

  -- state q4
  signal reg_q4        : std_logic;
  signal reg_q4_in     : std_logic;
  signal reg_q4_init   : std_logic;
		

  -- state q212
  signal reg_q212        : std_logic;
  signal reg_q212_in     : std_logic;
  signal reg_q212_init   : std_logic;
		

  -- state q2419
  signal reg_q2419        : std_logic;
  signal reg_q2419_in     : std_logic;
  signal reg_q2419_init   : std_logic;
		

  -- state q276
  signal reg_q276        : std_logic;
  signal reg_q276_in     : std_logic;
  signal reg_q276_init   : std_logic;
		

  -- state q345
  signal reg_q345        : std_logic;
  signal reg_q345_in     : std_logic;
  signal reg_q345_init   : std_logic;
		

  -- state q1290
  signal reg_q1290        : std_logic;
  signal reg_q1290_in     : std_logic;
  signal reg_q1290_init   : std_logic;
		

  -- state q1292
  signal reg_q1292        : std_logic;
  signal reg_q1292_in     : std_logic;
  signal reg_q1292_init   : std_logic;
		

  -- state q2078
  signal reg_q2078        : std_logic;
  signal reg_q2078_in     : std_logic;
  signal reg_q2078_init   : std_logic;
		

  -- state q2080
  signal reg_q2080        : std_logic;
  signal reg_q2080_in     : std_logic;
  signal reg_q2080_init   : std_logic;
		

  -- state q1830
  signal reg_q1830        : std_logic;
  signal reg_q1830_in     : std_logic;
  signal reg_q1830_init   : std_logic;
		

  -- state q1798
  signal reg_q1798        : std_logic;
  signal reg_q1798_in     : std_logic;
  signal reg_q1798_init   : std_logic;
		

  -- state q2020
  signal reg_q2020        : std_logic;
  signal reg_q2020_in     : std_logic;
  signal reg_q2020_init   : std_logic;
		

  -- state q2539
  signal reg_q2539        : std_logic;
  signal reg_q2539_in     : std_logic;
  signal reg_q2539_init   : std_logic;
		

  -- state q2541
  signal reg_q2541        : std_logic;
  signal reg_q2541_in     : std_logic;
  signal reg_q2541_init   : std_logic;
		

  -- state q2316
  signal reg_q2316        : std_logic;
  signal reg_q2316_in     : std_logic;
  signal reg_q2316_init   : std_logic;
		

  -- state q2318
  signal reg_q2318        : std_logic;
  signal reg_q2318_in     : std_logic;
  signal reg_q2318_init   : std_logic;
		

  -- state q931
  signal reg_q931        : std_logic;
  signal reg_q931_in     : std_logic;
  signal reg_q931_init   : std_logic;
		

  -- state q1629
  signal reg_q1629        : std_logic;
  signal reg_q1629_in     : std_logic;
  signal reg_q1629_init   : std_logic;
		

  -- state q2465
  signal reg_q2465        : std_logic;
  signal reg_q2465_in     : std_logic;
  signal reg_q2465_init   : std_logic;
		

  -- state q2056
  signal reg_q2056        : std_logic;
  signal reg_q2056_in     : std_logic;
  signal reg_q2056_init   : std_logic;
		

  -- state q2058
  signal reg_q2058        : std_logic;
  signal reg_q2058_in     : std_logic;
  signal reg_q2058_init   : std_logic;
		

  -- state q2022
  signal reg_q2022        : std_logic;
  signal reg_q2022_in     : std_logic;
  signal reg_q2022_init   : std_logic;
		

  -- state q1948
  signal reg_q1948        : std_logic;
  signal reg_q1948_in     : std_logic;
  signal reg_q1948_init   : std_logic;
		

  -- state q1950
  signal reg_q1950        : std_logic;
  signal reg_q1950_in     : std_logic;
  signal reg_q1950_init   : std_logic;
		

  -- state q2168
  signal reg_q2168        : std_logic;
  signal reg_q2168_in     : std_logic;
  signal reg_q2168_init   : std_logic;
		

  -- state q636
  signal reg_q636        : std_logic;
  signal reg_q636_in     : std_logic;
  signal reg_q636_init   : std_logic;
		

  -- state q1484
  signal reg_q1484        : std_logic;
  signal reg_q1484_in     : std_logic;
  signal reg_q1484_init   : std_logic;
		

  -- state q929
  signal reg_q929        : std_logic;
  signal reg_q929_in     : std_logic;
  signal reg_q929_init   : std_logic;
		

  -- state q460
  signal reg_q460        : std_logic;
  signal reg_q460_in     : std_logic;
  signal reg_q460_init   : std_logic;
		

  -- state q1700
  signal reg_q1700        : std_logic;
  signal reg_q1700_in     : std_logic;
  signal reg_q1700_init   : std_logic;
		

  -- state q2084
  signal reg_q2084        : std_logic;
  signal reg_q2084_in     : std_logic;
  signal reg_q2084_init   : std_logic;
		

  -- state q2086
  signal reg_q2086        : std_logic;
  signal reg_q2086_in     : std_logic;
  signal reg_q2086_init   : std_logic;
		

  -- state q1474
  signal reg_q1474        : std_logic;
  signal reg_q1474_in     : std_logic;
  signal reg_q1474_init   : std_logic;
		

  -- state q1476
  signal reg_q1476        : std_logic;
  signal reg_q1476_in     : std_logic;
  signal reg_q1476_init   : std_logic;
		

  -- state q1052
  signal reg_q1052        : std_logic;
  signal reg_q1052_in     : std_logic;
  signal reg_q1052_init   : std_logic;
		

  -- state q1054
  signal reg_q1054        : std_logic;
  signal reg_q1054_in     : std_logic;
  signal reg_q1054_init   : std_logic;
		

  -- state q2619
  signal reg_q2619        : std_logic;
  signal reg_q2619_in     : std_logic;
  signal reg_q2619_init   : std_logic;
		

  -- state q1856
  signal reg_q1856        : std_logic;
  signal reg_q1856_in     : std_logic;
  signal reg_q1856_init   : std_logic;
		

  -- state q2363
  signal reg_q2363        : std_logic;
  signal reg_q2363_in     : std_logic;
  signal reg_q2363_init   : std_logic;
		

  -- state q2327
  signal reg_q2327        : std_logic;
  signal reg_q2327_in     : std_logic;
  signal reg_q2327_init   : std_logic;
		

  -- state q222
  signal reg_q222        : std_logic;
  signal reg_q222_in     : std_logic;
  signal reg_q222_init   : std_logic;
		

  -- state q1155
  signal reg_q1155        : std_logic;
  signal reg_q1155_in     : std_logic;
  signal reg_q1155_init   : std_logic;
		

  -- state q1746
  signal reg_q1746        : std_logic;
  signal reg_q1746_in     : std_logic;
  signal reg_q1746_init   : std_logic;
		

  -- state q1262
  signal reg_q1262        : std_logic;
  signal reg_q1262_in     : std_logic;
  signal reg_q1262_init   : std_logic;
		

  -- state q2389
  signal reg_q2389        : std_logic;
  signal reg_q2389_in     : std_logic;
  signal reg_q2389_init   : std_logic;
		

  -- state q2391
  signal reg_q2391        : std_logic;
  signal reg_q2391_in     : std_logic;
  signal reg_q2391_init   : std_logic;
		

  -- state q2359
  signal reg_q2359        : std_logic;
  signal reg_q2359_in     : std_logic;
  signal reg_q2359_init   : std_logic;
		

  -- state q1952
  signal reg_q1952        : std_logic;
  signal reg_q1952_in     : std_logic;
  signal reg_q1952_init   : std_logic;
		

  -- state q2563
  signal reg_q2563        : std_logic;
  signal reg_q2563_in     : std_logic;
  signal reg_q2563_init   : std_logic;
		

  -- state q2593
  signal reg_q2593        : std_logic;
  signal reg_q2593_in     : std_logic;
  signal reg_q2593_init   : std_logic;
		

  -- state q2595
  signal reg_q2595        : std_logic;
  signal reg_q2595_in     : std_logic;
  signal reg_q2595_init   : std_logic;
		

  -- state q313
  signal reg_q313        : std_logic;
  signal reg_q313_in     : std_logic;
  signal reg_q313_init   : std_logic;
		

  -- state q315
  signal reg_q315        : std_logic;
  signal reg_q315_in     : std_logic;
  signal reg_q315_init   : std_logic;
		

  -- state q576
  signal reg_q576        : std_logic;
  signal reg_q576_in     : std_logic;
  signal reg_q576_init   : std_logic;
		

  -- state q578
  signal reg_q578        : std_logic;
  signal reg_q578_in     : std_logic;
  signal reg_q578_init   : std_logic;
		

  -- state q1472
  signal reg_q1472        : std_logic;
  signal reg_q1472_in     : std_logic;
  signal reg_q1472_init   : std_logic;
		

  -- state q2603
  signal reg_q2603        : std_logic;
  signal reg_q2603_in     : std_logic;
  signal reg_q2603_init   : std_logic;
		

  -- state q1588
  signal reg_q1588        : std_logic;
  signal reg_q1588_in     : std_logic;
  signal reg_q1588_init   : std_logic;
		

  -- state q2076
  signal reg_q2076        : std_logic;
  signal reg_q2076_in     : std_logic;
  signal reg_q2076_init   : std_logic;
		

  -- state q2206
  signal reg_q2206        : std_logic;
  signal reg_q2206_in     : std_logic;
  signal reg_q2206_init   : std_logic;
		

  -- state q2212
  signal reg_q2212        : std_logic;
  signal reg_q2212_in     : std_logic;
  signal reg_q2212_init   : std_logic;
		

  -- state q2006
  signal reg_q2006        : std_logic;
  signal reg_q2006_in     : std_logic;
  signal reg_q2006_init   : std_logic;
		

  -- state q2008
  signal reg_q2008        : std_logic;
  signal reg_q2008_in     : std_logic;
  signal reg_q2008_init   : std_logic;
		

  -- state q355
  signal reg_q355        : std_logic;
  signal reg_q355_in     : std_logic;
  signal reg_q355_init   : std_logic;
		

  -- state q1074
  signal reg_q1074        : std_logic;
  signal reg_q1074_in     : std_logic;
  signal reg_q1074_init   : std_logic;
		

  -- state q2225
  signal reg_q2225        : std_logic;
  signal reg_q2225_in     : std_logic;
  signal reg_q2225_init   : std_logic;
		

  -- state q1385
  signal reg_q1385        : std_logic;
  signal reg_q1385_in     : std_logic;
  signal reg_q1385_init   : std_logic;
		

  -- state q1119
  signal reg_q1119        : std_logic;
  signal reg_q1119_in     : std_logic;
  signal reg_q1119_init   : std_logic;
		

  -- state q274
  signal reg_q274        : std_logic;
  signal reg_q274_in     : std_logic;
  signal reg_q274_init   : std_logic;
		

  -- state q650
  signal reg_q650        : std_logic;
  signal reg_q650_in     : std_logic;
  signal reg_q650_init   : std_logic;
		

  -- state q652
  signal reg_q652        : std_logic;
  signal reg_q652_in     : std_logic;
  signal reg_q652_init   : std_logic;
		

  -- state q2609
  signal reg_q2609        : std_logic;
  signal reg_q2609_in     : std_logic;
  signal reg_q2609_init   : std_logic;
		

  -- state q1635
  signal reg_q1635        : std_logic;
  signal reg_q1635_in     : std_logic;
  signal reg_q1635_init   : std_logic;
		

  -- state q667
  signal reg_q667        : std_logic;
  signal reg_q667_in     : std_logic;
  signal reg_q667_init   : std_logic;
		

  -- state q1912
  signal reg_q1912        : std_logic;
  signal reg_q1912_in     : std_logic;
  signal reg_q1912_init   : std_logic;
		

  -- state q1514
  signal reg_q1514        : std_logic;
  signal reg_q1514_in     : std_logic;
  signal reg_q1514_init   : std_logic;
		

  -- state q1516
  signal reg_q1516        : std_logic;
  signal reg_q1516_in     : std_logic;
  signal reg_q1516_init   : std_logic;
		

  -- state q1940
  signal reg_q1940        : std_logic;
  signal reg_q1940_in     : std_logic;
  signal reg_q1940_init   : std_logic;
		

  -- state q1100
  signal reg_q1100        : std_logic;
  signal reg_q1100_in     : std_logic;
  signal reg_q1100_init   : std_logic;
		

  -- state q227
  signal reg_q227        : std_logic;
  signal reg_q227_in     : std_logic;
  signal reg_q227_init   : std_logic;
		

  -- state q506
  signal reg_q506        : std_logic;
  signal reg_q506_in     : std_logic;
  signal reg_q506_init   : std_logic;
		

  -- state q682
  signal reg_q682        : std_logic;
  signal reg_q682_in     : std_logic;
  signal reg_q682_init   : std_logic;
		

  -- state q1021
  signal reg_q1021        : std_logic;
  signal reg_q1021_in     : std_logic;
  signal reg_q1021_init   : std_logic;
		

  -- state q190
  signal reg_q190        : std_logic;
  signal reg_q190_in     : std_logic;
  signal reg_q190_init   : std_logic;
		

  -- state q192
  signal reg_q192        : std_logic;
  signal reg_q192_in     : std_logic;
  signal reg_q192_init   : std_logic;
		

  -- state q2433
  signal reg_q2433        : std_logic;
  signal reg_q2433_in     : std_logic;
  signal reg_q2433_init   : std_logic;
		

  -- state q921
  signal reg_q921        : std_logic;
  signal reg_q921_in     : std_logic;
  signal reg_q921_init   : std_logic;
		

  -- state q1278
  signal reg_q1278        : std_logic;
  signal reg_q1278_in     : std_logic;
  signal reg_q1278_init   : std_logic;
		

  -- state q214
  signal reg_q214        : std_logic;
  signal reg_q214_in     : std_logic;
  signal reg_q214_init   : std_logic;
		

  -- state q347
  signal reg_q347        : std_logic;
  signal reg_q347_in     : std_logic;
  signal reg_q347_init   : std_logic;
		

  -- state q2664
  signal reg_q2664        : std_logic;
  signal reg_q2664_in     : std_logic;
  signal reg_q2664_init   : std_logic;
		

  -- state q2676
  signal reg_q2676        : std_logic;
  signal reg_q2676_in     : std_logic;
  signal reg_q2676_init   : std_logic;
		

  -- state q2666
  signal reg_q2666        : std_logic;
  signal reg_q2666_in     : std_logic;
  signal reg_q2666_init   : std_logic;
		

  -- state q428
  signal reg_q428        : std_logic;
  signal reg_q428_in     : std_logic;
  signal reg_q428_init   : std_logic;
		

  -- state q2485
  signal reg_q2485        : std_logic;
  signal reg_q2485_in     : std_logic;
  signal reg_q2485_init   : std_logic;
		

  -- state q1637
  signal reg_q1637        : std_logic;
  signal reg_q1637_in     : std_logic;
  signal reg_q1637_init   : std_logic;
		

  -- state q2361
  signal reg_q2361        : std_logic;
  signal reg_q2361_in     : std_logic;
  signal reg_q2361_init   : std_logic;
		

  -- state q1187
  signal reg_q1187        : std_logic;
  signal reg_q1187_in     : std_logic;
  signal reg_q1187_init   : std_logic;
		

  -- state q1294
  signal reg_q1294        : std_logic;
  signal reg_q1294_in     : std_logic;
  signal reg_q1294_init   : std_logic;
		

  -- state q478
  signal reg_q478        : std_logic;
  signal reg_q478_in     : std_logic;
  signal reg_q478_init   : std_logic;
		

  -- state q1864
  signal reg_q1864        : std_logic;
  signal reg_q1864_in     : std_logic;
  signal reg_q1864_init   : std_logic;
		

  -- state q1203
  signal reg_q1203        : std_logic;
  signal reg_q1203_in     : std_logic;
  signal reg_q1203_init   : std_logic;
		

  -- state q500
  signal reg_q500        : std_logic;
  signal reg_q500_in     : std_logic;
  signal reg_q500_init   : std_logic;
		

  -- state q998
  signal reg_q998        : std_logic;
  signal reg_q998_in     : std_logic;
  signal reg_q998_init   : std_logic;
		

  -- state q171
  signal reg_q171        : std_logic;
  signal reg_q171_in     : std_logic;
  signal reg_q171_init   : std_logic;
		

  -- state q2561
  signal reg_q2561        : std_logic;
  signal reg_q2561_in     : std_logic;
  signal reg_q2561_init   : std_logic;
		

  -- state q1586
  signal reg_q1586        : std_logic;
  signal reg_q1586_in     : std_logic;
  signal reg_q1586_init   : std_logic;
		

  -- state q2320
  signal reg_q2320        : std_logic;
  signal reg_q2320_in     : std_logic;
  signal reg_q2320_init   : std_logic;
		

  -- state q42
  signal reg_q42        : std_logic;
  signal reg_q42_in     : std_logic;
  signal reg_q42_init   : std_logic;
		

  -- state q44
  signal reg_q44        : std_logic;
  signal reg_q44_in     : std_logic;
  signal reg_q44_init   : std_logic;
		

  -- state q1518
  signal reg_q1518        : std_logic;
  signal reg_q1518_in     : std_logic;
  signal reg_q1518_init   : std_logic;
		

  -- state q2626
  signal reg_q2626        : std_logic;
  signal reg_q2626_in     : std_logic;
  signal reg_q2626_init   : std_logic;
		

  -- state q2589
  signal reg_q2589        : std_logic;
  signal reg_q2589_in     : std_logic;
  signal reg_q2589_init   : std_logic;
		

  -- state q2591
  signal reg_q2591        : std_logic;
  signal reg_q2591_in     : std_logic;
  signal reg_q2591_init   : std_logic;
		

  -- state q1870
  signal reg_q1870        : std_logic;
  signal reg_q1870_in     : std_logic;
  signal reg_q1870_init   : std_logic;
		

  -- state q1157
  signal reg_q1157        : std_logic;
  signal reg_q1157_in     : std_logic;
  signal reg_q1157_init   : std_logic;
		

  -- state q776
  signal reg_q776        : std_logic;
  signal reg_q776_in     : std_logic;
  signal reg_q776_init   : std_logic;
		

  -- state q2186
  signal reg_q2186        : std_logic;
  signal reg_q2186_in     : std_logic;
  signal reg_q2186_init   : std_logic;
		

  -- state q480
  signal reg_q480        : std_logic;
  signal reg_q480_in     : std_logic;
  signal reg_q480_init   : std_logic;
		

  -- state q97
  signal reg_q97        : std_logic;
  signal reg_q97_in     : std_logic;
  signal reg_q97_init   : std_logic;
		

  -- state q1080
  signal reg_q1080        : std_logic;
  signal reg_q1080_in     : std_logic;
  signal reg_q1080_init   : std_logic;
		

  -- state q1121
  signal reg_q1121        : std_logic;
  signal reg_q1121_in     : std_logic;
  signal reg_q1121_init   : std_logic;
		

  -- state q1486
  signal reg_q1486        : std_logic;
  signal reg_q1486_in     : std_logic;
  signal reg_q1486_init   : std_logic;
		

  -- state q2082
  signal reg_q2082        : std_logic;
  signal reg_q2082_in     : std_logic;
  signal reg_q2082_init   : std_logic;
		

  -- state q492
  signal reg_q492        : std_logic;
  signal reg_q492_in     : std_logic;
  signal reg_q492_init   : std_logic;
		

  -- state q544
  signal reg_q544        : std_logic;
  signal reg_q544_in     : std_logic;
  signal reg_q544_init   : std_logic;
		

  -- state q2099
  signal reg_q2099        : std_logic;
  signal reg_q2099_in     : std_logic;
  signal reg_q2099_init   : std_logic;
		

  -- state q216
  signal reg_q216        : std_logic;
  signal reg_q216_in     : std_logic;
  signal reg_q216_init   : std_logic;
		

  -- state q1639
  signal reg_q1639        : std_logic;
  signal reg_q1639_in     : std_logic;
  signal reg_q1639_init   : std_logic;
		

  -- state q2393
  signal reg_q2393        : std_logic;
  signal reg_q2393_in     : std_logic;
  signal reg_q2393_init   : std_logic;
		

  -- state q542
  signal reg_q542        : std_logic;
  signal reg_q542_in     : std_logic;
  signal reg_q542_init   : std_logic;
		

  -- state q2504
  signal reg_q2504        : std_logic;
  signal reg_q2504_in     : std_logic;
  signal reg_q2504_init   : std_logic;
		

  -- state q1066
  signal reg_q1066        : std_logic;
  signal reg_q1066_in     : std_logic;
  signal reg_q1066_init   : std_logic;
		

  -- state q180
  signal reg_q180        : std_logic;
  signal reg_q180_in     : std_logic;
  signal reg_q180_init   : std_logic;
		

  -- state q574
  signal reg_q574        : std_logic;
  signal reg_q574_in     : std_logic;
  signal reg_q574_init   : std_logic;
		

  -- state q272
  signal reg_q272        : std_logic;
  signal reg_q272_in     : std_logic;
  signal reg_q272_init   : std_logic;
		

  -- state q1010
  signal reg_q1010        : std_logic;
  signal reg_q1010_in     : std_logic;
  signal reg_q1010_init   : std_logic;
		

  -- state q508
  signal reg_q508        : std_logic;
  signal reg_q508_in     : std_logic;
  signal reg_q508_init   : std_logic;
		

  -- state q259
  signal reg_q259        : std_logic;
  signal reg_q259_in     : std_logic;
  signal reg_q259_init   : std_logic;
		

  -- state q554
  signal reg_q554        : std_logic;
  signal reg_q554_in     : std_logic;
  signal reg_q554_init   : std_logic;
		

  -- state q2495
  signal reg_q2495        : std_logic;
  signal reg_q2495_in     : std_logic;
  signal reg_q2495_init   : std_logic;
		

  -- state q2184
  signal reg_q2184        : std_logic;
  signal reg_q2184_in     : std_logic;
  signal reg_q2184_init   : std_logic;
		

  -- state q2068
  signal reg_q2068        : std_logic;
  signal reg_q2068_in     : std_logic;
  signal reg_q2068_init   : std_logic;
		

  -- state q572
  signal reg_q572        : std_logic;
  signal reg_q572_in     : std_logic;
  signal reg_q572_init   : std_logic;
		

  -- state q2004
  signal reg_q2004        : std_logic;
  signal reg_q2004_in     : std_logic;
  signal reg_q2004_init   : std_logic;
		

  -- state q30
  signal reg_q30        : std_logic;
  signal reg_q30_in     : std_logic;
  signal reg_q30_init   : std_logic;
		

  -- state q2478
  signal reg_q2478        : std_logic;
  signal reg_q2478_in     : std_logic;
  signal reg_q2478_init   : std_logic;
		

  -- state q482
  signal reg_q482        : std_logic;
  signal reg_q482_in     : std_logic;
  signal reg_q482_init   : std_logic;
		

  -- state q484
  signal reg_q484        : std_logic;
  signal reg_q484_in     : std_logic;
  signal reg_q484_init   : std_logic;
		

  -- state q490
  signal reg_q490        : std_logic;
  signal reg_q490_in     : std_logic;
  signal reg_q490_init   : std_logic;
		

  -- state q2449
  signal reg_q2449        : std_logic;
  signal reg_q2449_in     : std_logic;
  signal reg_q2449_init   : std_logic;
		

  -- state q2547
  signal reg_q2547        : std_logic;
  signal reg_q2547_in     : std_logic;
  signal reg_q2547_init   : std_logic;
		

  -- state q953
  signal reg_q953        : std_logic;
  signal reg_q953_in     : std_logic;
  signal reg_q953_init   : std_logic;
		

  -- state q2060
  signal reg_q2060        : std_logic;
  signal reg_q2060_in     : std_logic;
  signal reg_q2060_init   : std_logic;
		

  -- state q783
  signal reg_q783        : std_logic;
  signal reg_q783_in     : std_logic;
  signal reg_q783_init   : std_logic;
		

  -- state q893
  signal reg_q893        : std_logic;
  signal reg_q893_in     : std_logic;
  signal reg_q893_init   : std_logic;
		

  -- state q886
  signal reg_q886        : std_logic;
  signal reg_q886_in     : std_logic;
  signal reg_q886_init   : std_logic;
		

  -- state q2062
  signal reg_q2062        : std_logic;
  signal reg_q2062_in     : std_logic;
  signal reg_q2062_init   : std_logic;
		

  -- state q2381
  signal reg_q2381        : std_logic;
  signal reg_q2381_in     : std_logic;
  signal reg_q2381_init   : std_logic;
		

  -- state q648
  signal reg_q648        : std_logic;
  signal reg_q648_in     : std_logic;
  signal reg_q648_init   : std_logic;
		

  -- state q811
  signal reg_q811        : std_logic;
  signal reg_q811_in     : std_logic;
  signal reg_q811_init   : std_logic;
		

  -- state q1641
  signal reg_q1641        : std_logic;
  signal reg_q1641_in     : std_logic;
  signal reg_q1641_init   : std_logic;
		

  -- state q677
  signal reg_q677        : std_logic;
  signal reg_q677_in     : std_logic;
  signal reg_q677_init   : std_logic;
		

  -- state q662
  signal reg_q662        : std_logic;
  signal reg_q662_in     : std_logic;
  signal reg_q662_init   : std_logic;
		

  -- state q846
  signal reg_q846        : std_logic;
  signal reg_q846_in     : std_logic;
  signal reg_q846_init   : std_logic;
		

  -- state q2690
  signal reg_q2690        : std_logic;
  signal reg_q2690_in     : std_logic;
  signal reg_q2690_init   : std_logic;
		

  -- state q2088
  signal reg_q2088        : std_logic;
  signal reg_q2088_in     : std_logic;
  signal reg_q2088_init   : std_logic;
		

  -- symbol decoder
  signal symb_decoder : std_logic_vector(2**DATA_WIDTH - 1 downto 0);

  -- intialization signal
  signal initialize   : std_logic;


	begin
	-- initialization
  	initialize <= INIT OR INPUT_EOF; 
	 
		symb_decoder(16#b3#) <= '1' when (INPUT = X"b3") else
                          '0';
		symb_decoder(16#a1#) <= '1' when (INPUT = X"a1") else
                          '0';
		symb_decoder(16#7f#) <= '1' when (INPUT = X"7f") else
                          '0';
		symb_decoder(16#0f#) <= '1' when (INPUT = X"0f") else
                          '0';
		symb_decoder(16#7d#) <= '1' when (INPUT = X"7d") else
                          '0';
		symb_decoder(16#15#) <= '1' when (INPUT = X"15") else
                          '0';
		symb_decoder(16#fe#) <= '1' when (INPUT = X"fe") else
                          '0';
		symb_decoder(16#1a#) <= '1' when (INPUT = X"1a") else
                          '0';
		symb_decoder(16#5a#) <= '1' when (INPUT = X"5a") else
                          '0';
		symb_decoder(16#e3#) <= '1' when (INPUT = X"e3") else
                          '0';
		symb_decoder(16#30#) <= '1' when (INPUT = X"30") else
                          '0';
		symb_decoder(16#b5#) <= '1' when (INPUT = X"b5") else
                          '0';
		symb_decoder(16#4f#) <= '1' when (INPUT = X"4f") else
                          '0';
		symb_decoder(16#55#) <= '1' when (INPUT = X"55") else
                          '0';
		symb_decoder(16#19#) <= '1' when (INPUT = X"19") else
                          '0';
		symb_decoder(16#45#) <= '1' when (INPUT = X"45") else
                          '0';
		symb_decoder(16#af#) <= '1' when (INPUT = X"af") else
                          '0';
		symb_decoder(16#ff#) <= '1' when (INPUT = X"ff") else
                          '0';
		symb_decoder(16#ea#) <= '1' when (INPUT = X"ea") else
                          '0';
		symb_decoder(16#ce#) <= '1' when (INPUT = X"ce") else
                          '0';
		symb_decoder(16#07#) <= '1' when (INPUT = X"07") else
                          '0';
		symb_decoder(16#cd#) <= '1' when (INPUT = X"cd") else
                          '0';
		symb_decoder(16#13#) <= '1' when (INPUT = X"13") else
                          '0';
		symb_decoder(16#41#) <= '1' when (INPUT = X"41") else
                          '0';
		symb_decoder(16#3d#) <= '1' when (INPUT = X"3d") else
                          '0';
		symb_decoder(16#50#) <= '1' when (INPUT = X"50") else
                          '0';
		symb_decoder(16#f3#) <= '1' when (INPUT = X"f3") else
                          '0';
		symb_decoder(16#8e#) <= '1' when (INPUT = X"8e") else
                          '0';
		symb_decoder(16#bf#) <= '1' when (INPUT = X"bf") else
                          '0';
		symb_decoder(16#ba#) <= '1' when (INPUT = X"ba") else
                          '0';
		symb_decoder(16#17#) <= '1' when (INPUT = X"17") else
                          '0';
		symb_decoder(16#08#) <= '1' when (INPUT = X"08") else
                          '0';
		symb_decoder(16#67#) <= '1' when (INPUT = X"67") else
                          '0';
		symb_decoder(16#c1#) <= '1' when (INPUT = X"c1") else
                          '0';
		symb_decoder(16#be#) <= '1' when (INPUT = X"be") else
                          '0';
		symb_decoder(16#25#) <= '1' when (INPUT = X"25") else
                          '0';
		symb_decoder(16#29#) <= '1' when (INPUT = X"29") else
                          '0';
		symb_decoder(16#28#) <= '1' when (INPUT = X"28") else
                          '0';
		symb_decoder(16#c2#) <= '1' when (INPUT = X"c2") else
                          '0';
		symb_decoder(16#a4#) <= '1' when (INPUT = X"a4") else
                          '0';
		symb_decoder(16#ab#) <= '1' when (INPUT = X"ab") else
                          '0';
		symb_decoder(16#c3#) <= '1' when (INPUT = X"c3") else
                          '0';
		symb_decoder(16#40#) <= '1' when (INPUT = X"40") else
                          '0';
		symb_decoder(16#ed#) <= '1' when (INPUT = X"ed") else
                          '0';
		symb_decoder(16#23#) <= '1' when (INPUT = X"23") else
                          '0';
		symb_decoder(16#87#) <= '1' when (INPUT = X"87") else
                          '0';
		symb_decoder(16#b8#) <= '1' when (INPUT = X"b8") else
                          '0';
		symb_decoder(16#66#) <= '1' when (INPUT = X"66") else
                          '0';
		symb_decoder(16#70#) <= '1' when (INPUT = X"70") else
                          '0';
		symb_decoder(16#20#) <= '1' when (INPUT = X"20") else
                          '0';
		symb_decoder(16#bb#) <= '1' when (INPUT = X"bb") else
                          '0';
		symb_decoder(16#10#) <= '1' when (INPUT = X"10") else
                          '0';
		symb_decoder(16#f9#) <= '1' when (INPUT = X"f9") else
                          '0';
		symb_decoder(16#ca#) <= '1' when (INPUT = X"ca") else
                          '0';
		symb_decoder(16#c5#) <= '1' when (INPUT = X"c5") else
                          '0';
		symb_decoder(16#5f#) <= '1' when (INPUT = X"5f") else
                          '0';
		symb_decoder(16#9d#) <= '1' when (INPUT = X"9d") else
                          '0';
		symb_decoder(16#3b#) <= '1' when (INPUT = X"3b") else
                          '0';
		symb_decoder(16#3c#) <= '1' when (INPUT = X"3c") else
                          '0';
		symb_decoder(16#57#) <= '1' when (INPUT = X"57") else
                          '0';
		symb_decoder(16#58#) <= '1' when (INPUT = X"58") else
                          '0';
		symb_decoder(16#0e#) <= '1' when (INPUT = X"0e") else
                          '0';
		symb_decoder(16#04#) <= '1' when (INPUT = X"04") else
                          '0';
		symb_decoder(16#84#) <= '1' when (INPUT = X"84") else
                          '0';
		symb_decoder(16#6c#) <= '1' when (INPUT = X"6c") else
                          '0';
		symb_decoder(16#61#) <= '1' when (INPUT = X"61") else
                          '0';
		symb_decoder(16#da#) <= '1' when (INPUT = X"da") else
                          '0';
		symb_decoder(16#9e#) <= '1' when (INPUT = X"9e") else
                          '0';
		symb_decoder(16#7c#) <= '1' when (INPUT = X"7c") else
                          '0';
		symb_decoder(16#44#) <= '1' when (INPUT = X"44") else
                          '0';
		symb_decoder(16#33#) <= '1' when (INPUT = X"33") else
                          '0';
		symb_decoder(16#cf#) <= '1' when (INPUT = X"cf") else
                          '0';
		symb_decoder(16#5d#) <= '1' when (INPUT = X"5d") else
                          '0';
		symb_decoder(16#6b#) <= '1' when (INPUT = X"6b") else
                          '0';
		symb_decoder(16#74#) <= '1' when (INPUT = X"74") else
                          '0';
		symb_decoder(16#f0#) <= '1' when (INPUT = X"f0") else
                          '0';
		symb_decoder(16#00#) <= '1' when (INPUT = X"00") else
                          '0';
		symb_decoder(16#fd#) <= '1' when (INPUT = X"fd") else
                          '0';
		symb_decoder(16#7e#) <= '1' when (INPUT = X"7e") else
                          '0';
		symb_decoder(16#79#) <= '1' when (INPUT = X"79") else
                          '0';
		symb_decoder(16#2f#) <= '1' when (INPUT = X"2f") else
                          '0';
		symb_decoder(16#7a#) <= '1' when (INPUT = X"7a") else
                          '0';
		symb_decoder(16#b6#) <= '1' when (INPUT = X"b6") else
                          '0';
		symb_decoder(16#8c#) <= '1' when (INPUT = X"8c") else
                          '0';
		symb_decoder(16#9a#) <= '1' when (INPUT = X"9a") else
                          '0';
		symb_decoder(16#06#) <= '1' when (INPUT = X"06") else
                          '0';
		symb_decoder(16#0b#) <= '1' when (INPUT = X"0b") else
                          '0';
		symb_decoder(16#8f#) <= '1' when (INPUT = X"8f") else
                          '0';
		symb_decoder(16#d5#) <= '1' when (INPUT = X"d5") else
                          '0';
		symb_decoder(16#99#) <= '1' when (INPUT = X"99") else
                          '0';
		symb_decoder(16#4a#) <= '1' when (INPUT = X"4a") else
                          '0';
		symb_decoder(16#5b#) <= '1' when (INPUT = X"5b") else
                          '0';
		symb_decoder(16#4b#) <= '1' when (INPUT = X"4b") else
                          '0';
		symb_decoder(16#96#) <= '1' when (INPUT = X"96") else
                          '0';
		symb_decoder(16#03#) <= '1' when (INPUT = X"03") else
                          '0';
		symb_decoder(16#dd#) <= '1' when (INPUT = X"dd") else
                          '0';
		symb_decoder(16#52#) <= '1' when (INPUT = X"52") else
                          '0';
		symb_decoder(16#94#) <= '1' when (INPUT = X"94") else
                          '0';
		symb_decoder(16#3f#) <= '1' when (INPUT = X"3f") else
                          '0';
		symb_decoder(16#65#) <= '1' when (INPUT = X"65") else
                          '0';
		symb_decoder(16#3a#) <= '1' when (INPUT = X"3a") else
                          '0';
		symb_decoder(16#d1#) <= '1' when (INPUT = X"d1") else
                          '0';
		symb_decoder(16#1e#) <= '1' when (INPUT = X"1e") else
                          '0';
		symb_decoder(16#db#) <= '1' when (INPUT = X"db") else
                          '0';
		symb_decoder(16#c6#) <= '1' when (INPUT = X"c6") else
                          '0';
		symb_decoder(16#9c#) <= '1' when (INPUT = X"9c") else
                          '0';
		symb_decoder(16#8d#) <= '1' when (INPUT = X"8d") else
                          '0';
		symb_decoder(16#a3#) <= '1' when (INPUT = X"a3") else
                          '0';
		symb_decoder(16#4c#) <= '1' when (INPUT = X"4c") else
                          '0';
		symb_decoder(16#de#) <= '1' when (INPUT = X"de") else
                          '0';
		symb_decoder(16#9b#) <= '1' when (INPUT = X"9b") else
                          '0';
		symb_decoder(16#eb#) <= '1' when (INPUT = X"eb") else
                          '0';
		symb_decoder(16#6e#) <= '1' when (INPUT = X"6e") else
                          '0';
		symb_decoder(16#62#) <= '1' when (INPUT = X"62") else
                          '0';
		symb_decoder(16#d0#) <= '1' when (INPUT = X"d0") else
                          '0';
		symb_decoder(16#ad#) <= '1' when (INPUT = X"ad") else
                          '0';
		symb_decoder(16#76#) <= '1' when (INPUT = X"76") else
                          '0';
		symb_decoder(16#aa#) <= '1' when (INPUT = X"aa") else
                          '0';
		symb_decoder(16#a6#) <= '1' when (INPUT = X"a6") else
                          '0';
		symb_decoder(16#31#) <= '1' when (INPUT = X"31") else
                          '0';
		symb_decoder(16#26#) <= '1' when (INPUT = X"26") else
                          '0';
		symb_decoder(16#f5#) <= '1' when (INPUT = X"f5") else
                          '0';
		symb_decoder(16#ef#) <= '1' when (INPUT = X"ef") else
                          '0';
		symb_decoder(16#1c#) <= '1' when (INPUT = X"1c") else
                          '0';
		symb_decoder(16#ee#) <= '1' when (INPUT = X"ee") else
                          '0';
		symb_decoder(16#73#) <= '1' when (INPUT = X"73") else
                          '0';
		symb_decoder(16#77#) <= '1' when (INPUT = X"77") else
                          '0';
		symb_decoder(16#e7#) <= '1' when (INPUT = X"e7") else
                          '0';
		symb_decoder(16#4d#) <= '1' when (INPUT = X"4d") else
                          '0';
		symb_decoder(16#38#) <= '1' when (INPUT = X"38") else
                          '0';
		symb_decoder(16#ae#) <= '1' when (INPUT = X"ae") else
                          '0';
		symb_decoder(16#02#) <= '1' when (INPUT = X"02") else
                          '0';
		symb_decoder(16#e5#) <= '1' when (INPUT = X"e5") else
                          '0';
		symb_decoder(16#ec#) <= '1' when (INPUT = X"ec") else
                          '0';
		symb_decoder(16#8b#) <= '1' when (INPUT = X"8b") else
                          '0';
		symb_decoder(16#2a#) <= '1' when (INPUT = X"2a") else
                          '0';
		symb_decoder(16#f4#) <= '1' when (INPUT = X"f4") else
                          '0';
		symb_decoder(16#0a#) <= '1' when (INPUT = X"0a") else
                          '0';
		symb_decoder(16#bd#) <= '1' when (INPUT = X"bd") else
                          '0';
		symb_decoder(16#48#) <= '1' when (INPUT = X"48") else
                          '0';
		symb_decoder(16#86#) <= '1' when (INPUT = X"86") else
                          '0';
		symb_decoder(16#39#) <= '1' when (INPUT = X"39") else
                          '0';
		symb_decoder(16#92#) <= '1' when (INPUT = X"92") else
                          '0';
		symb_decoder(16#2b#) <= '1' when (INPUT = X"2b") else
                          '0';
		symb_decoder(16#d6#) <= '1' when (INPUT = X"d6") else
                          '0';
		symb_decoder(16#05#) <= '1' when (INPUT = X"05") else
                          '0';
		symb_decoder(16#2c#) <= '1' when (INPUT = X"2c") else
                          '0';
		symb_decoder(16#97#) <= '1' when (INPUT = X"97") else
                          '0';
		symb_decoder(16#e0#) <= '1' when (INPUT = X"e0") else
                          '0';
		symb_decoder(16#82#) <= '1' when (INPUT = X"82") else
                          '0';
		symb_decoder(16#43#) <= '1' when (INPUT = X"43") else
                          '0';
		symb_decoder(16#3e#) <= '1' when (INPUT = X"3e") else
                          '0';
		symb_decoder(16#14#) <= '1' when (INPUT = X"14") else
                          '0';
		symb_decoder(16#5c#) <= '1' when (INPUT = X"5c") else
                          '0';
		symb_decoder(16#54#) <= '1' when (INPUT = X"54") else
                          '0';
		symb_decoder(16#64#) <= '1' when (INPUT = X"64") else
                          '0';
		symb_decoder(16#a2#) <= '1' when (INPUT = X"a2") else
                          '0';
		symb_decoder(16#f6#) <= '1' when (INPUT = X"f6") else
                          '0';
		symb_decoder(16#a5#) <= '1' when (INPUT = X"a5") else
                          '0';
		symb_decoder(16#c9#) <= '1' when (INPUT = X"c9") else
                          '0';
		symb_decoder(16#1b#) <= '1' when (INPUT = X"1b") else
                          '0';
		symb_decoder(16#98#) <= '1' when (INPUT = X"98") else
                          '0';
		symb_decoder(16#b1#) <= '1' when (INPUT = X"b1") else
                          '0';
		symb_decoder(16#32#) <= '1' when (INPUT = X"32") else
                          '0';
		symb_decoder(16#47#) <= '1' when (INPUT = X"47") else
                          '0';
		symb_decoder(16#1d#) <= '1' when (INPUT = X"1d") else
                          '0';
		symb_decoder(16#24#) <= '1' when (INPUT = X"24") else
                          '0';
		symb_decoder(16#d2#) <= '1' when (INPUT = X"d2") else
                          '0';
		symb_decoder(16#b7#) <= '1' when (INPUT = X"b7") else
                          '0';
		symb_decoder(16#df#) <= '1' when (INPUT = X"df") else
                          '0';
		symb_decoder(16#b4#) <= '1' when (INPUT = X"b4") else
                          '0';
		symb_decoder(16#e2#) <= '1' when (INPUT = X"e2") else
                          '0';
		symb_decoder(16#0c#) <= '1' when (INPUT = X"0c") else
                          '0';
		symb_decoder(16#81#) <= '1' when (INPUT = X"81") else
                          '0';
		symb_decoder(16#35#) <= '1' when (INPUT = X"35") else
                          '0';
		symb_decoder(16#12#) <= '1' when (INPUT = X"12") else
                          '0';
		symb_decoder(16#69#) <= '1' when (INPUT = X"69") else
                          '0';
		symb_decoder(16#59#) <= '1' when (INPUT = X"59") else
                          '0';
		symb_decoder(16#f7#) <= '1' when (INPUT = X"f7") else
                          '0';
		symb_decoder(16#fa#) <= '1' when (INPUT = X"fa") else
                          '0';
		symb_decoder(16#56#) <= '1' when (INPUT = X"56") else
                          '0';
		symb_decoder(16#75#) <= '1' when (INPUT = X"75") else
                          '0';
		symb_decoder(16#d3#) <= '1' when (INPUT = X"d3") else
                          '0';
		symb_decoder(16#cc#) <= '1' when (INPUT = X"cc") else
                          '0';
		symb_decoder(16#b0#) <= '1' when (INPUT = X"b0") else
                          '0';
		symb_decoder(16#11#) <= '1' when (INPUT = X"11") else
                          '0';
		symb_decoder(16#fb#) <= '1' when (INPUT = X"fb") else
                          '0';
		symb_decoder(16#80#) <= '1' when (INPUT = X"80") else
                          '0';
		symb_decoder(16#d7#) <= '1' when (INPUT = X"d7") else
                          '0';
		symb_decoder(16#90#) <= '1' when (INPUT = X"90") else
                          '0';
		symb_decoder(16#18#) <= '1' when (INPUT = X"18") else
                          '0';
		symb_decoder(16#34#) <= '1' when (INPUT = X"34") else
                          '0';
		symb_decoder(16#63#) <= '1' when (INPUT = X"63") else
                          '0';
		symb_decoder(16#60#) <= '1' when (INPUT = X"60") else
                          '0';
		symb_decoder(16#53#) <= '1' when (INPUT = X"53") else
                          '0';
		symb_decoder(16#16#) <= '1' when (INPUT = X"16") else
                          '0';
		symb_decoder(16#46#) <= '1' when (INPUT = X"46") else
                          '0';
		symb_decoder(16#d8#) <= '1' when (INPUT = X"d8") else
                          '0';
		symb_decoder(16#72#) <= '1' when (INPUT = X"72") else
                          '0';
		symb_decoder(16#a7#) <= '1' when (INPUT = X"a7") else
                          '0';
		symb_decoder(16#91#) <= '1' when (INPUT = X"91") else
                          '0';
		symb_decoder(16#4e#) <= '1' when (INPUT = X"4e") else
                          '0';
		symb_decoder(16#51#) <= '1' when (INPUT = X"51") else
                          '0';
		symb_decoder(16#01#) <= '1' when (INPUT = X"01") else
                          '0';
		symb_decoder(16#0d#) <= '1' when (INPUT = X"0d") else
                          '0';
		symb_decoder(16#1f#) <= '1' when (INPUT = X"1f") else
                          '0';
		symb_decoder(16#89#) <= '1' when (INPUT = X"89") else
                          '0';
		symb_decoder(16#e9#) <= '1' when (INPUT = X"e9") else
                          '0';
		symb_decoder(16#49#) <= '1' when (INPUT = X"49") else
                          '0';
		symb_decoder(16#ac#) <= '1' when (INPUT = X"ac") else
                          '0';
		symb_decoder(16#93#) <= '1' when (INPUT = X"93") else
                          '0';
		symb_decoder(16#c0#) <= '1' when (INPUT = X"c0") else
                          '0';
		symb_decoder(16#68#) <= '1' when (INPUT = X"68") else
                          '0';
		symb_decoder(16#e6#) <= '1' when (INPUT = X"e6") else
                          '0';
		symb_decoder(16#6a#) <= '1' when (INPUT = X"6a") else
                          '0';
		symb_decoder(16#c7#) <= '1' when (INPUT = X"c7") else
                          '0';
		symb_decoder(16#fc#) <= '1' when (INPUT = X"fc") else
                          '0';
		symb_decoder(16#42#) <= '1' when (INPUT = X"42") else
                          '0';
		symb_decoder(16#dc#) <= '1' when (INPUT = X"dc") else
                          '0';
		symb_decoder(16#95#) <= '1' when (INPUT = X"95") else
                          '0';
		symb_decoder(16#27#) <= '1' when (INPUT = X"27") else
                          '0';
		symb_decoder(16#b2#) <= '1' when (INPUT = X"b2") else
                          '0';
		symb_decoder(16#5e#) <= '1' when (INPUT = X"5e") else
                          '0';
		symb_decoder(16#09#) <= '1' when (INPUT = X"09") else
                          '0';
		symb_decoder(16#c4#) <= '1' when (INPUT = X"c4") else
                          '0';
		symb_decoder(16#a0#) <= '1' when (INPUT = X"a0") else
                          '0';
		symb_decoder(16#6d#) <= '1' when (INPUT = X"6d") else
                          '0';
		symb_decoder(16#83#) <= '1' when (INPUT = X"83") else
                          '0';
		symb_decoder(16#b9#) <= '1' when (INPUT = X"b9") else
                          '0';
		symb_decoder(16#88#) <= '1' when (INPUT = X"88") else
                          '0';
		symb_decoder(16#a9#) <= '1' when (INPUT = X"a9") else
                          '0';
		symb_decoder(16#cb#) <= '1' when (INPUT = X"cb") else
                          '0';
		symb_decoder(16#f8#) <= '1' when (INPUT = X"f8") else
                          '0';
		symb_decoder(16#85#) <= '1' when (INPUT = X"85") else
                          '0';
		symb_decoder(16#f2#) <= '1' when (INPUT = X"f2") else
                          '0';
		symb_decoder(16#71#) <= '1' when (INPUT = X"71") else
                          '0';
		symb_decoder(16#36#) <= '1' when (INPUT = X"36") else
                          '0';
		symb_decoder(16#21#) <= '1' when (INPUT = X"21") else
                          '0';
		symb_decoder(16#d4#) <= '1' when (INPUT = X"d4") else
                          '0';
		symb_decoder(16#2d#) <= '1' when (INPUT = X"2d") else
                          '0';
		symb_decoder(16#f1#) <= '1' when (INPUT = X"f1") else
                          '0';
		symb_decoder(16#bc#) <= '1' when (INPUT = X"bc") else
                          '0';
		symb_decoder(16#c8#) <= '1' when (INPUT = X"c8") else
                          '0';
		symb_decoder(16#37#) <= '1' when (INPUT = X"37") else
                          '0';
		symb_decoder(16#9f#) <= '1' when (INPUT = X"9f") else
                          '0';
		symb_decoder(16#a8#) <= '1' when (INPUT = X"a8") else
                          '0';
		symb_decoder(16#e8#) <= '1' when (INPUT = X"e8") else
                          '0';
		symb_decoder(16#22#) <= '1' when (INPUT = X"22") else
                          '0';
		symb_decoder(16#8a#) <= '1' when (INPUT = X"8a") else
                          '0';
		symb_decoder(16#d9#) <= '1' when (INPUT = X"d9") else
                          '0';
		symb_decoder(16#e1#) <= '1' when (INPUT = X"e1") else
                          '0';
		symb_decoder(16#2e#) <= '1' when (INPUT = X"2e") else
                          '0';
		symb_decoder(16#6f#) <= '1' when (INPUT = X"6f") else
                          '0';
		symb_decoder(16#e4#) <= '1' when (INPUT = X"e4") else
                          '0';
		symb_decoder(16#7b#) <= '1' when (INPUT = X"7b") else
                          '0';
		symb_decoder(16#78#) <= '1' when (INPUT = X"78") else
                          '0';


reg_q889_in <= (reg_q887 AND symb_decoder(16#5b#));
reg_q889_init <= '0' ;
	p_reg_q889: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q889 <= reg_q889_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q889 <= reg_q889_init;
        else
          reg_q889 <= reg_q889_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q896_in <= (reg_q889 AND symb_decoder(16#b3#)) OR
 					(reg_q889 AND symb_decoder(16#a1#)) OR
 					(reg_q889 AND symb_decoder(16#7f#)) OR
 					(reg_q889 AND symb_decoder(16#0f#)) OR
 					(reg_q889 AND symb_decoder(16#7d#)) OR
 					(reg_q889 AND symb_decoder(16#15#)) OR
 					(reg_q889 AND symb_decoder(16#fe#)) OR
 					(reg_q889 AND symb_decoder(16#1a#)) OR
 					(reg_q889 AND symb_decoder(16#5a#)) OR
 					(reg_q889 AND symb_decoder(16#e3#)) OR
 					(reg_q889 AND symb_decoder(16#30#)) OR
 					(reg_q889 AND symb_decoder(16#b5#)) OR
 					(reg_q889 AND symb_decoder(16#4f#)) OR
 					(reg_q889 AND symb_decoder(16#55#)) OR
 					(reg_q889 AND symb_decoder(16#19#)) OR
 					(reg_q889 AND symb_decoder(16#45#)) OR
 					(reg_q889 AND symb_decoder(16#af#)) OR
 					(reg_q889 AND symb_decoder(16#ff#)) OR
 					(reg_q889 AND symb_decoder(16#ea#)) OR
 					(reg_q889 AND symb_decoder(16#ce#)) OR
 					(reg_q889 AND symb_decoder(16#07#)) OR
 					(reg_q889 AND symb_decoder(16#cd#)) OR
 					(reg_q889 AND symb_decoder(16#13#)) OR
 					(reg_q889 AND symb_decoder(16#41#)) OR
 					(reg_q889 AND symb_decoder(16#3d#)) OR
 					(reg_q889 AND symb_decoder(16#50#)) OR
 					(reg_q889 AND symb_decoder(16#f3#)) OR
 					(reg_q889 AND symb_decoder(16#8e#)) OR
 					(reg_q889 AND symb_decoder(16#bf#)) OR
 					(reg_q889 AND symb_decoder(16#ba#)) OR
 					(reg_q889 AND symb_decoder(16#17#)) OR
 					(reg_q889 AND symb_decoder(16#08#)) OR
 					(reg_q889 AND symb_decoder(16#67#)) OR
 					(reg_q889 AND symb_decoder(16#c1#)) OR
 					(reg_q889 AND symb_decoder(16#be#)) OR
 					(reg_q889 AND symb_decoder(16#25#)) OR
 					(reg_q889 AND symb_decoder(16#29#)) OR
 					(reg_q889 AND symb_decoder(16#28#)) OR
 					(reg_q889 AND symb_decoder(16#c2#)) OR
 					(reg_q889 AND symb_decoder(16#a4#)) OR
 					(reg_q889 AND symb_decoder(16#ab#)) OR
 					(reg_q889 AND symb_decoder(16#c3#)) OR
 					(reg_q889 AND symb_decoder(16#40#)) OR
 					(reg_q889 AND symb_decoder(16#ed#)) OR
 					(reg_q889 AND symb_decoder(16#23#)) OR
 					(reg_q889 AND symb_decoder(16#87#)) OR
 					(reg_q889 AND symb_decoder(16#b8#)) OR
 					(reg_q889 AND symb_decoder(16#66#)) OR
 					(reg_q889 AND symb_decoder(16#70#)) OR
 					(reg_q889 AND symb_decoder(16#20#)) OR
 					(reg_q889 AND symb_decoder(16#bb#)) OR
 					(reg_q889 AND symb_decoder(16#10#)) OR
 					(reg_q889 AND symb_decoder(16#f9#)) OR
 					(reg_q889 AND symb_decoder(16#ca#)) OR
 					(reg_q889 AND symb_decoder(16#c5#)) OR
 					(reg_q889 AND symb_decoder(16#5f#)) OR
 					(reg_q889 AND symb_decoder(16#9d#)) OR
 					(reg_q889 AND symb_decoder(16#3b#)) OR
 					(reg_q889 AND symb_decoder(16#3c#)) OR
 					(reg_q889 AND symb_decoder(16#57#)) OR
 					(reg_q889 AND symb_decoder(16#58#)) OR
 					(reg_q889 AND symb_decoder(16#0e#)) OR
 					(reg_q889 AND symb_decoder(16#04#)) OR
 					(reg_q889 AND symb_decoder(16#84#)) OR
 					(reg_q889 AND symb_decoder(16#6c#)) OR
 					(reg_q889 AND symb_decoder(16#61#)) OR
 					(reg_q889 AND symb_decoder(16#da#)) OR
 					(reg_q889 AND symb_decoder(16#9e#)) OR
 					(reg_q889 AND symb_decoder(16#7c#)) OR
 					(reg_q889 AND symb_decoder(16#44#)) OR
 					(reg_q889 AND symb_decoder(16#33#)) OR
 					(reg_q889 AND symb_decoder(16#cf#)) OR
 					(reg_q889 AND symb_decoder(16#5d#)) OR
 					(reg_q889 AND symb_decoder(16#6b#)) OR
 					(reg_q889 AND symb_decoder(16#74#)) OR
 					(reg_q889 AND symb_decoder(16#f0#)) OR
 					(reg_q889 AND symb_decoder(16#00#)) OR
 					(reg_q889 AND symb_decoder(16#fd#)) OR
 					(reg_q889 AND symb_decoder(16#7e#)) OR
 					(reg_q889 AND symb_decoder(16#79#)) OR
 					(reg_q889 AND symb_decoder(16#2f#)) OR
 					(reg_q889 AND symb_decoder(16#7a#)) OR
 					(reg_q889 AND symb_decoder(16#b6#)) OR
 					(reg_q889 AND symb_decoder(16#8c#)) OR
 					(reg_q889 AND symb_decoder(16#9a#)) OR
 					(reg_q889 AND symb_decoder(16#06#)) OR
 					(reg_q889 AND symb_decoder(16#0b#)) OR
 					(reg_q889 AND symb_decoder(16#8f#)) OR
 					(reg_q889 AND symb_decoder(16#d5#)) OR
 					(reg_q889 AND symb_decoder(16#99#)) OR
 					(reg_q889 AND symb_decoder(16#4a#)) OR
 					(reg_q889 AND symb_decoder(16#5b#)) OR
 					(reg_q889 AND symb_decoder(16#4b#)) OR
 					(reg_q889 AND symb_decoder(16#96#)) OR
 					(reg_q889 AND symb_decoder(16#03#)) OR
 					(reg_q889 AND symb_decoder(16#dd#)) OR
 					(reg_q889 AND symb_decoder(16#52#)) OR
 					(reg_q889 AND symb_decoder(16#94#)) OR
 					(reg_q889 AND symb_decoder(16#3f#)) OR
 					(reg_q889 AND symb_decoder(16#65#)) OR
 					(reg_q889 AND symb_decoder(16#3a#)) OR
 					(reg_q889 AND symb_decoder(16#d1#)) OR
 					(reg_q889 AND symb_decoder(16#1e#)) OR
 					(reg_q889 AND symb_decoder(16#db#)) OR
 					(reg_q889 AND symb_decoder(16#c6#)) OR
 					(reg_q889 AND symb_decoder(16#9c#)) OR
 					(reg_q889 AND symb_decoder(16#8d#)) OR
 					(reg_q889 AND symb_decoder(16#a3#)) OR
 					(reg_q889 AND symb_decoder(16#4c#)) OR
 					(reg_q889 AND symb_decoder(16#de#)) OR
 					(reg_q889 AND symb_decoder(16#9b#)) OR
 					(reg_q889 AND symb_decoder(16#eb#)) OR
 					(reg_q889 AND symb_decoder(16#6e#)) OR
 					(reg_q889 AND symb_decoder(16#62#)) OR
 					(reg_q889 AND symb_decoder(16#d0#)) OR
 					(reg_q889 AND symb_decoder(16#ad#)) OR
 					(reg_q889 AND symb_decoder(16#76#)) OR
 					(reg_q889 AND symb_decoder(16#aa#)) OR
 					(reg_q889 AND symb_decoder(16#a6#)) OR
 					(reg_q889 AND symb_decoder(16#31#)) OR
 					(reg_q889 AND symb_decoder(16#26#)) OR
 					(reg_q889 AND symb_decoder(16#f5#)) OR
 					(reg_q889 AND symb_decoder(16#ef#)) OR
 					(reg_q889 AND symb_decoder(16#1c#)) OR
 					(reg_q889 AND symb_decoder(16#ee#)) OR
 					(reg_q889 AND symb_decoder(16#73#)) OR
 					(reg_q889 AND symb_decoder(16#77#)) OR
 					(reg_q889 AND symb_decoder(16#e7#)) OR
 					(reg_q889 AND symb_decoder(16#4d#)) OR
 					(reg_q889 AND symb_decoder(16#38#)) OR
 					(reg_q889 AND symb_decoder(16#ae#)) OR
 					(reg_q889 AND symb_decoder(16#02#)) OR
 					(reg_q889 AND symb_decoder(16#e5#)) OR
 					(reg_q889 AND symb_decoder(16#ec#)) OR
 					(reg_q889 AND symb_decoder(16#8b#)) OR
 					(reg_q889 AND symb_decoder(16#2a#)) OR
 					(reg_q889 AND symb_decoder(16#f4#)) OR
 					(reg_q889 AND symb_decoder(16#0a#)) OR
 					(reg_q889 AND symb_decoder(16#bd#)) OR
 					(reg_q889 AND symb_decoder(16#48#)) OR
 					(reg_q889 AND symb_decoder(16#86#)) OR
 					(reg_q889 AND symb_decoder(16#39#)) OR
 					(reg_q889 AND symb_decoder(16#92#)) OR
 					(reg_q889 AND symb_decoder(16#2b#)) OR
 					(reg_q889 AND symb_decoder(16#d6#)) OR
 					(reg_q889 AND symb_decoder(16#05#)) OR
 					(reg_q889 AND symb_decoder(16#2c#)) OR
 					(reg_q889 AND symb_decoder(16#97#)) OR
 					(reg_q889 AND symb_decoder(16#e0#)) OR
 					(reg_q889 AND symb_decoder(16#82#)) OR
 					(reg_q889 AND symb_decoder(16#43#)) OR
 					(reg_q889 AND symb_decoder(16#3e#)) OR
 					(reg_q889 AND symb_decoder(16#14#)) OR
 					(reg_q889 AND symb_decoder(16#5c#)) OR
 					(reg_q889 AND symb_decoder(16#54#)) OR
 					(reg_q889 AND symb_decoder(16#64#)) OR
 					(reg_q889 AND symb_decoder(16#a2#)) OR
 					(reg_q889 AND symb_decoder(16#f6#)) OR
 					(reg_q889 AND symb_decoder(16#a5#)) OR
 					(reg_q889 AND symb_decoder(16#c9#)) OR
 					(reg_q889 AND symb_decoder(16#1b#)) OR
 					(reg_q889 AND symb_decoder(16#98#)) OR
 					(reg_q889 AND symb_decoder(16#b1#)) OR
 					(reg_q889 AND symb_decoder(16#32#)) OR
 					(reg_q889 AND symb_decoder(16#47#)) OR
 					(reg_q889 AND symb_decoder(16#1d#)) OR
 					(reg_q889 AND symb_decoder(16#24#)) OR
 					(reg_q889 AND symb_decoder(16#d2#)) OR
 					(reg_q889 AND symb_decoder(16#b7#)) OR
 					(reg_q889 AND symb_decoder(16#df#)) OR
 					(reg_q889 AND symb_decoder(16#b4#)) OR
 					(reg_q889 AND symb_decoder(16#e2#)) OR
 					(reg_q889 AND symb_decoder(16#0c#)) OR
 					(reg_q889 AND symb_decoder(16#81#)) OR
 					(reg_q889 AND symb_decoder(16#35#)) OR
 					(reg_q889 AND symb_decoder(16#12#)) OR
 					(reg_q889 AND symb_decoder(16#69#)) OR
 					(reg_q889 AND symb_decoder(16#59#)) OR
 					(reg_q889 AND symb_decoder(16#f7#)) OR
 					(reg_q889 AND symb_decoder(16#fa#)) OR
 					(reg_q889 AND symb_decoder(16#56#)) OR
 					(reg_q889 AND symb_decoder(16#75#)) OR
 					(reg_q889 AND symb_decoder(16#d3#)) OR
 					(reg_q889 AND symb_decoder(16#cc#)) OR
 					(reg_q889 AND symb_decoder(16#b0#)) OR
 					(reg_q889 AND symb_decoder(16#11#)) OR
 					(reg_q889 AND symb_decoder(16#fb#)) OR
 					(reg_q889 AND symb_decoder(16#80#)) OR
 					(reg_q889 AND symb_decoder(16#d7#)) OR
 					(reg_q889 AND symb_decoder(16#90#)) OR
 					(reg_q889 AND symb_decoder(16#18#)) OR
 					(reg_q889 AND symb_decoder(16#34#)) OR
 					(reg_q889 AND symb_decoder(16#63#)) OR
 					(reg_q889 AND symb_decoder(16#60#)) OR
 					(reg_q889 AND symb_decoder(16#53#)) OR
 					(reg_q889 AND symb_decoder(16#16#)) OR
 					(reg_q889 AND symb_decoder(16#46#)) OR
 					(reg_q889 AND symb_decoder(16#d8#)) OR
 					(reg_q889 AND symb_decoder(16#72#)) OR
 					(reg_q889 AND symb_decoder(16#a7#)) OR
 					(reg_q889 AND symb_decoder(16#91#)) OR
 					(reg_q889 AND symb_decoder(16#4e#)) OR
 					(reg_q889 AND symb_decoder(16#51#)) OR
 					(reg_q889 AND symb_decoder(16#01#)) OR
 					(reg_q889 AND symb_decoder(16#0d#)) OR
 					(reg_q889 AND symb_decoder(16#1f#)) OR
 					(reg_q889 AND symb_decoder(16#89#)) OR
 					(reg_q889 AND symb_decoder(16#e9#)) OR
 					(reg_q889 AND symb_decoder(16#49#)) OR
 					(reg_q889 AND symb_decoder(16#ac#)) OR
 					(reg_q889 AND symb_decoder(16#93#)) OR
 					(reg_q889 AND symb_decoder(16#c0#)) OR
 					(reg_q889 AND symb_decoder(16#68#)) OR
 					(reg_q889 AND symb_decoder(16#e6#)) OR
 					(reg_q889 AND symb_decoder(16#6a#)) OR
 					(reg_q889 AND symb_decoder(16#c7#)) OR
 					(reg_q889 AND symb_decoder(16#fc#)) OR
 					(reg_q889 AND symb_decoder(16#42#)) OR
 					(reg_q889 AND symb_decoder(16#dc#)) OR
 					(reg_q889 AND symb_decoder(16#95#)) OR
 					(reg_q889 AND symb_decoder(16#27#)) OR
 					(reg_q889 AND symb_decoder(16#b2#)) OR
 					(reg_q889 AND symb_decoder(16#5e#)) OR
 					(reg_q889 AND symb_decoder(16#09#)) OR
 					(reg_q889 AND symb_decoder(16#c4#)) OR
 					(reg_q889 AND symb_decoder(16#a0#)) OR
 					(reg_q889 AND symb_decoder(16#6d#)) OR
 					(reg_q889 AND symb_decoder(16#83#)) OR
 					(reg_q889 AND symb_decoder(16#b9#)) OR
 					(reg_q889 AND symb_decoder(16#88#)) OR
 					(reg_q889 AND symb_decoder(16#a9#)) OR
 					(reg_q889 AND symb_decoder(16#cb#)) OR
 					(reg_q889 AND symb_decoder(16#f8#)) OR
 					(reg_q889 AND symb_decoder(16#85#)) OR
 					(reg_q889 AND symb_decoder(16#f2#)) OR
 					(reg_q889 AND symb_decoder(16#71#)) OR
 					(reg_q889 AND symb_decoder(16#36#)) OR
 					(reg_q889 AND symb_decoder(16#21#)) OR
 					(reg_q889 AND symb_decoder(16#d4#)) OR
 					(reg_q889 AND symb_decoder(16#2d#)) OR
 					(reg_q889 AND symb_decoder(16#f1#)) OR
 					(reg_q889 AND symb_decoder(16#bc#)) OR
 					(reg_q889 AND symb_decoder(16#c8#)) OR
 					(reg_q889 AND symb_decoder(16#37#)) OR
 					(reg_q889 AND symb_decoder(16#9f#)) OR
 					(reg_q889 AND symb_decoder(16#a8#)) OR
 					(reg_q889 AND symb_decoder(16#e8#)) OR
 					(reg_q889 AND symb_decoder(16#22#)) OR
 					(reg_q889 AND symb_decoder(16#8a#)) OR
 					(reg_q889 AND symb_decoder(16#d9#)) OR
 					(reg_q889 AND symb_decoder(16#e1#)) OR
 					(reg_q889 AND symb_decoder(16#2e#)) OR
 					(reg_q889 AND symb_decoder(16#6f#)) OR
 					(reg_q889 AND symb_decoder(16#e4#)) OR
 					(reg_q889 AND symb_decoder(16#7b#)) OR
 					(reg_q889 AND symb_decoder(16#78#)) OR
 					(reg_q896 AND symb_decoder(16#f9#)) OR
 					(reg_q896 AND symb_decoder(16#81#)) OR
 					(reg_q896 AND symb_decoder(16#7c#)) OR
 					(reg_q896 AND symb_decoder(16#00#)) OR
 					(reg_q896 AND symb_decoder(16#80#)) OR
 					(reg_q896 AND symb_decoder(16#8a#)) OR
 					(reg_q896 AND symb_decoder(16#4b#)) OR
 					(reg_q896 AND symb_decoder(16#95#)) OR
 					(reg_q896 AND symb_decoder(16#8d#)) OR
 					(reg_q896 AND symb_decoder(16#fb#)) OR
 					(reg_q896 AND symb_decoder(16#4e#)) OR
 					(reg_q896 AND symb_decoder(16#fd#)) OR
 					(reg_q896 AND symb_decoder(16#49#)) OR
 					(reg_q896 AND symb_decoder(16#83#)) OR
 					(reg_q896 AND symb_decoder(16#02#)) OR
 					(reg_q896 AND symb_decoder(16#ba#)) OR
 					(reg_q896 AND symb_decoder(16#31#)) OR
 					(reg_q896 AND symb_decoder(16#a6#)) OR
 					(reg_q896 AND symb_decoder(16#a9#)) OR
 					(reg_q896 AND symb_decoder(16#a4#)) OR
 					(reg_q896 AND symb_decoder(16#10#)) OR
 					(reg_q896 AND symb_decoder(16#37#)) OR
 					(reg_q896 AND symb_decoder(16#f8#)) OR
 					(reg_q896 AND symb_decoder(16#f2#)) OR
 					(reg_q896 AND symb_decoder(16#51#)) OR
 					(reg_q896 AND symb_decoder(16#52#)) OR
 					(reg_q896 AND symb_decoder(16#30#)) OR
 					(reg_q896 AND symb_decoder(16#c3#)) OR
 					(reg_q896 AND symb_decoder(16#21#)) OR
 					(reg_q896 AND symb_decoder(16#5b#)) OR
 					(reg_q896 AND symb_decoder(16#f5#)) OR
 					(reg_q896 AND symb_decoder(16#89#)) OR
 					(reg_q896 AND symb_decoder(16#0a#)) OR
 					(reg_q896 AND symb_decoder(16#e6#)) OR
 					(reg_q896 AND symb_decoder(16#ea#)) OR
 					(reg_q896 AND symb_decoder(16#3f#)) OR
 					(reg_q896 AND symb_decoder(16#0e#)) OR
 					(reg_q896 AND symb_decoder(16#22#)) OR
 					(reg_q896 AND symb_decoder(16#ac#)) OR
 					(reg_q896 AND symb_decoder(16#64#)) OR
 					(reg_q896 AND symb_decoder(16#c8#)) OR
 					(reg_q896 AND symb_decoder(16#84#)) OR
 					(reg_q896 AND symb_decoder(16#c6#)) OR
 					(reg_q896 AND symb_decoder(16#13#)) OR
 					(reg_q896 AND symb_decoder(16#2a#)) OR
 					(reg_q896 AND symb_decoder(16#fe#)) OR
 					(reg_q896 AND symb_decoder(16#bb#)) OR
 					(reg_q896 AND symb_decoder(16#d0#)) OR
 					(reg_q896 AND symb_decoder(16#dc#)) OR
 					(reg_q896 AND symb_decoder(16#05#)) OR
 					(reg_q896 AND symb_decoder(16#f3#)) OR
 					(reg_q896 AND symb_decoder(16#3a#)) OR
 					(reg_q896 AND symb_decoder(16#1d#)) OR
 					(reg_q896 AND symb_decoder(16#8e#)) OR
 					(reg_q896 AND symb_decoder(16#de#)) OR
 					(reg_q896 AND symb_decoder(16#b6#)) OR
 					(reg_q896 AND symb_decoder(16#29#)) OR
 					(reg_q896 AND symb_decoder(16#b5#)) OR
 					(reg_q896 AND symb_decoder(16#90#)) OR
 					(reg_q896 AND symb_decoder(16#71#)) OR
 					(reg_q896 AND symb_decoder(16#b4#)) OR
 					(reg_q896 AND symb_decoder(16#ad#)) OR
 					(reg_q896 AND symb_decoder(16#85#)) OR
 					(reg_q896 AND symb_decoder(16#27#)) OR
 					(reg_q896 AND symb_decoder(16#e0#)) OR
 					(reg_q896 AND symb_decoder(16#69#)) OR
 					(reg_q896 AND symb_decoder(16#fc#)) OR
 					(reg_q896 AND symb_decoder(16#d8#)) OR
 					(reg_q896 AND symb_decoder(16#53#)) OR
 					(reg_q896 AND symb_decoder(16#0c#)) OR
 					(reg_q896 AND symb_decoder(16#3c#)) OR
 					(reg_q896 AND symb_decoder(16#af#)) OR
 					(reg_q896 AND symb_decoder(16#2c#)) OR
 					(reg_q896 AND symb_decoder(16#25#)) OR
 					(reg_q896 AND symb_decoder(16#f7#)) OR
 					(reg_q896 AND symb_decoder(16#61#)) OR
 					(reg_q896 AND symb_decoder(16#9e#)) OR
 					(reg_q896 AND symb_decoder(16#2b#)) OR
 					(reg_q896 AND symb_decoder(16#09#)) OR
 					(reg_q896 AND symb_decoder(16#56#)) OR
 					(reg_q896 AND symb_decoder(16#07#)) OR
 					(reg_q896 AND symb_decoder(16#d2#)) OR
 					(reg_q896 AND symb_decoder(16#a3#)) OR
 					(reg_q896 AND symb_decoder(16#46#)) OR
 					(reg_q896 AND symb_decoder(16#41#)) OR
 					(reg_q896 AND symb_decoder(16#58#)) OR
 					(reg_q896 AND symb_decoder(16#5c#)) OR
 					(reg_q896 AND symb_decoder(16#4f#)) OR
 					(reg_q896 AND symb_decoder(16#39#)) OR
 					(reg_q896 AND symb_decoder(16#94#)) OR
 					(reg_q896 AND symb_decoder(16#19#)) OR
 					(reg_q896 AND symb_decoder(16#96#)) OR
 					(reg_q896 AND symb_decoder(16#ab#)) OR
 					(reg_q896 AND symb_decoder(16#2e#)) OR
 					(reg_q896 AND symb_decoder(16#df#)) OR
 					(reg_q896 AND symb_decoder(16#a7#)) OR
 					(reg_q896 AND symb_decoder(16#cd#)) OR
 					(reg_q896 AND symb_decoder(16#5d#)) OR
 					(reg_q896 AND symb_decoder(16#14#)) OR
 					(reg_q896 AND symb_decoder(16#4d#)) OR
 					(reg_q896 AND symb_decoder(16#7b#)) OR
 					(reg_q896 AND symb_decoder(16#0d#)) OR
 					(reg_q896 AND symb_decoder(16#ee#)) OR
 					(reg_q896 AND symb_decoder(16#97#)) OR
 					(reg_q896 AND symb_decoder(16#92#)) OR
 					(reg_q896 AND symb_decoder(16#7a#)) OR
 					(reg_q896 AND symb_decoder(16#67#)) OR
 					(reg_q896 AND symb_decoder(16#91#)) OR
 					(reg_q896 AND symb_decoder(16#3b#)) OR
 					(reg_q896 AND symb_decoder(16#dd#)) OR
 					(reg_q896 AND symb_decoder(16#cb#)) OR
 					(reg_q896 AND symb_decoder(16#38#)) OR
 					(reg_q896 AND symb_decoder(16#cf#)) OR
 					(reg_q896 AND symb_decoder(16#c2#)) OR
 					(reg_q896 AND symb_decoder(16#c7#)) OR
 					(reg_q896 AND symb_decoder(16#bf#)) OR
 					(reg_q896 AND symb_decoder(16#7e#)) OR
 					(reg_q896 AND symb_decoder(16#0f#)) OR
 					(reg_q896 AND symb_decoder(16#ff#)) OR
 					(reg_q896 AND symb_decoder(16#c9#)) OR
 					(reg_q896 AND symb_decoder(16#a0#)) OR
 					(reg_q896 AND symb_decoder(16#18#)) OR
 					(reg_q896 AND symb_decoder(16#9b#)) OR
 					(reg_q896 AND symb_decoder(16#74#)) OR
 					(reg_q896 AND symb_decoder(16#aa#)) OR
 					(reg_q896 AND symb_decoder(16#47#)) OR
 					(reg_q896 AND symb_decoder(16#15#)) OR
 					(reg_q896 AND symb_decoder(16#b2#)) OR
 					(reg_q896 AND symb_decoder(16#1e#)) OR
 					(reg_q896 AND symb_decoder(16#cc#)) OR
 					(reg_q896 AND symb_decoder(16#06#)) OR
 					(reg_q896 AND symb_decoder(16#28#)) OR
 					(reg_q896 AND symb_decoder(16#ae#)) OR
 					(reg_q896 AND symb_decoder(16#da#)) OR
 					(reg_q896 AND symb_decoder(16#3d#)) OR
 					(reg_q896 AND symb_decoder(16#04#)) OR
 					(reg_q896 AND symb_decoder(16#c0#)) OR
 					(reg_q896 AND symb_decoder(16#2f#)) OR
 					(reg_q896 AND symb_decoder(16#12#)) OR
 					(reg_q896 AND symb_decoder(16#62#)) OR
 					(reg_q896 AND symb_decoder(16#57#)) OR
 					(reg_q896 AND symb_decoder(16#9a#)) OR
 					(reg_q896 AND symb_decoder(16#55#)) OR
 					(reg_q896 AND symb_decoder(16#f4#)) OR
 					(reg_q896 AND symb_decoder(16#5f#)) OR
 					(reg_q896 AND symb_decoder(16#e4#)) OR
 					(reg_q896 AND symb_decoder(16#01#)) OR
 					(reg_q896 AND symb_decoder(16#36#)) OR
 					(reg_q896 AND symb_decoder(16#be#)) OR
 					(reg_q896 AND symb_decoder(16#77#)) OR
 					(reg_q896 AND symb_decoder(16#75#)) OR
 					(reg_q896 AND symb_decoder(16#9c#)) OR
 					(reg_q896 AND symb_decoder(16#b3#)) OR
 					(reg_q896 AND symb_decoder(16#6a#)) OR
 					(reg_q896 AND symb_decoder(16#88#)) OR
 					(reg_q896 AND symb_decoder(16#8c#)) OR
 					(reg_q896 AND symb_decoder(16#f0#)) OR
 					(reg_q896 AND symb_decoder(16#60#)) OR
 					(reg_q896 AND symb_decoder(16#59#)) OR
 					(reg_q896 AND symb_decoder(16#1b#)) OR
 					(reg_q896 AND symb_decoder(16#9f#)) OR
 					(reg_q896 AND symb_decoder(16#08#)) OR
 					(reg_q896 AND symb_decoder(16#16#)) OR
 					(reg_q896 AND symb_decoder(16#b9#)) OR
 					(reg_q896 AND symb_decoder(16#24#)) OR
 					(reg_q896 AND symb_decoder(16#e3#)) OR
 					(reg_q896 AND symb_decoder(16#42#)) OR
 					(reg_q896 AND symb_decoder(16#1f#)) OR
 					(reg_q896 AND symb_decoder(16#2d#)) OR
 					(reg_q896 AND symb_decoder(16#e5#)) OR
 					(reg_q896 AND symb_decoder(16#a8#)) OR
 					(reg_q896 AND symb_decoder(16#5a#)) OR
 					(reg_q896 AND symb_decoder(16#48#)) OR
 					(reg_q896 AND symb_decoder(16#bd#)) OR
 					(reg_q896 AND symb_decoder(16#32#)) OR
 					(reg_q896 AND symb_decoder(16#e8#)) OR
 					(reg_q896 AND symb_decoder(16#ca#)) OR
 					(reg_q896 AND symb_decoder(16#d6#)) OR
 					(reg_q896 AND symb_decoder(16#1c#)) OR
 					(reg_q896 AND symb_decoder(16#ce#)) OR
 					(reg_q896 AND symb_decoder(16#68#)) OR
 					(reg_q896 AND symb_decoder(16#72#)) OR
 					(reg_q896 AND symb_decoder(16#f6#)) OR
 					(reg_q896 AND symb_decoder(16#6f#)) OR
 					(reg_q896 AND symb_decoder(16#fa#)) OR
 					(reg_q896 AND symb_decoder(16#40#)) OR
 					(reg_q896 AND symb_decoder(16#f1#)) OR
 					(reg_q896 AND symb_decoder(16#b8#)) OR
 					(reg_q896 AND symb_decoder(16#6b#)) OR
 					(reg_q896 AND symb_decoder(16#63#)) OR
 					(reg_q896 AND symb_decoder(16#5e#)) OR
 					(reg_q896 AND symb_decoder(16#a5#)) OR
 					(reg_q896 AND symb_decoder(16#7d#)) OR
 					(reg_q896 AND symb_decoder(16#d7#)) OR
 					(reg_q896 AND symb_decoder(16#50#)) OR
 					(reg_q896 AND symb_decoder(16#d3#)) OR
 					(reg_q896 AND symb_decoder(16#7f#)) OR
 					(reg_q896 AND symb_decoder(16#99#)) OR
 					(reg_q896 AND symb_decoder(16#86#)) OR
 					(reg_q896 AND symb_decoder(16#35#)) OR
 					(reg_q896 AND symb_decoder(16#eb#)) OR
 					(reg_q896 AND symb_decoder(16#b1#)) OR
 					(reg_q896 AND symb_decoder(16#0b#)) OR
 					(reg_q896 AND symb_decoder(16#11#)) OR
 					(reg_q896 AND symb_decoder(16#e1#)) OR
 					(reg_q896 AND symb_decoder(16#66#)) OR
 					(reg_q896 AND symb_decoder(16#87#)) OR
 					(reg_q896 AND symb_decoder(16#79#)) OR
 					(reg_q896 AND symb_decoder(16#73#)) OR
 					(reg_q896 AND symb_decoder(16#6c#)) OR
 					(reg_q896 AND symb_decoder(16#d1#)) OR
 					(reg_q896 AND symb_decoder(16#33#)) OR
 					(reg_q896 AND symb_decoder(16#70#)) OR
 					(reg_q896 AND symb_decoder(16#ed#)) OR
 					(reg_q896 AND symb_decoder(16#8b#)) OR
 					(reg_q896 AND symb_decoder(16#b7#)) OR
 					(reg_q896 AND symb_decoder(16#34#)) OR
 					(reg_q896 AND symb_decoder(16#1a#)) OR
 					(reg_q896 AND symb_decoder(16#93#)) OR
 					(reg_q896 AND symb_decoder(16#d9#)) OR
 					(reg_q896 AND symb_decoder(16#4c#)) OR
 					(reg_q896 AND symb_decoder(16#bc#)) OR
 					(reg_q896 AND symb_decoder(16#82#)) OR
 					(reg_q896 AND symb_decoder(16#db#)) OR
 					(reg_q896 AND symb_decoder(16#65#)) OR
 					(reg_q896 AND symb_decoder(16#d5#)) OR
 					(reg_q896 AND symb_decoder(16#17#)) OR
 					(reg_q896 AND symb_decoder(16#54#)) OR
 					(reg_q896 AND symb_decoder(16#44#)) OR
 					(reg_q896 AND symb_decoder(16#20#)) OR
 					(reg_q896 AND symb_decoder(16#ef#)) OR
 					(reg_q896 AND symb_decoder(16#76#)) OR
 					(reg_q896 AND symb_decoder(16#a1#)) OR
 					(reg_q896 AND symb_decoder(16#78#)) OR
 					(reg_q896 AND symb_decoder(16#98#)) OR
 					(reg_q896 AND symb_decoder(16#3e#)) OR
 					(reg_q896 AND symb_decoder(16#8f#)) OR
 					(reg_q896 AND symb_decoder(16#b0#)) OR
 					(reg_q896 AND symb_decoder(16#e7#)) OR
 					(reg_q896 AND symb_decoder(16#e9#)) OR
 					(reg_q896 AND symb_decoder(16#45#)) OR
 					(reg_q896 AND symb_decoder(16#c5#)) OR
 					(reg_q896 AND symb_decoder(16#a2#)) OR
 					(reg_q896 AND symb_decoder(16#6d#)) OR
 					(reg_q896 AND symb_decoder(16#c4#)) OR
 					(reg_q896 AND symb_decoder(16#9d#)) OR
 					(reg_q896 AND symb_decoder(16#d4#)) OR
 					(reg_q896 AND symb_decoder(16#6e#)) OR
 					(reg_q896 AND symb_decoder(16#c1#)) OR
 					(reg_q896 AND symb_decoder(16#43#)) OR
 					(reg_q896 AND symb_decoder(16#4a#)) OR
 					(reg_q896 AND symb_decoder(16#03#)) OR
 					(reg_q896 AND symb_decoder(16#ec#)) OR
 					(reg_q896 AND symb_decoder(16#26#)) OR
 					(reg_q896 AND symb_decoder(16#e2#)) OR
 					(reg_q896 AND symb_decoder(16#23#));
reg_q896_init <= '0' ;
	p_reg_q896: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q896 <= reg_q896_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q896 <= reg_q896_init;
        else
          reg_q896 <= reg_q896_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q178_in <= (reg_q178 AND symb_decoder(16#ef#)) OR
 					(reg_q178 AND symb_decoder(16#fd#)) OR
 					(reg_q178 AND symb_decoder(16#f5#)) OR
 					(reg_q178 AND symb_decoder(16#7a#)) OR
 					(reg_q178 AND symb_decoder(16#02#)) OR
 					(reg_q178 AND symb_decoder(16#74#)) OR
 					(reg_q178 AND symb_decoder(16#88#)) OR
 					(reg_q178 AND symb_decoder(16#3a#)) OR
 					(reg_q178 AND symb_decoder(16#6c#)) OR
 					(reg_q178 AND symb_decoder(16#a3#)) OR
 					(reg_q178 AND symb_decoder(16#14#)) OR
 					(reg_q178 AND symb_decoder(16#8b#)) OR
 					(reg_q178 AND symb_decoder(16#32#)) OR
 					(reg_q178 AND symb_decoder(16#04#)) OR
 					(reg_q178 AND symb_decoder(16#98#)) OR
 					(reg_q178 AND symb_decoder(16#0c#)) OR
 					(reg_q178 AND symb_decoder(16#30#)) OR
 					(reg_q178 AND symb_decoder(16#40#)) OR
 					(reg_q178 AND symb_decoder(16#8a#)) OR
 					(reg_q178 AND symb_decoder(16#0d#)) OR
 					(reg_q178 AND symb_decoder(16#c7#)) OR
 					(reg_q178 AND symb_decoder(16#70#)) OR
 					(reg_q178 AND symb_decoder(16#61#)) OR
 					(reg_q178 AND symb_decoder(16#a5#)) OR
 					(reg_q178 AND symb_decoder(16#51#)) OR
 					(reg_q178 AND symb_decoder(16#bd#)) OR
 					(reg_q178 AND symb_decoder(16#d2#)) OR
 					(reg_q178 AND symb_decoder(16#a8#)) OR
 					(reg_q178 AND symb_decoder(16#de#)) OR
 					(reg_q178 AND symb_decoder(16#bc#)) OR
 					(reg_q178 AND symb_decoder(16#c3#)) OR
 					(reg_q178 AND symb_decoder(16#76#)) OR
 					(reg_q178 AND symb_decoder(16#b0#)) OR
 					(reg_q178 AND symb_decoder(16#47#)) OR
 					(reg_q178 AND symb_decoder(16#28#)) OR
 					(reg_q178 AND symb_decoder(16#2f#)) OR
 					(reg_q178 AND symb_decoder(16#0b#)) OR
 					(reg_q178 AND symb_decoder(16#4d#)) OR
 					(reg_q178 AND symb_decoder(16#81#)) OR
 					(reg_q178 AND symb_decoder(16#ca#)) OR
 					(reg_q178 AND symb_decoder(16#1c#)) OR
 					(reg_q178 AND symb_decoder(16#df#)) OR
 					(reg_q178 AND symb_decoder(16#e5#)) OR
 					(reg_q178 AND symb_decoder(16#1d#)) OR
 					(reg_q178 AND symb_decoder(16#27#)) OR
 					(reg_q178 AND symb_decoder(16#49#)) OR
 					(reg_q178 AND symb_decoder(16#19#)) OR
 					(reg_q178 AND symb_decoder(16#8e#)) OR
 					(reg_q178 AND symb_decoder(16#94#)) OR
 					(reg_q178 AND symb_decoder(16#86#)) OR
 					(reg_q178 AND symb_decoder(16#0a#)) OR
 					(reg_q178 AND symb_decoder(16#66#)) OR
 					(reg_q178 AND symb_decoder(16#6e#)) OR
 					(reg_q178 AND symb_decoder(16#fa#)) OR
 					(reg_q178 AND symb_decoder(16#13#)) OR
 					(reg_q178 AND symb_decoder(16#80#)) OR
 					(reg_q178 AND symb_decoder(16#e4#)) OR
 					(reg_q178 AND symb_decoder(16#f2#)) OR
 					(reg_q178 AND symb_decoder(16#e7#)) OR
 					(reg_q178 AND symb_decoder(16#56#)) OR
 					(reg_q178 AND symb_decoder(16#99#)) OR
 					(reg_q178 AND symb_decoder(16#f0#)) OR
 					(reg_q178 AND symb_decoder(16#34#)) OR
 					(reg_q178 AND symb_decoder(16#43#)) OR
 					(reg_q178 AND symb_decoder(16#20#)) OR
 					(reg_q178 AND symb_decoder(16#39#)) OR
 					(reg_q178 AND symb_decoder(16#9e#)) OR
 					(reg_q178 AND symb_decoder(16#7e#)) OR
 					(reg_q178 AND symb_decoder(16#ff#)) OR
 					(reg_q178 AND symb_decoder(16#45#)) OR
 					(reg_q178 AND symb_decoder(16#5e#)) OR
 					(reg_q178 AND symb_decoder(16#bb#)) OR
 					(reg_q178 AND symb_decoder(16#8f#)) OR
 					(reg_q178 AND symb_decoder(16#01#)) OR
 					(reg_q178 AND symb_decoder(16#21#)) OR
 					(reg_q178 AND symb_decoder(16#4b#)) OR
 					(reg_q178 AND symb_decoder(16#b7#)) OR
 					(reg_q178 AND symb_decoder(16#a6#)) OR
 					(reg_q178 AND symb_decoder(16#b2#)) OR
 					(reg_q178 AND symb_decoder(16#50#)) OR
 					(reg_q178 AND symb_decoder(16#15#)) OR
 					(reg_q178 AND symb_decoder(16#e8#)) OR
 					(reg_q178 AND symb_decoder(16#78#)) OR
 					(reg_q178 AND symb_decoder(16#f8#)) OR
 					(reg_q178 AND symb_decoder(16#58#)) OR
 					(reg_q178 AND symb_decoder(16#c1#)) OR
 					(reg_q178 AND symb_decoder(16#18#)) OR
 					(reg_q178 AND symb_decoder(16#9c#)) OR
 					(reg_q178 AND symb_decoder(16#9a#)) OR
 					(reg_q178 AND symb_decoder(16#f9#)) OR
 					(reg_q178 AND symb_decoder(16#91#)) OR
 					(reg_q178 AND symb_decoder(16#92#)) OR
 					(reg_q178 AND symb_decoder(16#9b#)) OR
 					(reg_q178 AND symb_decoder(16#85#)) OR
 					(reg_q178 AND symb_decoder(16#fb#)) OR
 					(reg_q178 AND symb_decoder(16#07#)) OR
 					(reg_q178 AND symb_decoder(16#d4#)) OR
 					(reg_q178 AND symb_decoder(16#68#)) OR
 					(reg_q178 AND symb_decoder(16#37#)) OR
 					(reg_q178 AND symb_decoder(16#5d#)) OR
 					(reg_q178 AND symb_decoder(16#a0#)) OR
 					(reg_q178 AND symb_decoder(16#31#)) OR
 					(reg_q178 AND symb_decoder(16#a9#)) OR
 					(reg_q178 AND symb_decoder(16#cc#)) OR
 					(reg_q178 AND symb_decoder(16#8d#)) OR
 					(reg_q178 AND symb_decoder(16#ab#)) OR
 					(reg_q178 AND symb_decoder(16#9f#)) OR
 					(reg_q178 AND symb_decoder(16#33#)) OR
 					(reg_q178 AND symb_decoder(16#a4#)) OR
 					(reg_q178 AND symb_decoder(16#b1#)) OR
 					(reg_q178 AND symb_decoder(16#cf#)) OR
 					(reg_q178 AND symb_decoder(16#f7#)) OR
 					(reg_q178 AND symb_decoder(16#24#)) OR
 					(reg_q178 AND symb_decoder(16#97#)) OR
 					(reg_q178 AND symb_decoder(16#93#)) OR
 					(reg_q178 AND symb_decoder(16#6d#)) OR
 					(reg_q178 AND symb_decoder(16#11#)) OR
 					(reg_q178 AND symb_decoder(16#ce#)) OR
 					(reg_q178 AND symb_decoder(16#05#)) OR
 					(reg_q178 AND symb_decoder(16#55#)) OR
 					(reg_q178 AND symb_decoder(16#60#)) OR
 					(reg_q178 AND symb_decoder(16#c6#)) OR
 					(reg_q178 AND symb_decoder(16#7d#)) OR
 					(reg_q178 AND symb_decoder(16#7c#)) OR
 					(reg_q178 AND symb_decoder(16#0e#)) OR
 					(reg_q178 AND symb_decoder(16#54#)) OR
 					(reg_q178 AND symb_decoder(16#08#)) OR
 					(reg_q178 AND symb_decoder(16#96#)) OR
 					(reg_q178 AND symb_decoder(16#65#)) OR
 					(reg_q178 AND symb_decoder(16#a2#)) OR
 					(reg_q178 AND symb_decoder(16#48#)) OR
 					(reg_q178 AND symb_decoder(16#03#)) OR
 					(reg_q178 AND symb_decoder(16#c4#)) OR
 					(reg_q178 AND symb_decoder(16#d8#)) OR
 					(reg_q178 AND symb_decoder(16#f6#)) OR
 					(reg_q178 AND symb_decoder(16#2b#)) OR
 					(reg_q178 AND symb_decoder(16#44#)) OR
 					(reg_q178 AND symb_decoder(16#95#)) OR
 					(reg_q178 AND symb_decoder(16#3f#)) OR
 					(reg_q178 AND symb_decoder(16#4a#)) OR
 					(reg_q178 AND symb_decoder(16#3d#)) OR
 					(reg_q178 AND symb_decoder(16#36#)) OR
 					(reg_q178 AND symb_decoder(16#ed#)) OR
 					(reg_q178 AND symb_decoder(16#69#)) OR
 					(reg_q178 AND symb_decoder(16#b8#)) OR
 					(reg_q178 AND symb_decoder(16#90#)) OR
 					(reg_q178 AND symb_decoder(16#ea#)) OR
 					(reg_q178 AND symb_decoder(16#67#)) OR
 					(reg_q178 AND symb_decoder(16#e1#)) OR
 					(reg_q178 AND symb_decoder(16#6a#)) OR
 					(reg_q178 AND symb_decoder(16#7b#)) OR
 					(reg_q178 AND symb_decoder(16#b6#)) OR
 					(reg_q178 AND symb_decoder(16#29#)) OR
 					(reg_q178 AND symb_decoder(16#dd#)) OR
 					(reg_q178 AND symb_decoder(16#1f#)) OR
 					(reg_q178 AND symb_decoder(16#fe#)) OR
 					(reg_q178 AND symb_decoder(16#aa#)) OR
 					(reg_q178 AND symb_decoder(16#cb#)) OR
 					(reg_q178 AND symb_decoder(16#b5#)) OR
 					(reg_q178 AND symb_decoder(16#0f#)) OR
 					(reg_q178 AND symb_decoder(16#7f#)) OR
 					(reg_q178 AND symb_decoder(16#2c#)) OR
 					(reg_q178 AND symb_decoder(16#4f#)) OR
 					(reg_q178 AND symb_decoder(16#db#)) OR
 					(reg_q178 AND symb_decoder(16#ac#)) OR
 					(reg_q178 AND symb_decoder(16#d5#)) OR
 					(reg_q178 AND symb_decoder(16#1b#)) OR
 					(reg_q178 AND symb_decoder(16#cd#)) OR
 					(reg_q178 AND symb_decoder(16#d0#)) OR
 					(reg_q178 AND symb_decoder(16#b4#)) OR
 					(reg_q178 AND symb_decoder(16#6b#)) OR
 					(reg_q178 AND symb_decoder(16#9d#)) OR
 					(reg_q178 AND symb_decoder(16#63#)) OR
 					(reg_q178 AND symb_decoder(16#87#)) OR
 					(reg_q178 AND symb_decoder(16#5c#)) OR
 					(reg_q178 AND symb_decoder(16#e9#)) OR
 					(reg_q178 AND symb_decoder(16#35#)) OR
 					(reg_q178 AND symb_decoder(16#4c#)) OR
 					(reg_q178 AND symb_decoder(16#f4#)) OR
 					(reg_q178 AND symb_decoder(16#64#)) OR
 					(reg_q178 AND symb_decoder(16#d9#)) OR
 					(reg_q178 AND symb_decoder(16#17#)) OR
 					(reg_q178 AND symb_decoder(16#b9#)) OR
 					(reg_q178 AND symb_decoder(16#ec#)) OR
 					(reg_q178 AND symb_decoder(16#af#)) OR
 					(reg_q178 AND symb_decoder(16#f1#)) OR
 					(reg_q178 AND symb_decoder(16#83#)) OR
 					(reg_q178 AND symb_decoder(16#41#)) OR
 					(reg_q178 AND symb_decoder(16#c0#)) OR
 					(reg_q178 AND symb_decoder(16#d3#)) OR
 					(reg_q178 AND symb_decoder(16#53#)) OR
 					(reg_q178 AND symb_decoder(16#fc#)) OR
 					(reg_q178 AND symb_decoder(16#c8#)) OR
 					(reg_q178 AND symb_decoder(16#d6#)) OR
 					(reg_q178 AND symb_decoder(16#84#)) OR
 					(reg_q178 AND symb_decoder(16#d7#)) OR
 					(reg_q178 AND symb_decoder(16#8c#)) OR
 					(reg_q178 AND symb_decoder(16#77#)) OR
 					(reg_q178 AND symb_decoder(16#75#)) OR
 					(reg_q178 AND symb_decoder(16#3e#)) OR
 					(reg_q178 AND symb_decoder(16#52#)) OR
 					(reg_q178 AND symb_decoder(16#ba#)) OR
 					(reg_q178 AND symb_decoder(16#09#)) OR
 					(reg_q178 AND symb_decoder(16#25#)) OR
 					(reg_q178 AND symb_decoder(16#ad#)) OR
 					(reg_q178 AND symb_decoder(16#b3#)) OR
 					(reg_q178 AND symb_decoder(16#2e#)) OR
 					(reg_q178 AND symb_decoder(16#a1#)) OR
 					(reg_q178 AND symb_decoder(16#00#)) OR
 					(reg_q178 AND symb_decoder(16#f3#)) OR
 					(reg_q178 AND symb_decoder(16#be#)) OR
 					(reg_q178 AND symb_decoder(16#22#)) OR
 					(reg_q178 AND symb_decoder(16#82#)) OR
 					(reg_q178 AND symb_decoder(16#2d#)) OR
 					(reg_q178 AND symb_decoder(16#e3#)) OR
 					(reg_q178 AND symb_decoder(16#4e#)) OR
 					(reg_q178 AND symb_decoder(16#5a#)) OR
 					(reg_q178 AND symb_decoder(16#57#)) OR
 					(reg_q178 AND symb_decoder(16#bf#)) OR
 					(reg_q178 AND symb_decoder(16#16#)) OR
 					(reg_q178 AND symb_decoder(16#38#)) OR
 					(reg_q178 AND symb_decoder(16#89#)) OR
 					(reg_q178 AND symb_decoder(16#1a#)) OR
 					(reg_q178 AND symb_decoder(16#72#)) OR
 					(reg_q178 AND symb_decoder(16#10#)) OR
 					(reg_q178 AND symb_decoder(16#59#)) OR
 					(reg_q178 AND symb_decoder(16#a7#)) OR
 					(reg_q178 AND symb_decoder(16#46#)) OR
 					(reg_q178 AND symb_decoder(16#6f#)) OR
 					(reg_q178 AND symb_decoder(16#ee#)) OR
 					(reg_q178 AND symb_decoder(16#2a#)) OR
 					(reg_q178 AND symb_decoder(16#1e#)) OR
 					(reg_q178 AND symb_decoder(16#e2#)) OR
 					(reg_q178 AND symb_decoder(16#eb#)) OR
 					(reg_q178 AND symb_decoder(16#e6#)) OR
 					(reg_q178 AND symb_decoder(16#42#)) OR
 					(reg_q178 AND symb_decoder(16#ae#)) OR
 					(reg_q178 AND symb_decoder(16#d1#)) OR
 					(reg_q178 AND symb_decoder(16#73#)) OR
 					(reg_q178 AND symb_decoder(16#c9#)) OR
 					(reg_q178 AND symb_decoder(16#26#)) OR
 					(reg_q178 AND symb_decoder(16#3c#)) OR
 					(reg_q178 AND symb_decoder(16#71#)) OR
 					(reg_q178 AND symb_decoder(16#06#)) OR
 					(reg_q178 AND symb_decoder(16#79#)) OR
 					(reg_q178 AND symb_decoder(16#3b#)) OR
 					(reg_q178 AND symb_decoder(16#e0#)) OR
 					(reg_q178 AND symb_decoder(16#c5#)) OR
 					(reg_q178 AND symb_decoder(16#dc#)) OR
 					(reg_q178 AND symb_decoder(16#5b#)) OR
 					(reg_q178 AND symb_decoder(16#12#)) OR
 					(reg_q178 AND symb_decoder(16#da#)) OR
 					(reg_q178 AND symb_decoder(16#62#)) OR
 					(reg_q178 AND symb_decoder(16#23#)) OR
 					(reg_q178 AND symb_decoder(16#c2#)) OR
 					(reg_q178 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#));
reg_q178_init <= '0' ;
	p_reg_q178: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q178 <= reg_q178_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q178 <= reg_q178_init;
        else
          reg_q178 <= reg_q178_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1812_in <= (reg_q1810 AND symb_decoder(16#45#)) OR
 					(reg_q1810 AND symb_decoder(16#65#));
reg_q1812_init <= '0' ;
	p_reg_q1812: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1812 <= reg_q1812_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1812 <= reg_q1812_init;
        else
          reg_q1812 <= reg_q1812_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1814_in <= (reg_q1812 AND symb_decoder(16#72#)) OR
 					(reg_q1812 AND symb_decoder(16#52#));
reg_q1814_init <= '0' ;
	p_reg_q1814: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1814 <= reg_q1814_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1814 <= reg_q1814_init;
        else
          reg_q1814 <= reg_q1814_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1013_in <= (reg_q1013 AND symb_decoder(16#aa#)) OR
 					(reg_q1013 AND symb_decoder(16#30#)) OR
 					(reg_q1013 AND symb_decoder(16#62#)) OR
 					(reg_q1013 AND symb_decoder(16#3d#)) OR
 					(reg_q1013 AND symb_decoder(16#cd#)) OR
 					(reg_q1013 AND symb_decoder(16#e6#)) OR
 					(reg_q1013 AND symb_decoder(16#22#)) OR
 					(reg_q1013 AND symb_decoder(16#b7#)) OR
 					(reg_q1013 AND symb_decoder(16#d8#)) OR
 					(reg_q1013 AND symb_decoder(16#d6#)) OR
 					(reg_q1013 AND symb_decoder(16#b9#)) OR
 					(reg_q1013 AND symb_decoder(16#05#)) OR
 					(reg_q1013 AND symb_decoder(16#16#)) OR
 					(reg_q1013 AND symb_decoder(16#2b#)) OR
 					(reg_q1013 AND symb_decoder(16#55#)) OR
 					(reg_q1013 AND symb_decoder(16#95#)) OR
 					(reg_q1013 AND symb_decoder(16#e8#)) OR
 					(reg_q1013 AND symb_decoder(16#97#)) OR
 					(reg_q1013 AND symb_decoder(16#db#)) OR
 					(reg_q1013 AND symb_decoder(16#ff#)) OR
 					(reg_q1013 AND symb_decoder(16#4e#)) OR
 					(reg_q1013 AND symb_decoder(16#ab#)) OR
 					(reg_q1013 AND symb_decoder(16#57#)) OR
 					(reg_q1013 AND symb_decoder(16#5a#)) OR
 					(reg_q1013 AND symb_decoder(16#d3#)) OR
 					(reg_q1013 AND symb_decoder(16#70#)) OR
 					(reg_q1013 AND symb_decoder(16#7c#)) OR
 					(reg_q1013 AND symb_decoder(16#c1#)) OR
 					(reg_q1013 AND symb_decoder(16#6d#)) OR
 					(reg_q1013 AND symb_decoder(16#6e#)) OR
 					(reg_q1013 AND symb_decoder(16#53#)) OR
 					(reg_q1013 AND symb_decoder(16#c8#)) OR
 					(reg_q1013 AND symb_decoder(16#8c#)) OR
 					(reg_q1013 AND symb_decoder(16#35#)) OR
 					(reg_q1013 AND symb_decoder(16#18#)) OR
 					(reg_q1013 AND symb_decoder(16#74#)) OR
 					(reg_q1013 AND symb_decoder(16#49#)) OR
 					(reg_q1013 AND symb_decoder(16#76#)) OR
 					(reg_q1013 AND symb_decoder(16#cf#)) OR
 					(reg_q1013 AND symb_decoder(16#33#)) OR
 					(reg_q1013 AND symb_decoder(16#1a#)) OR
 					(reg_q1013 AND symb_decoder(16#cb#)) OR
 					(reg_q1013 AND symb_decoder(16#fd#)) OR
 					(reg_q1013 AND symb_decoder(16#82#)) OR
 					(reg_q1013 AND symb_decoder(16#7b#)) OR
 					(reg_q1013 AND symb_decoder(16#0d#)) OR
 					(reg_q1013 AND symb_decoder(16#d0#)) OR
 					(reg_q1013 AND symb_decoder(16#34#)) OR
 					(reg_q1013 AND symb_decoder(16#13#)) OR
 					(reg_q1013 AND symb_decoder(16#fc#)) OR
 					(reg_q1013 AND symb_decoder(16#66#)) OR
 					(reg_q1013 AND symb_decoder(16#bf#)) OR
 					(reg_q1013 AND symb_decoder(16#c2#)) OR
 					(reg_q1013 AND symb_decoder(16#b6#)) OR
 					(reg_q1013 AND symb_decoder(16#51#)) OR
 					(reg_q1013 AND symb_decoder(16#17#)) OR
 					(reg_q1013 AND symb_decoder(16#3a#)) OR
 					(reg_q1013 AND symb_decoder(16#10#)) OR
 					(reg_q1013 AND symb_decoder(16#7d#)) OR
 					(reg_q1013 AND symb_decoder(16#56#)) OR
 					(reg_q1013 AND symb_decoder(16#f9#)) OR
 					(reg_q1013 AND symb_decoder(16#e0#)) OR
 					(reg_q1013 AND symb_decoder(16#e9#)) OR
 					(reg_q1013 AND symb_decoder(16#ae#)) OR
 					(reg_q1013 AND symb_decoder(16#fb#)) OR
 					(reg_q1013 AND symb_decoder(16#48#)) OR
 					(reg_q1013 AND symb_decoder(16#89#)) OR
 					(reg_q1013 AND symb_decoder(16#ce#)) OR
 					(reg_q1013 AND symb_decoder(16#b8#)) OR
 					(reg_q1013 AND symb_decoder(16#e1#)) OR
 					(reg_q1013 AND symb_decoder(16#c4#)) OR
 					(reg_q1013 AND symb_decoder(16#a6#)) OR
 					(reg_q1013 AND symb_decoder(16#26#)) OR
 					(reg_q1013 AND symb_decoder(16#a9#)) OR
 					(reg_q1013 AND symb_decoder(16#6b#)) OR
 					(reg_q1013 AND symb_decoder(16#94#)) OR
 					(reg_q1013 AND symb_decoder(16#cc#)) OR
 					(reg_q1013 AND symb_decoder(16#0c#)) OR
 					(reg_q1013 AND symb_decoder(16#38#)) OR
 					(reg_q1013 AND symb_decoder(16#bb#)) OR
 					(reg_q1013 AND symb_decoder(16#84#)) OR
 					(reg_q1013 AND symb_decoder(16#8e#)) OR
 					(reg_q1013 AND symb_decoder(16#93#)) OR
 					(reg_q1013 AND symb_decoder(16#06#)) OR
 					(reg_q1013 AND symb_decoder(16#91#)) OR
 					(reg_q1013 AND symb_decoder(16#04#)) OR
 					(reg_q1013 AND symb_decoder(16#f7#)) OR
 					(reg_q1013 AND symb_decoder(16#41#)) OR
 					(reg_q1013 AND symb_decoder(16#80#)) OR
 					(reg_q1013 AND symb_decoder(16#b3#)) OR
 					(reg_q1013 AND symb_decoder(16#0b#)) OR
 					(reg_q1013 AND symb_decoder(16#3f#)) OR
 					(reg_q1013 AND symb_decoder(16#00#)) OR
 					(reg_q1013 AND symb_decoder(16#12#)) OR
 					(reg_q1013 AND symb_decoder(16#8d#)) OR
 					(reg_q1013 AND symb_decoder(16#e7#)) OR
 					(reg_q1013 AND symb_decoder(16#9a#)) OR
 					(reg_q1013 AND symb_decoder(16#61#)) OR
 					(reg_q1013 AND symb_decoder(16#0f#)) OR
 					(reg_q1013 AND symb_decoder(16#40#)) OR
 					(reg_q1013 AND symb_decoder(16#1c#)) OR
 					(reg_q1013 AND symb_decoder(16#08#)) OR
 					(reg_q1013 AND symb_decoder(16#e4#)) OR
 					(reg_q1013 AND symb_decoder(16#eb#)) OR
 					(reg_q1013 AND symb_decoder(16#ba#)) OR
 					(reg_q1013 AND symb_decoder(16#f8#)) OR
 					(reg_q1013 AND symb_decoder(16#c5#)) OR
 					(reg_q1013 AND symb_decoder(16#ee#)) OR
 					(reg_q1013 AND symb_decoder(16#a0#)) OR
 					(reg_q1013 AND symb_decoder(16#52#)) OR
 					(reg_q1013 AND symb_decoder(16#c9#)) OR
 					(reg_q1013 AND symb_decoder(16#de#)) OR
 					(reg_q1013 AND symb_decoder(16#b1#)) OR
 					(reg_q1013 AND symb_decoder(16#fa#)) OR
 					(reg_q1013 AND symb_decoder(16#b2#)) OR
 					(reg_q1013 AND symb_decoder(16#a4#)) OR
 					(reg_q1013 AND symb_decoder(16#fe#)) OR
 					(reg_q1013 AND symb_decoder(16#8f#)) OR
 					(reg_q1013 AND symb_decoder(16#ad#)) OR
 					(reg_q1013 AND symb_decoder(16#9b#)) OR
 					(reg_q1013 AND symb_decoder(16#23#)) OR
 					(reg_q1013 AND symb_decoder(16#2e#)) OR
 					(reg_q1013 AND symb_decoder(16#54#)) OR
 					(reg_q1013 AND symb_decoder(16#f6#)) OR
 					(reg_q1013 AND symb_decoder(16#77#)) OR
 					(reg_q1013 AND symb_decoder(16#d4#)) OR
 					(reg_q1013 AND symb_decoder(16#0a#)) OR
 					(reg_q1013 AND symb_decoder(16#8b#)) OR
 					(reg_q1013 AND symb_decoder(16#50#)) OR
 					(reg_q1013 AND symb_decoder(16#32#)) OR
 					(reg_q1013 AND symb_decoder(16#a3#)) OR
 					(reg_q1013 AND symb_decoder(16#a2#)) OR
 					(reg_q1013 AND symb_decoder(16#6f#)) OR
 					(reg_q1013 AND symb_decoder(16#11#)) OR
 					(reg_q1013 AND symb_decoder(16#ec#)) OR
 					(reg_q1013 AND symb_decoder(16#9c#)) OR
 					(reg_q1013 AND symb_decoder(16#da#)) OR
 					(reg_q1013 AND symb_decoder(16#d9#)) OR
 					(reg_q1013 AND symb_decoder(16#dd#)) OR
 					(reg_q1013 AND symb_decoder(16#7f#)) OR
 					(reg_q1013 AND symb_decoder(16#21#)) OR
 					(reg_q1013 AND symb_decoder(16#58#)) OR
 					(reg_q1013 AND symb_decoder(16#5d#)) OR
 					(reg_q1013 AND symb_decoder(16#71#)) OR
 					(reg_q1013 AND symb_decoder(16#5b#)) OR
 					(reg_q1013 AND symb_decoder(16#14#)) OR
 					(reg_q1013 AND symb_decoder(16#87#)) OR
 					(reg_q1013 AND symb_decoder(16#39#)) OR
 					(reg_q1013 AND symb_decoder(16#e5#)) OR
 					(reg_q1013 AND symb_decoder(16#59#)) OR
 					(reg_q1013 AND symb_decoder(16#a5#)) OR
 					(reg_q1013 AND symb_decoder(16#6c#)) OR
 					(reg_q1013 AND symb_decoder(16#09#)) OR
 					(reg_q1013 AND symb_decoder(16#46#)) OR
 					(reg_q1013 AND symb_decoder(16#f3#)) OR
 					(reg_q1013 AND symb_decoder(16#1e#)) OR
 					(reg_q1013 AND symb_decoder(16#bd#)) OR
 					(reg_q1013 AND symb_decoder(16#72#)) OR
 					(reg_q1013 AND symb_decoder(16#ef#)) OR
 					(reg_q1013 AND symb_decoder(16#b4#)) OR
 					(reg_q1013 AND symb_decoder(16#dc#)) OR
 					(reg_q1013 AND symb_decoder(16#07#)) OR
 					(reg_q1013 AND symb_decoder(16#86#)) OR
 					(reg_q1013 AND symb_decoder(16#44#)) OR
 					(reg_q1013 AND symb_decoder(16#47#)) OR
 					(reg_q1013 AND symb_decoder(16#28#)) OR
 					(reg_q1013 AND symb_decoder(16#b5#)) OR
 					(reg_q1013 AND symb_decoder(16#c3#)) OR
 					(reg_q1013 AND symb_decoder(16#02#)) OR
 					(reg_q1013 AND symb_decoder(16#ea#)) OR
 					(reg_q1013 AND symb_decoder(16#6a#)) OR
 					(reg_q1013 AND symb_decoder(16#7a#)) OR
 					(reg_q1013 AND symb_decoder(16#42#)) OR
 					(reg_q1013 AND symb_decoder(16#36#)) OR
 					(reg_q1013 AND symb_decoder(16#5e#)) OR
 					(reg_q1013 AND symb_decoder(16#73#)) OR
 					(reg_q1013 AND symb_decoder(16#f5#)) OR
 					(reg_q1013 AND symb_decoder(16#19#)) OR
 					(reg_q1013 AND symb_decoder(16#e2#)) OR
 					(reg_q1013 AND symb_decoder(16#2a#)) OR
 					(reg_q1013 AND symb_decoder(16#4c#)) OR
 					(reg_q1013 AND symb_decoder(16#9e#)) OR
 					(reg_q1013 AND symb_decoder(16#f4#)) OR
 					(reg_q1013 AND symb_decoder(16#bc#)) OR
 					(reg_q1013 AND symb_decoder(16#27#)) OR
 					(reg_q1013 AND symb_decoder(16#3e#)) OR
 					(reg_q1013 AND symb_decoder(16#a1#)) OR
 					(reg_q1013 AND symb_decoder(16#90#)) OR
 					(reg_q1013 AND symb_decoder(16#64#)) OR
 					(reg_q1013 AND symb_decoder(16#d2#)) OR
 					(reg_q1013 AND symb_decoder(16#20#)) OR
 					(reg_q1013 AND symb_decoder(16#63#)) OR
 					(reg_q1013 AND symb_decoder(16#8a#)) OR
 					(reg_q1013 AND symb_decoder(16#ed#)) OR
 					(reg_q1013 AND symb_decoder(16#9d#)) OR
 					(reg_q1013 AND symb_decoder(16#7e#)) OR
 					(reg_q1013 AND symb_decoder(16#a7#)) OR
 					(reg_q1013 AND symb_decoder(16#2f#)) OR
 					(reg_q1013 AND symb_decoder(16#c7#)) OR
 					(reg_q1013 AND symb_decoder(16#c0#)) OR
 					(reg_q1013 AND symb_decoder(16#ca#)) OR
 					(reg_q1013 AND symb_decoder(16#15#)) OR
 					(reg_q1013 AND symb_decoder(16#43#)) OR
 					(reg_q1013 AND symb_decoder(16#85#)) OR
 					(reg_q1013 AND symb_decoder(16#45#)) OR
 					(reg_q1013 AND symb_decoder(16#67#)) OR
 					(reg_q1013 AND symb_decoder(16#4b#)) OR
 					(reg_q1013 AND symb_decoder(16#24#)) OR
 					(reg_q1013 AND symb_decoder(16#d7#)) OR
 					(reg_q1013 AND symb_decoder(16#d5#)) OR
 					(reg_q1013 AND symb_decoder(16#f0#)) OR
 					(reg_q1013 AND symb_decoder(16#ac#)) OR
 					(reg_q1013 AND symb_decoder(16#25#)) OR
 					(reg_q1013 AND symb_decoder(16#df#)) OR
 					(reg_q1013 AND symb_decoder(16#9f#)) OR
 					(reg_q1013 AND symb_decoder(16#c6#)) OR
 					(reg_q1013 AND symb_decoder(16#1d#)) OR
 					(reg_q1013 AND symb_decoder(16#78#)) OR
 					(reg_q1013 AND symb_decoder(16#88#)) OR
 					(reg_q1013 AND symb_decoder(16#29#)) OR
 					(reg_q1013 AND symb_decoder(16#01#)) OR
 					(reg_q1013 AND symb_decoder(16#d1#)) OR
 					(reg_q1013 AND symb_decoder(16#79#)) OR
 					(reg_q1013 AND symb_decoder(16#5c#)) OR
 					(reg_q1013 AND symb_decoder(16#1b#)) OR
 					(reg_q1013 AND symb_decoder(16#af#)) OR
 					(reg_q1013 AND symb_decoder(16#31#)) OR
 					(reg_q1013 AND symb_decoder(16#92#)) OR
 					(reg_q1013 AND symb_decoder(16#75#)) OR
 					(reg_q1013 AND symb_decoder(16#81#)) OR
 					(reg_q1013 AND symb_decoder(16#3c#)) OR
 					(reg_q1013 AND symb_decoder(16#5f#)) OR
 					(reg_q1013 AND symb_decoder(16#3b#)) OR
 					(reg_q1013 AND symb_decoder(16#0e#)) OR
 					(reg_q1013 AND symb_decoder(16#96#)) OR
 					(reg_q1013 AND symb_decoder(16#2c#)) OR
 					(reg_q1013 AND symb_decoder(16#69#)) OR
 					(reg_q1013 AND symb_decoder(16#a8#)) OR
 					(reg_q1013 AND symb_decoder(16#99#)) OR
 					(reg_q1013 AND symb_decoder(16#b0#)) OR
 					(reg_q1013 AND symb_decoder(16#60#)) OR
 					(reg_q1013 AND symb_decoder(16#4d#)) OR
 					(reg_q1013 AND symb_decoder(16#e3#)) OR
 					(reg_q1013 AND symb_decoder(16#4f#)) OR
 					(reg_q1013 AND symb_decoder(16#be#)) OR
 					(reg_q1013 AND symb_decoder(16#f2#)) OR
 					(reg_q1013 AND symb_decoder(16#4a#)) OR
 					(reg_q1013 AND symb_decoder(16#03#)) OR
 					(reg_q1013 AND symb_decoder(16#2d#)) OR
 					(reg_q1013 AND symb_decoder(16#37#)) OR
 					(reg_q1013 AND symb_decoder(16#68#)) OR
 					(reg_q1013 AND symb_decoder(16#1f#)) OR
 					(reg_q1013 AND symb_decoder(16#98#)) OR
 					(reg_q1013 AND symb_decoder(16#65#)) OR
 					(reg_q1013 AND symb_decoder(16#83#)) OR
 					(reg_q1013 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#));
reg_q1013_init <= '0' ;
	p_reg_q1013: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1013 <= reg_q1013_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1013 <= reg_q1013_init;
        else
          reg_q1013 <= reg_q1013_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2695_in <= '0' ;
reg_q2695_init <= '1' ;
	p_reg_q2695: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2695 <= reg_q2695_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2695 <= reg_q2695_init;
        else
          reg_q2695 <= reg_q2695_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q779_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q779 AND symb_decoder(16#e6#)) OR
 					(reg_q779 AND symb_decoder(16#f4#)) OR
 					(reg_q779 AND symb_decoder(16#5e#)) OR
 					(reg_q779 AND symb_decoder(16#3d#)) OR
 					(reg_q779 AND symb_decoder(16#a2#)) OR
 					(reg_q779 AND symb_decoder(16#37#)) OR
 					(reg_q779 AND symb_decoder(16#da#)) OR
 					(reg_q779 AND symb_decoder(16#30#)) OR
 					(reg_q779 AND symb_decoder(16#70#)) OR
 					(reg_q779 AND symb_decoder(16#0e#)) OR
 					(reg_q779 AND symb_decoder(16#0d#)) OR
 					(reg_q779 AND symb_decoder(16#42#)) OR
 					(reg_q779 AND symb_decoder(16#54#)) OR
 					(reg_q779 AND symb_decoder(16#cf#)) OR
 					(reg_q779 AND symb_decoder(16#f1#)) OR
 					(reg_q779 AND symb_decoder(16#5d#)) OR
 					(reg_q779 AND symb_decoder(16#fd#)) OR
 					(reg_q779 AND symb_decoder(16#0b#)) OR
 					(reg_q779 AND symb_decoder(16#01#)) OR
 					(reg_q779 AND symb_decoder(16#ec#)) OR
 					(reg_q779 AND symb_decoder(16#0a#)) OR
 					(reg_q779 AND symb_decoder(16#2a#)) OR
 					(reg_q779 AND symb_decoder(16#5c#)) OR
 					(reg_q779 AND symb_decoder(16#b1#)) OR
 					(reg_q779 AND symb_decoder(16#75#)) OR
 					(reg_q779 AND symb_decoder(16#81#)) OR
 					(reg_q779 AND symb_decoder(16#08#)) OR
 					(reg_q779 AND symb_decoder(16#04#)) OR
 					(reg_q779 AND symb_decoder(16#4a#)) OR
 					(reg_q779 AND symb_decoder(16#b4#)) OR
 					(reg_q779 AND symb_decoder(16#8a#)) OR
 					(reg_q779 AND symb_decoder(16#c1#)) OR
 					(reg_q779 AND symb_decoder(16#a3#)) OR
 					(reg_q779 AND symb_decoder(16#ae#)) OR
 					(reg_q779 AND symb_decoder(16#5a#)) OR
 					(reg_q779 AND symb_decoder(16#bf#)) OR
 					(reg_q779 AND symb_decoder(16#26#)) OR
 					(reg_q779 AND symb_decoder(16#45#)) OR
 					(reg_q779 AND symb_decoder(16#eb#)) OR
 					(reg_q779 AND symb_decoder(16#05#)) OR
 					(reg_q779 AND symb_decoder(16#31#)) OR
 					(reg_q779 AND symb_decoder(16#ef#)) OR
 					(reg_q779 AND symb_decoder(16#60#)) OR
 					(reg_q779 AND symb_decoder(16#d3#)) OR
 					(reg_q779 AND symb_decoder(16#3b#)) OR
 					(reg_q779 AND symb_decoder(16#46#)) OR
 					(reg_q779 AND symb_decoder(16#89#)) OR
 					(reg_q779 AND symb_decoder(16#80#)) OR
 					(reg_q779 AND symb_decoder(16#f9#)) OR
 					(reg_q779 AND symb_decoder(16#d8#)) OR
 					(reg_q779 AND symb_decoder(16#02#)) OR
 					(reg_q779 AND symb_decoder(16#50#)) OR
 					(reg_q779 AND symb_decoder(16#7d#)) OR
 					(reg_q779 AND symb_decoder(16#4e#)) OR
 					(reg_q779 AND symb_decoder(16#aa#)) OR
 					(reg_q779 AND symb_decoder(16#90#)) OR
 					(reg_q779 AND symb_decoder(16#9e#)) OR
 					(reg_q779 AND symb_decoder(16#68#)) OR
 					(reg_q779 AND symb_decoder(16#5b#)) OR
 					(reg_q779 AND symb_decoder(16#d0#)) OR
 					(reg_q779 AND symb_decoder(16#cd#)) OR
 					(reg_q779 AND symb_decoder(16#ee#)) OR
 					(reg_q779 AND symb_decoder(16#17#)) OR
 					(reg_q779 AND symb_decoder(16#fe#)) OR
 					(reg_q779 AND symb_decoder(16#58#)) OR
 					(reg_q779 AND symb_decoder(16#c6#)) OR
 					(reg_q779 AND symb_decoder(16#d5#)) OR
 					(reg_q779 AND symb_decoder(16#b2#)) OR
 					(reg_q779 AND symb_decoder(16#78#)) OR
 					(reg_q779 AND symb_decoder(16#6a#)) OR
 					(reg_q779 AND symb_decoder(16#12#)) OR
 					(reg_q779 AND symb_decoder(16#cb#)) OR
 					(reg_q779 AND symb_decoder(16#ea#)) OR
 					(reg_q779 AND symb_decoder(16#51#)) OR
 					(reg_q779 AND symb_decoder(16#82#)) OR
 					(reg_q779 AND symb_decoder(16#0c#)) OR
 					(reg_q779 AND symb_decoder(16#77#)) OR
 					(reg_q779 AND symb_decoder(16#b7#)) OR
 					(reg_q779 AND symb_decoder(16#d6#)) OR
 					(reg_q779 AND symb_decoder(16#74#)) OR
 					(reg_q779 AND symb_decoder(16#39#)) OR
 					(reg_q779 AND symb_decoder(16#63#)) OR
 					(reg_q779 AND symb_decoder(16#dc#)) OR
 					(reg_q779 AND symb_decoder(16#35#)) OR
 					(reg_q779 AND symb_decoder(16#8b#)) OR
 					(reg_q779 AND symb_decoder(16#ca#)) OR
 					(reg_q779 AND symb_decoder(16#a5#)) OR
 					(reg_q779 AND symb_decoder(16#e1#)) OR
 					(reg_q779 AND symb_decoder(16#7c#)) OR
 					(reg_q779 AND symb_decoder(16#22#)) OR
 					(reg_q779 AND symb_decoder(16#3c#)) OR
 					(reg_q779 AND symb_decoder(16#34#)) OR
 					(reg_q779 AND symb_decoder(16#4f#)) OR
 					(reg_q779 AND symb_decoder(16#69#)) OR
 					(reg_q779 AND symb_decoder(16#41#)) OR
 					(reg_q779 AND symb_decoder(16#40#)) OR
 					(reg_q779 AND symb_decoder(16#e4#)) OR
 					(reg_q779 AND symb_decoder(16#47#)) OR
 					(reg_q779 AND symb_decoder(16#4d#)) OR
 					(reg_q779 AND symb_decoder(16#3e#)) OR
 					(reg_q779 AND symb_decoder(16#6c#)) OR
 					(reg_q779 AND symb_decoder(16#10#)) OR
 					(reg_q779 AND symb_decoder(16#bd#)) OR
 					(reg_q779 AND symb_decoder(16#dd#)) OR
 					(reg_q779 AND symb_decoder(16#32#)) OR
 					(reg_q779 AND symb_decoder(16#66#)) OR
 					(reg_q779 AND symb_decoder(16#f8#)) OR
 					(reg_q779 AND symb_decoder(16#59#)) OR
 					(reg_q779 AND symb_decoder(16#a1#)) OR
 					(reg_q779 AND symb_decoder(16#1d#)) OR
 					(reg_q779 AND symb_decoder(16#97#)) OR
 					(reg_q779 AND symb_decoder(16#2c#)) OR
 					(reg_q779 AND symb_decoder(16#df#)) OR
 					(reg_q779 AND symb_decoder(16#1a#)) OR
 					(reg_q779 AND symb_decoder(16#6b#)) OR
 					(reg_q779 AND symb_decoder(16#73#)) OR
 					(reg_q779 AND symb_decoder(16#6d#)) OR
 					(reg_q779 AND symb_decoder(16#1f#)) OR
 					(reg_q779 AND symb_decoder(16#a7#)) OR
 					(reg_q779 AND symb_decoder(16#c5#)) OR
 					(reg_q779 AND symb_decoder(16#28#)) OR
 					(reg_q779 AND symb_decoder(16#d1#)) OR
 					(reg_q779 AND symb_decoder(16#07#)) OR
 					(reg_q779 AND symb_decoder(16#7b#)) OR
 					(reg_q779 AND symb_decoder(16#18#)) OR
 					(reg_q779 AND symb_decoder(16#94#)) OR
 					(reg_q779 AND symb_decoder(16#a9#)) OR
 					(reg_q779 AND symb_decoder(16#9d#)) OR
 					(reg_q779 AND symb_decoder(16#49#)) OR
 					(reg_q779 AND symb_decoder(16#ab#)) OR
 					(reg_q779 AND symb_decoder(16#88#)) OR
 					(reg_q779 AND symb_decoder(16#e3#)) OR
 					(reg_q779 AND symb_decoder(16#86#)) OR
 					(reg_q779 AND symb_decoder(16#23#)) OR
 					(reg_q779 AND symb_decoder(16#cc#)) OR
 					(reg_q779 AND symb_decoder(16#fa#)) OR
 					(reg_q779 AND symb_decoder(16#16#)) OR
 					(reg_q779 AND symb_decoder(16#c4#)) OR
 					(reg_q779 AND symb_decoder(16#b8#)) OR
 					(reg_q779 AND symb_decoder(16#27#)) OR
 					(reg_q779 AND symb_decoder(16#f6#)) OR
 					(reg_q779 AND symb_decoder(16#84#)) OR
 					(reg_q779 AND symb_decoder(16#fc#)) OR
 					(reg_q779 AND symb_decoder(16#67#)) OR
 					(reg_q779 AND symb_decoder(16#e9#)) OR
 					(reg_q779 AND symb_decoder(16#e0#)) OR
 					(reg_q779 AND symb_decoder(16#ce#)) OR
 					(reg_q779 AND symb_decoder(16#c2#)) OR
 					(reg_q779 AND symb_decoder(16#f3#)) OR
 					(reg_q779 AND symb_decoder(16#a0#)) OR
 					(reg_q779 AND symb_decoder(16#76#)) OR
 					(reg_q779 AND symb_decoder(16#b3#)) OR
 					(reg_q779 AND symb_decoder(16#38#)) OR
 					(reg_q779 AND symb_decoder(16#b6#)) OR
 					(reg_q779 AND symb_decoder(16#87#)) OR
 					(reg_q779 AND symb_decoder(16#af#)) OR
 					(reg_q779 AND symb_decoder(16#9c#)) OR
 					(reg_q779 AND symb_decoder(16#ff#)) OR
 					(reg_q779 AND symb_decoder(16#9a#)) OR
 					(reg_q779 AND symb_decoder(16#d7#)) OR
 					(reg_q779 AND symb_decoder(16#ed#)) OR
 					(reg_q779 AND symb_decoder(16#c8#)) OR
 					(reg_q779 AND symb_decoder(16#1e#)) OR
 					(reg_q779 AND symb_decoder(16#8c#)) OR
 					(reg_q779 AND symb_decoder(16#06#)) OR
 					(reg_q779 AND symb_decoder(16#24#)) OR
 					(reg_q779 AND symb_decoder(16#ba#)) OR
 					(reg_q779 AND symb_decoder(16#4c#)) OR
 					(reg_q779 AND symb_decoder(16#20#)) OR
 					(reg_q779 AND symb_decoder(16#a6#)) OR
 					(reg_q779 AND symb_decoder(16#8d#)) OR
 					(reg_q779 AND symb_decoder(16#c0#)) OR
 					(reg_q779 AND symb_decoder(16#7f#)) OR
 					(reg_q779 AND symb_decoder(16#e2#)) OR
 					(reg_q779 AND symb_decoder(16#64#)) OR
 					(reg_q779 AND symb_decoder(16#55#)) OR
 					(reg_q779 AND symb_decoder(16#85#)) OR
 					(reg_q779 AND symb_decoder(16#25#)) OR
 					(reg_q779 AND symb_decoder(16#19#)) OR
 					(reg_q779 AND symb_decoder(16#72#)) OR
 					(reg_q779 AND symb_decoder(16#9b#)) OR
 					(reg_q779 AND symb_decoder(16#6e#)) OR
 					(reg_q779 AND symb_decoder(16#e7#)) OR
 					(reg_q779 AND symb_decoder(16#09#)) OR
 					(reg_q779 AND symb_decoder(16#36#)) OR
 					(reg_q779 AND symb_decoder(16#15#)) OR
 					(reg_q779 AND symb_decoder(16#db#)) OR
 					(reg_q779 AND symb_decoder(16#f2#)) OR
 					(reg_q779 AND symb_decoder(16#53#)) OR
 					(reg_q779 AND symb_decoder(16#2d#)) OR
 					(reg_q779 AND symb_decoder(16#8e#)) OR
 					(reg_q779 AND symb_decoder(16#b5#)) OR
 					(reg_q779 AND symb_decoder(16#bc#)) OR
 					(reg_q779 AND symb_decoder(16#c3#)) OR
 					(reg_q779 AND symb_decoder(16#1b#)) OR
 					(reg_q779 AND symb_decoder(16#48#)) OR
 					(reg_q779 AND symb_decoder(16#43#)) OR
 					(reg_q779 AND symb_decoder(16#00#)) OR
 					(reg_q779 AND symb_decoder(16#e5#)) OR
 					(reg_q779 AND symb_decoder(16#9f#)) OR
 					(reg_q779 AND symb_decoder(16#99#)) OR
 					(reg_q779 AND symb_decoder(16#61#)) OR
 					(reg_q779 AND symb_decoder(16#bb#)) OR
 					(reg_q779 AND symb_decoder(16#7a#)) OR
 					(reg_q779 AND symb_decoder(16#ad#)) OR
 					(reg_q779 AND symb_decoder(16#d4#)) OR
 					(reg_q779 AND symb_decoder(16#57#)) OR
 					(reg_q779 AND symb_decoder(16#c9#)) OR
 					(reg_q779 AND symb_decoder(16#d9#)) OR
 					(reg_q779 AND symb_decoder(16#e8#)) OR
 					(reg_q779 AND symb_decoder(16#f7#)) OR
 					(reg_q779 AND symb_decoder(16#44#)) OR
 					(reg_q779 AND symb_decoder(16#62#)) OR
 					(reg_q779 AND symb_decoder(16#d2#)) OR
 					(reg_q779 AND symb_decoder(16#95#)) OR
 					(reg_q779 AND symb_decoder(16#13#)) OR
 					(reg_q779 AND symb_decoder(16#a8#)) OR
 					(reg_q779 AND symb_decoder(16#3a#)) OR
 					(reg_q779 AND symb_decoder(16#96#)) OR
 					(reg_q779 AND symb_decoder(16#3f#)) OR
 					(reg_q779 AND symb_decoder(16#4b#)) OR
 					(reg_q779 AND symb_decoder(16#8f#)) OR
 					(reg_q779 AND symb_decoder(16#33#)) OR
 					(reg_q779 AND symb_decoder(16#5f#)) OR
 					(reg_q779 AND symb_decoder(16#a4#)) OR
 					(reg_q779 AND symb_decoder(16#ac#)) OR
 					(reg_q779 AND symb_decoder(16#14#)) OR
 					(reg_q779 AND symb_decoder(16#65#)) OR
 					(reg_q779 AND symb_decoder(16#7e#)) OR
 					(reg_q779 AND symb_decoder(16#1c#)) OR
 					(reg_q779 AND symb_decoder(16#79#)) OR
 					(reg_q779 AND symb_decoder(16#93#)) OR
 					(reg_q779 AND symb_decoder(16#b9#)) OR
 					(reg_q779 AND symb_decoder(16#2f#)) OR
 					(reg_q779 AND symb_decoder(16#0f#)) OR
 					(reg_q779 AND symb_decoder(16#98#)) OR
 					(reg_q779 AND symb_decoder(16#21#)) OR
 					(reg_q779 AND symb_decoder(16#92#)) OR
 					(reg_q779 AND symb_decoder(16#f0#)) OR
 					(reg_q779 AND symb_decoder(16#2b#)) OR
 					(reg_q779 AND symb_decoder(16#71#)) OR
 					(reg_q779 AND symb_decoder(16#c7#)) OR
 					(reg_q779 AND symb_decoder(16#f5#)) OR
 					(reg_q779 AND symb_decoder(16#de#)) OR
 					(reg_q779 AND symb_decoder(16#83#)) OR
 					(reg_q779 AND symb_decoder(16#be#)) OR
 					(reg_q779 AND symb_decoder(16#b0#)) OR
 					(reg_q779 AND symb_decoder(16#91#)) OR
 					(reg_q779 AND symb_decoder(16#29#)) OR
 					(reg_q779 AND symb_decoder(16#fb#)) OR
 					(reg_q779 AND symb_decoder(16#6f#)) OR
 					(reg_q779 AND symb_decoder(16#52#)) OR
 					(reg_q779 AND symb_decoder(16#56#)) OR
 					(reg_q779 AND symb_decoder(16#2e#)) OR
 					(reg_q779 AND symb_decoder(16#03#)) OR
 					(reg_q779 AND symb_decoder(16#11#));
reg_q779_init <= '0' ;
	p_reg_q779: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q779 <= reg_q779_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q779 <= reg_q779_init;
        else
          reg_q779 <= reg_q779_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2124_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2124 AND symb_decoder(16#9f#)) OR
 					(reg_q2124 AND symb_decoder(16#52#)) OR
 					(reg_q2124 AND symb_decoder(16#c5#)) OR
 					(reg_q2124 AND symb_decoder(16#c6#)) OR
 					(reg_q2124 AND symb_decoder(16#14#)) OR
 					(reg_q2124 AND symb_decoder(16#24#)) OR
 					(reg_q2124 AND symb_decoder(16#99#)) OR
 					(reg_q2124 AND symb_decoder(16#0f#)) OR
 					(reg_q2124 AND symb_decoder(16#86#)) OR
 					(reg_q2124 AND symb_decoder(16#8e#)) OR
 					(reg_q2124 AND symb_decoder(16#7f#)) OR
 					(reg_q2124 AND symb_decoder(16#75#)) OR
 					(reg_q2124 AND symb_decoder(16#cc#)) OR
 					(reg_q2124 AND symb_decoder(16#b4#)) OR
 					(reg_q2124 AND symb_decoder(16#9a#)) OR
 					(reg_q2124 AND symb_decoder(16#03#)) OR
 					(reg_q2124 AND symb_decoder(16#f8#)) OR
 					(reg_q2124 AND symb_decoder(16#31#)) OR
 					(reg_q2124 AND symb_decoder(16#95#)) OR
 					(reg_q2124 AND symb_decoder(16#c0#)) OR
 					(reg_q2124 AND symb_decoder(16#89#)) OR
 					(reg_q2124 AND symb_decoder(16#42#)) OR
 					(reg_q2124 AND symb_decoder(16#8b#)) OR
 					(reg_q2124 AND symb_decoder(16#59#)) OR
 					(reg_q2124 AND symb_decoder(16#07#)) OR
 					(reg_q2124 AND symb_decoder(16#a2#)) OR
 					(reg_q2124 AND symb_decoder(16#6e#)) OR
 					(reg_q2124 AND symb_decoder(16#10#)) OR
 					(reg_q2124 AND symb_decoder(16#58#)) OR
 					(reg_q2124 AND symb_decoder(16#5c#)) OR
 					(reg_q2124 AND symb_decoder(16#5b#)) OR
 					(reg_q2124 AND symb_decoder(16#20#)) OR
 					(reg_q2124 AND symb_decoder(16#00#)) OR
 					(reg_q2124 AND symb_decoder(16#bf#)) OR
 					(reg_q2124 AND symb_decoder(16#cf#)) OR
 					(reg_q2124 AND symb_decoder(16#98#)) OR
 					(reg_q2124 AND symb_decoder(16#90#)) OR
 					(reg_q2124 AND symb_decoder(16#1a#)) OR
 					(reg_q2124 AND symb_decoder(16#26#)) OR
 					(reg_q2124 AND symb_decoder(16#a5#)) OR
 					(reg_q2124 AND symb_decoder(16#7b#)) OR
 					(reg_q2124 AND symb_decoder(16#60#)) OR
 					(reg_q2124 AND symb_decoder(16#6b#)) OR
 					(reg_q2124 AND symb_decoder(16#87#)) OR
 					(reg_q2124 AND symb_decoder(16#ae#)) OR
 					(reg_q2124 AND symb_decoder(16#56#)) OR
 					(reg_q2124 AND symb_decoder(16#0b#)) OR
 					(reg_q2124 AND symb_decoder(16#04#)) OR
 					(reg_q2124 AND symb_decoder(16#c3#)) OR
 					(reg_q2124 AND symb_decoder(16#2c#)) OR
 					(reg_q2124 AND symb_decoder(16#1b#)) OR
 					(reg_q2124 AND symb_decoder(16#b8#)) OR
 					(reg_q2124 AND symb_decoder(16#09#)) OR
 					(reg_q2124 AND symb_decoder(16#aa#)) OR
 					(reg_q2124 AND symb_decoder(16#12#)) OR
 					(reg_q2124 AND symb_decoder(16#b6#)) OR
 					(reg_q2124 AND symb_decoder(16#17#)) OR
 					(reg_q2124 AND symb_decoder(16#8d#)) OR
 					(reg_q2124 AND symb_decoder(16#18#)) OR
 					(reg_q2124 AND symb_decoder(16#57#)) OR
 					(reg_q2124 AND symb_decoder(16#16#)) OR
 					(reg_q2124 AND symb_decoder(16#3b#)) OR
 					(reg_q2124 AND symb_decoder(16#7e#)) OR
 					(reg_q2124 AND symb_decoder(16#a7#)) OR
 					(reg_q2124 AND symb_decoder(16#ee#)) OR
 					(reg_q2124 AND symb_decoder(16#de#)) OR
 					(reg_q2124 AND symb_decoder(16#93#)) OR
 					(reg_q2124 AND symb_decoder(16#d1#)) OR
 					(reg_q2124 AND symb_decoder(16#7a#)) OR
 					(reg_q2124 AND symb_decoder(16#c1#)) OR
 					(reg_q2124 AND symb_decoder(16#6a#)) OR
 					(reg_q2124 AND symb_decoder(16#db#)) OR
 					(reg_q2124 AND symb_decoder(16#92#)) OR
 					(reg_q2124 AND symb_decoder(16#71#)) OR
 					(reg_q2124 AND symb_decoder(16#0c#)) OR
 					(reg_q2124 AND symb_decoder(16#4e#)) OR
 					(reg_q2124 AND symb_decoder(16#f6#)) OR
 					(reg_q2124 AND symb_decoder(16#69#)) OR
 					(reg_q2124 AND symb_decoder(16#a0#)) OR
 					(reg_q2124 AND symb_decoder(16#b1#)) OR
 					(reg_q2124 AND symb_decoder(16#61#)) OR
 					(reg_q2124 AND symb_decoder(16#fd#)) OR
 					(reg_q2124 AND symb_decoder(16#9b#)) OR
 					(reg_q2124 AND symb_decoder(16#0e#)) OR
 					(reg_q2124 AND symb_decoder(16#c2#)) OR
 					(reg_q2124 AND symb_decoder(16#d9#)) OR
 					(reg_q2124 AND symb_decoder(16#5d#)) OR
 					(reg_q2124 AND symb_decoder(16#cb#)) OR
 					(reg_q2124 AND symb_decoder(16#19#)) OR
 					(reg_q2124 AND symb_decoder(16#30#)) OR
 					(reg_q2124 AND symb_decoder(16#84#)) OR
 					(reg_q2124 AND symb_decoder(16#9e#)) OR
 					(reg_q2124 AND symb_decoder(16#54#)) OR
 					(reg_q2124 AND symb_decoder(16#a3#)) OR
 					(reg_q2124 AND symb_decoder(16#bb#)) OR
 					(reg_q2124 AND symb_decoder(16#50#)) OR
 					(reg_q2124 AND symb_decoder(16#13#)) OR
 					(reg_q2124 AND symb_decoder(16#ca#)) OR
 					(reg_q2124 AND symb_decoder(16#b5#)) OR
 					(reg_q2124 AND symb_decoder(16#9d#)) OR
 					(reg_q2124 AND symb_decoder(16#ad#)) OR
 					(reg_q2124 AND symb_decoder(16#d6#)) OR
 					(reg_q2124 AND symb_decoder(16#a1#)) OR
 					(reg_q2124 AND symb_decoder(16#63#)) OR
 					(reg_q2124 AND symb_decoder(16#88#)) OR
 					(reg_q2124 AND symb_decoder(16#70#)) OR
 					(reg_q2124 AND symb_decoder(16#7d#)) OR
 					(reg_q2124 AND symb_decoder(16#37#)) OR
 					(reg_q2124 AND symb_decoder(16#72#)) OR
 					(reg_q2124 AND symb_decoder(16#5e#)) OR
 					(reg_q2124 AND symb_decoder(16#28#)) OR
 					(reg_q2124 AND symb_decoder(16#29#)) OR
 					(reg_q2124 AND symb_decoder(16#96#)) OR
 					(reg_q2124 AND symb_decoder(16#38#)) OR
 					(reg_q2124 AND symb_decoder(16#f9#)) OR
 					(reg_q2124 AND symb_decoder(16#ff#)) OR
 					(reg_q2124 AND symb_decoder(16#66#)) OR
 					(reg_q2124 AND symb_decoder(16#c4#)) OR
 					(reg_q2124 AND symb_decoder(16#45#)) OR
 					(reg_q2124 AND symb_decoder(16#2f#)) OR
 					(reg_q2124 AND symb_decoder(16#67#)) OR
 					(reg_q2124 AND symb_decoder(16#33#)) OR
 					(reg_q2124 AND symb_decoder(16#46#)) OR
 					(reg_q2124 AND symb_decoder(16#0d#)) OR
 					(reg_q2124 AND symb_decoder(16#f5#)) OR
 					(reg_q2124 AND symb_decoder(16#41#)) OR
 					(reg_q2124 AND symb_decoder(16#73#)) OR
 					(reg_q2124 AND symb_decoder(16#32#)) OR
 					(reg_q2124 AND symb_decoder(16#3e#)) OR
 					(reg_q2124 AND symb_decoder(16#80#)) OR
 					(reg_q2124 AND symb_decoder(16#ed#)) OR
 					(reg_q2124 AND symb_decoder(16#d3#)) OR
 					(reg_q2124 AND symb_decoder(16#b7#)) OR
 					(reg_q2124 AND symb_decoder(16#b9#)) OR
 					(reg_q2124 AND symb_decoder(16#ac#)) OR
 					(reg_q2124 AND symb_decoder(16#2e#)) OR
 					(reg_q2124 AND symb_decoder(16#eb#)) OR
 					(reg_q2124 AND symb_decoder(16#0a#)) OR
 					(reg_q2124 AND symb_decoder(16#7c#)) OR
 					(reg_q2124 AND symb_decoder(16#76#)) OR
 					(reg_q2124 AND symb_decoder(16#47#)) OR
 					(reg_q2124 AND symb_decoder(16#74#)) OR
 					(reg_q2124 AND symb_decoder(16#cd#)) OR
 					(reg_q2124 AND symb_decoder(16#f0#)) OR
 					(reg_q2124 AND symb_decoder(16#f7#)) OR
 					(reg_q2124 AND symb_decoder(16#64#)) OR
 					(reg_q2124 AND symb_decoder(16#a6#)) OR
 					(reg_q2124 AND symb_decoder(16#bd#)) OR
 					(reg_q2124 AND symb_decoder(16#82#)) OR
 					(reg_q2124 AND symb_decoder(16#85#)) OR
 					(reg_q2124 AND symb_decoder(16#53#)) OR
 					(reg_q2124 AND symb_decoder(16#4b#)) OR
 					(reg_q2124 AND symb_decoder(16#3d#)) OR
 					(reg_q2124 AND symb_decoder(16#c7#)) OR
 					(reg_q2124 AND symb_decoder(16#34#)) OR
 					(reg_q2124 AND symb_decoder(16#ec#)) OR
 					(reg_q2124 AND symb_decoder(16#4c#)) OR
 					(reg_q2124 AND symb_decoder(16#e9#)) OR
 					(reg_q2124 AND symb_decoder(16#e5#)) OR
 					(reg_q2124 AND symb_decoder(16#02#)) OR
 					(reg_q2124 AND symb_decoder(16#d0#)) OR
 					(reg_q2124 AND symb_decoder(16#d4#)) OR
 					(reg_q2124 AND symb_decoder(16#51#)) OR
 					(reg_q2124 AND symb_decoder(16#2a#)) OR
 					(reg_q2124 AND symb_decoder(16#1e#)) OR
 					(reg_q2124 AND symb_decoder(16#4a#)) OR
 					(reg_q2124 AND symb_decoder(16#fb#)) OR
 					(reg_q2124 AND symb_decoder(16#22#)) OR
 					(reg_q2124 AND symb_decoder(16#44#)) OR
 					(reg_q2124 AND symb_decoder(16#fa#)) OR
 					(reg_q2124 AND symb_decoder(16#21#)) OR
 					(reg_q2124 AND symb_decoder(16#be#)) OR
 					(reg_q2124 AND symb_decoder(16#2b#)) OR
 					(reg_q2124 AND symb_decoder(16#e7#)) OR
 					(reg_q2124 AND symb_decoder(16#a8#)) OR
 					(reg_q2124 AND symb_decoder(16#43#)) OR
 					(reg_q2124 AND symb_decoder(16#fc#)) OR
 					(reg_q2124 AND symb_decoder(16#4d#)) OR
 					(reg_q2124 AND symb_decoder(16#d2#)) OR
 					(reg_q2124 AND symb_decoder(16#c8#)) OR
 					(reg_q2124 AND symb_decoder(16#ba#)) OR
 					(reg_q2124 AND symb_decoder(16#e8#)) OR
 					(reg_q2124 AND symb_decoder(16#e2#)) OR
 					(reg_q2124 AND symb_decoder(16#fe#)) OR
 					(reg_q2124 AND symb_decoder(16#39#)) OR
 					(reg_q2124 AND symb_decoder(16#9c#)) OR
 					(reg_q2124 AND symb_decoder(16#65#)) OR
 					(reg_q2124 AND symb_decoder(16#35#)) OR
 					(reg_q2124 AND symb_decoder(16#36#)) OR
 					(reg_q2124 AND symb_decoder(16#15#)) OR
 					(reg_q2124 AND symb_decoder(16#94#)) OR
 					(reg_q2124 AND symb_decoder(16#05#)) OR
 					(reg_q2124 AND symb_decoder(16#b0#)) OR
 					(reg_q2124 AND symb_decoder(16#97#)) OR
 					(reg_q2124 AND symb_decoder(16#dc#)) OR
 					(reg_q2124 AND symb_decoder(16#e4#)) OR
 					(reg_q2124 AND symb_decoder(16#08#)) OR
 					(reg_q2124 AND symb_decoder(16#3a#)) OR
 					(reg_q2124 AND symb_decoder(16#b2#)) OR
 					(reg_q2124 AND symb_decoder(16#40#)) OR
 					(reg_q2124 AND symb_decoder(16#ab#)) OR
 					(reg_q2124 AND symb_decoder(16#77#)) OR
 					(reg_q2124 AND symb_decoder(16#ef#)) OR
 					(reg_q2124 AND symb_decoder(16#68#)) OR
 					(reg_q2124 AND symb_decoder(16#81#)) OR
 					(reg_q2124 AND symb_decoder(16#91#)) OR
 					(reg_q2124 AND symb_decoder(16#79#)) OR
 					(reg_q2124 AND symb_decoder(16#a4#)) OR
 					(reg_q2124 AND symb_decoder(16#11#)) OR
 					(reg_q2124 AND symb_decoder(16#c9#)) OR
 					(reg_q2124 AND symb_decoder(16#d7#)) OR
 					(reg_q2124 AND symb_decoder(16#1d#)) OR
 					(reg_q2124 AND symb_decoder(16#5a#)) OR
 					(reg_q2124 AND symb_decoder(16#3c#)) OR
 					(reg_q2124 AND symb_decoder(16#48#)) OR
 					(reg_q2124 AND symb_decoder(16#e1#)) OR
 					(reg_q2124 AND symb_decoder(16#e6#)) OR
 					(reg_q2124 AND symb_decoder(16#8f#)) OR
 					(reg_q2124 AND symb_decoder(16#1c#)) OR
 					(reg_q2124 AND symb_decoder(16#4f#)) OR
 					(reg_q2124 AND symb_decoder(16#ce#)) OR
 					(reg_q2124 AND symb_decoder(16#8a#)) OR
 					(reg_q2124 AND symb_decoder(16#a9#)) OR
 					(reg_q2124 AND symb_decoder(16#1f#)) OR
 					(reg_q2124 AND symb_decoder(16#d8#)) OR
 					(reg_q2124 AND symb_decoder(16#2d#)) OR
 					(reg_q2124 AND symb_decoder(16#01#)) OR
 					(reg_q2124 AND symb_decoder(16#df#)) OR
 					(reg_q2124 AND symb_decoder(16#dd#)) OR
 					(reg_q2124 AND symb_decoder(16#f2#)) OR
 					(reg_q2124 AND symb_decoder(16#3f#)) OR
 					(reg_q2124 AND symb_decoder(16#62#)) OR
 					(reg_q2124 AND symb_decoder(16#da#)) OR
 					(reg_q2124 AND symb_decoder(16#06#)) OR
 					(reg_q2124 AND symb_decoder(16#49#)) OR
 					(reg_q2124 AND symb_decoder(16#55#)) OR
 					(reg_q2124 AND symb_decoder(16#6d#)) OR
 					(reg_q2124 AND symb_decoder(16#ea#)) OR
 					(reg_q2124 AND symb_decoder(16#e0#)) OR
 					(reg_q2124 AND symb_decoder(16#f4#)) OR
 					(reg_q2124 AND symb_decoder(16#8c#)) OR
 					(reg_q2124 AND symb_decoder(16#25#)) OR
 					(reg_q2124 AND symb_decoder(16#e3#)) OR
 					(reg_q2124 AND symb_decoder(16#78#)) OR
 					(reg_q2124 AND symb_decoder(16#27#)) OR
 					(reg_q2124 AND symb_decoder(16#6c#)) OR
 					(reg_q2124 AND symb_decoder(16#f3#)) OR
 					(reg_q2124 AND symb_decoder(16#af#)) OR
 					(reg_q2124 AND symb_decoder(16#6f#)) OR
 					(reg_q2124 AND symb_decoder(16#83#)) OR
 					(reg_q2124 AND symb_decoder(16#5f#)) OR
 					(reg_q2124 AND symb_decoder(16#bc#)) OR
 					(reg_q2124 AND symb_decoder(16#f1#)) OR
 					(reg_q2124 AND symb_decoder(16#b3#)) OR
 					(reg_q2124 AND symb_decoder(16#d5#)) OR
 					(reg_q2124 AND symb_decoder(16#23#));
reg_q2124_init <= '0' ;
	p_reg_q2124: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2124 <= reg_q2124_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2124 <= reg_q2124_init;
        else
          reg_q2124 <= reg_q2124_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q665_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q665 AND symb_decoder(16#2e#)) OR
 					(reg_q665 AND symb_decoder(16#24#)) OR
 					(reg_q665 AND symb_decoder(16#37#)) OR
 					(reg_q665 AND symb_decoder(16#cb#)) OR
 					(reg_q665 AND symb_decoder(16#c8#)) OR
 					(reg_q665 AND symb_decoder(16#0b#)) OR
 					(reg_q665 AND symb_decoder(16#d0#)) OR
 					(reg_q665 AND symb_decoder(16#6d#)) OR
 					(reg_q665 AND symb_decoder(16#cc#)) OR
 					(reg_q665 AND symb_decoder(16#89#)) OR
 					(reg_q665 AND symb_decoder(16#be#)) OR
 					(reg_q665 AND symb_decoder(16#ca#)) OR
 					(reg_q665 AND symb_decoder(16#fd#)) OR
 					(reg_q665 AND symb_decoder(16#d8#)) OR
 					(reg_q665 AND symb_decoder(16#ae#)) OR
 					(reg_q665 AND symb_decoder(16#5b#)) OR
 					(reg_q665 AND symb_decoder(16#b4#)) OR
 					(reg_q665 AND symb_decoder(16#57#)) OR
 					(reg_q665 AND symb_decoder(16#d1#)) OR
 					(reg_q665 AND symb_decoder(16#9e#)) OR
 					(reg_q665 AND symb_decoder(16#b2#)) OR
 					(reg_q665 AND symb_decoder(16#75#)) OR
 					(reg_q665 AND symb_decoder(16#e8#)) OR
 					(reg_q665 AND symb_decoder(16#6c#)) OR
 					(reg_q665 AND symb_decoder(16#3d#)) OR
 					(reg_q665 AND symb_decoder(16#25#)) OR
 					(reg_q665 AND symb_decoder(16#f5#)) OR
 					(reg_q665 AND symb_decoder(16#f7#)) OR
 					(reg_q665 AND symb_decoder(16#98#)) OR
 					(reg_q665 AND symb_decoder(16#ef#)) OR
 					(reg_q665 AND symb_decoder(16#19#)) OR
 					(reg_q665 AND symb_decoder(16#c0#)) OR
 					(reg_q665 AND symb_decoder(16#86#)) OR
 					(reg_q665 AND symb_decoder(16#d3#)) OR
 					(reg_q665 AND symb_decoder(16#d4#)) OR
 					(reg_q665 AND symb_decoder(16#dc#)) OR
 					(reg_q665 AND symb_decoder(16#8d#)) OR
 					(reg_q665 AND symb_decoder(16#9b#)) OR
 					(reg_q665 AND symb_decoder(16#32#)) OR
 					(reg_q665 AND symb_decoder(16#77#)) OR
 					(reg_q665 AND symb_decoder(16#bc#)) OR
 					(reg_q665 AND symb_decoder(16#a1#)) OR
 					(reg_q665 AND symb_decoder(16#90#)) OR
 					(reg_q665 AND symb_decoder(16#91#)) OR
 					(reg_q665 AND symb_decoder(16#f3#)) OR
 					(reg_q665 AND symb_decoder(16#79#)) OR
 					(reg_q665 AND symb_decoder(16#eb#)) OR
 					(reg_q665 AND symb_decoder(16#bf#)) OR
 					(reg_q665 AND symb_decoder(16#44#)) OR
 					(reg_q665 AND symb_decoder(16#e9#)) OR
 					(reg_q665 AND symb_decoder(16#d7#)) OR
 					(reg_q665 AND symb_decoder(16#40#)) OR
 					(reg_q665 AND symb_decoder(16#95#)) OR
 					(reg_q665 AND symb_decoder(16#2f#)) OR
 					(reg_q665 AND symb_decoder(16#7d#)) OR
 					(reg_q665 AND symb_decoder(16#ec#)) OR
 					(reg_q665 AND symb_decoder(16#f4#)) OR
 					(reg_q665 AND symb_decoder(16#cf#)) OR
 					(reg_q665 AND symb_decoder(16#3b#)) OR
 					(reg_q665 AND symb_decoder(16#4b#)) OR
 					(reg_q665 AND symb_decoder(16#3e#)) OR
 					(reg_q665 AND symb_decoder(16#5e#)) OR
 					(reg_q665 AND symb_decoder(16#7a#)) OR
 					(reg_q665 AND symb_decoder(16#01#)) OR
 					(reg_q665 AND symb_decoder(16#36#)) OR
 					(reg_q665 AND symb_decoder(16#38#)) OR
 					(reg_q665 AND symb_decoder(16#b0#)) OR
 					(reg_q665 AND symb_decoder(16#15#)) OR
 					(reg_q665 AND symb_decoder(16#0f#)) OR
 					(reg_q665 AND symb_decoder(16#b3#)) OR
 					(reg_q665 AND symb_decoder(16#97#)) OR
 					(reg_q665 AND symb_decoder(16#6b#)) OR
 					(reg_q665 AND symb_decoder(16#1a#)) OR
 					(reg_q665 AND symb_decoder(16#54#)) OR
 					(reg_q665 AND symb_decoder(16#0a#)) OR
 					(reg_q665 AND symb_decoder(16#ea#)) OR
 					(reg_q665 AND symb_decoder(16#03#)) OR
 					(reg_q665 AND symb_decoder(16#74#)) OR
 					(reg_q665 AND symb_decoder(16#72#)) OR
 					(reg_q665 AND symb_decoder(16#18#)) OR
 					(reg_q665 AND symb_decoder(16#2a#)) OR
 					(reg_q665 AND symb_decoder(16#60#)) OR
 					(reg_q665 AND symb_decoder(16#c6#)) OR
 					(reg_q665 AND symb_decoder(16#6a#)) OR
 					(reg_q665 AND symb_decoder(16#8a#)) OR
 					(reg_q665 AND symb_decoder(16#17#)) OR
 					(reg_q665 AND symb_decoder(16#e5#)) OR
 					(reg_q665 AND symb_decoder(16#a9#)) OR
 					(reg_q665 AND symb_decoder(16#12#)) OR
 					(reg_q665 AND symb_decoder(16#5c#)) OR
 					(reg_q665 AND symb_decoder(16#82#)) OR
 					(reg_q665 AND symb_decoder(16#14#)) OR
 					(reg_q665 AND symb_decoder(16#ac#)) OR
 					(reg_q665 AND symb_decoder(16#31#)) OR
 					(reg_q665 AND symb_decoder(16#51#)) OR
 					(reg_q665 AND symb_decoder(16#1c#)) OR
 					(reg_q665 AND symb_decoder(16#87#)) OR
 					(reg_q665 AND symb_decoder(16#b9#)) OR
 					(reg_q665 AND symb_decoder(16#06#)) OR
 					(reg_q665 AND symb_decoder(16#35#)) OR
 					(reg_q665 AND symb_decoder(16#d9#)) OR
 					(reg_q665 AND symb_decoder(16#2c#)) OR
 					(reg_q665 AND symb_decoder(16#b6#)) OR
 					(reg_q665 AND symb_decoder(16#1f#)) OR
 					(reg_q665 AND symb_decoder(16#ba#)) OR
 					(reg_q665 AND symb_decoder(16#00#)) OR
 					(reg_q665 AND symb_decoder(16#c9#)) OR
 					(reg_q665 AND symb_decoder(16#df#)) OR
 					(reg_q665 AND symb_decoder(16#7b#)) OR
 					(reg_q665 AND symb_decoder(16#a0#)) OR
 					(reg_q665 AND symb_decoder(16#1b#)) OR
 					(reg_q665 AND symb_decoder(16#64#)) OR
 					(reg_q665 AND symb_decoder(16#73#)) OR
 					(reg_q665 AND symb_decoder(16#f9#)) OR
 					(reg_q665 AND symb_decoder(16#b8#)) OR
 					(reg_q665 AND symb_decoder(16#9d#)) OR
 					(reg_q665 AND symb_decoder(16#af#)) OR
 					(reg_q665 AND symb_decoder(16#9f#)) OR
 					(reg_q665 AND symb_decoder(16#8c#)) OR
 					(reg_q665 AND symb_decoder(16#22#)) OR
 					(reg_q665 AND symb_decoder(16#0d#)) OR
 					(reg_q665 AND symb_decoder(16#05#)) OR
 					(reg_q665 AND symb_decoder(16#2b#)) OR
 					(reg_q665 AND symb_decoder(16#21#)) OR
 					(reg_q665 AND symb_decoder(16#5d#)) OR
 					(reg_q665 AND symb_decoder(16#8b#)) OR
 					(reg_q665 AND symb_decoder(16#78#)) OR
 					(reg_q665 AND symb_decoder(16#26#)) OR
 					(reg_q665 AND symb_decoder(16#96#)) OR
 					(reg_q665 AND symb_decoder(16#63#)) OR
 					(reg_q665 AND symb_decoder(16#71#)) OR
 					(reg_q665 AND symb_decoder(16#7e#)) OR
 					(reg_q665 AND symb_decoder(16#41#)) OR
 					(reg_q665 AND symb_decoder(16#76#)) OR
 					(reg_q665 AND symb_decoder(16#93#)) OR
 					(reg_q665 AND symb_decoder(16#80#)) OR
 					(reg_q665 AND symb_decoder(16#a5#)) OR
 					(reg_q665 AND symb_decoder(16#59#)) OR
 					(reg_q665 AND symb_decoder(16#c2#)) OR
 					(reg_q665 AND symb_decoder(16#2d#)) OR
 					(reg_q665 AND symb_decoder(16#67#)) OR
 					(reg_q665 AND symb_decoder(16#d5#)) OR
 					(reg_q665 AND symb_decoder(16#7f#)) OR
 					(reg_q665 AND symb_decoder(16#3c#)) OR
 					(reg_q665 AND symb_decoder(16#5f#)) OR
 					(reg_q665 AND symb_decoder(16#48#)) OR
 					(reg_q665 AND symb_decoder(16#e6#)) OR
 					(reg_q665 AND symb_decoder(16#13#)) OR
 					(reg_q665 AND symb_decoder(16#ff#)) OR
 					(reg_q665 AND symb_decoder(16#66#)) OR
 					(reg_q665 AND symb_decoder(16#8f#)) OR
 					(reg_q665 AND symb_decoder(16#c7#)) OR
 					(reg_q665 AND symb_decoder(16#b1#)) OR
 					(reg_q665 AND symb_decoder(16#04#)) OR
 					(reg_q665 AND symb_decoder(16#fc#)) OR
 					(reg_q665 AND symb_decoder(16#ab#)) OR
 					(reg_q665 AND symb_decoder(16#fb#)) OR
 					(reg_q665 AND symb_decoder(16#92#)) OR
 					(reg_q665 AND symb_decoder(16#4d#)) OR
 					(reg_q665 AND symb_decoder(16#94#)) OR
 					(reg_q665 AND symb_decoder(16#65#)) OR
 					(reg_q665 AND symb_decoder(16#f1#)) OR
 					(reg_q665 AND symb_decoder(16#0c#)) OR
 					(reg_q665 AND symb_decoder(16#45#)) OR
 					(reg_q665 AND symb_decoder(16#85#)) OR
 					(reg_q665 AND symb_decoder(16#e3#)) OR
 					(reg_q665 AND symb_decoder(16#3a#)) OR
 					(reg_q665 AND symb_decoder(16#34#)) OR
 					(reg_q665 AND symb_decoder(16#39#)) OR
 					(reg_q665 AND symb_decoder(16#e1#)) OR
 					(reg_q665 AND symb_decoder(16#3f#)) OR
 					(reg_q665 AND symb_decoder(16#e7#)) OR
 					(reg_q665 AND symb_decoder(16#99#)) OR
 					(reg_q665 AND symb_decoder(16#81#)) OR
 					(reg_q665 AND symb_decoder(16#62#)) OR
 					(reg_q665 AND symb_decoder(16#bb#)) OR
 					(reg_q665 AND symb_decoder(16#a2#)) OR
 					(reg_q665 AND symb_decoder(16#30#)) OR
 					(reg_q665 AND symb_decoder(16#a4#)) OR
 					(reg_q665 AND symb_decoder(16#33#)) OR
 					(reg_q665 AND symb_decoder(16#b5#)) OR
 					(reg_q665 AND symb_decoder(16#f2#)) OR
 					(reg_q665 AND symb_decoder(16#a6#)) OR
 					(reg_q665 AND symb_decoder(16#43#)) OR
 					(reg_q665 AND symb_decoder(16#f8#)) OR
 					(reg_q665 AND symb_decoder(16#27#)) OR
 					(reg_q665 AND symb_decoder(16#e4#)) OR
 					(reg_q665 AND symb_decoder(16#cd#)) OR
 					(reg_q665 AND symb_decoder(16#07#)) OR
 					(reg_q665 AND symb_decoder(16#55#)) OR
 					(reg_q665 AND symb_decoder(16#c1#)) OR
 					(reg_q665 AND symb_decoder(16#d2#)) OR
 					(reg_q665 AND symb_decoder(16#ce#)) OR
 					(reg_q665 AND symb_decoder(16#4f#)) OR
 					(reg_q665 AND symb_decoder(16#0e#)) OR
 					(reg_q665 AND symb_decoder(16#a8#)) OR
 					(reg_q665 AND symb_decoder(16#61#)) OR
 					(reg_q665 AND symb_decoder(16#f0#)) OR
 					(reg_q665 AND symb_decoder(16#20#)) OR
 					(reg_q665 AND symb_decoder(16#84#)) OR
 					(reg_q665 AND symb_decoder(16#c5#)) OR
 					(reg_q665 AND symb_decoder(16#53#)) OR
 					(reg_q665 AND symb_decoder(16#29#)) OR
 					(reg_q665 AND symb_decoder(16#23#)) OR
 					(reg_q665 AND symb_decoder(16#1d#)) OR
 					(reg_q665 AND symb_decoder(16#bd#)) OR
 					(reg_q665 AND symb_decoder(16#a3#)) OR
 					(reg_q665 AND symb_decoder(16#52#)) OR
 					(reg_q665 AND symb_decoder(16#ee#)) OR
 					(reg_q665 AND symb_decoder(16#4c#)) OR
 					(reg_q665 AND symb_decoder(16#fe#)) OR
 					(reg_q665 AND symb_decoder(16#fa#)) OR
 					(reg_q665 AND symb_decoder(16#9a#)) OR
 					(reg_q665 AND symb_decoder(16#da#)) OR
 					(reg_q665 AND symb_decoder(16#d6#)) OR
 					(reg_q665 AND symb_decoder(16#db#)) OR
 					(reg_q665 AND symb_decoder(16#a7#)) OR
 					(reg_q665 AND symb_decoder(16#f6#)) OR
 					(reg_q665 AND symb_decoder(16#dd#)) OR
 					(reg_q665 AND symb_decoder(16#83#)) OR
 					(reg_q665 AND symb_decoder(16#5a#)) OR
 					(reg_q665 AND symb_decoder(16#28#)) OR
 					(reg_q665 AND symb_decoder(16#58#)) OR
 					(reg_q665 AND symb_decoder(16#88#)) OR
 					(reg_q665 AND symb_decoder(16#ad#)) OR
 					(reg_q665 AND symb_decoder(16#ed#)) OR
 					(reg_q665 AND symb_decoder(16#42#)) OR
 					(reg_q665 AND symb_decoder(16#4a#)) OR
 					(reg_q665 AND symb_decoder(16#e2#)) OR
 					(reg_q665 AND symb_decoder(16#11#)) OR
 					(reg_q665 AND symb_decoder(16#9c#)) OR
 					(reg_q665 AND symb_decoder(16#68#)) OR
 					(reg_q665 AND symb_decoder(16#c3#)) OR
 					(reg_q665 AND symb_decoder(16#b7#)) OR
 					(reg_q665 AND symb_decoder(16#6e#)) OR
 					(reg_q665 AND symb_decoder(16#69#)) OR
 					(reg_q665 AND symb_decoder(16#47#)) OR
 					(reg_q665 AND symb_decoder(16#aa#)) OR
 					(reg_q665 AND symb_decoder(16#16#)) OR
 					(reg_q665 AND symb_decoder(16#7c#)) OR
 					(reg_q665 AND symb_decoder(16#46#)) OR
 					(reg_q665 AND symb_decoder(16#10#)) OR
 					(reg_q665 AND symb_decoder(16#56#)) OR
 					(reg_q665 AND symb_decoder(16#09#)) OR
 					(reg_q665 AND symb_decoder(16#08#)) OR
 					(reg_q665 AND symb_decoder(16#49#)) OR
 					(reg_q665 AND symb_decoder(16#02#)) OR
 					(reg_q665 AND symb_decoder(16#8e#)) OR
 					(reg_q665 AND symb_decoder(16#de#)) OR
 					(reg_q665 AND symb_decoder(16#e0#)) OR
 					(reg_q665 AND symb_decoder(16#1e#)) OR
 					(reg_q665 AND symb_decoder(16#50#)) OR
 					(reg_q665 AND symb_decoder(16#70#)) OR
 					(reg_q665 AND symb_decoder(16#c4#)) OR
 					(reg_q665 AND symb_decoder(16#4e#)) OR
 					(reg_q665 AND symb_decoder(16#6f#));
reg_q665_init <= '0' ;
	p_reg_q665: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q665 <= reg_q665_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q665 <= reg_q665_init;
        else
          reg_q665 <= reg_q665_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q816_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q816 AND symb_decoder(16#dc#)) OR
 					(reg_q816 AND symb_decoder(16#14#)) OR
 					(reg_q816 AND symb_decoder(16#08#)) OR
 					(reg_q816 AND symb_decoder(16#ea#)) OR
 					(reg_q816 AND symb_decoder(16#a2#)) OR
 					(reg_q816 AND symb_decoder(16#7b#)) OR
 					(reg_q816 AND symb_decoder(16#80#)) OR
 					(reg_q816 AND symb_decoder(16#70#)) OR
 					(reg_q816 AND symb_decoder(16#87#)) OR
 					(reg_q816 AND symb_decoder(16#28#)) OR
 					(reg_q816 AND symb_decoder(16#d7#)) OR
 					(reg_q816 AND symb_decoder(16#32#)) OR
 					(reg_q816 AND symb_decoder(16#81#)) OR
 					(reg_q816 AND symb_decoder(16#27#)) OR
 					(reg_q816 AND symb_decoder(16#fd#)) OR
 					(reg_q816 AND symb_decoder(16#74#)) OR
 					(reg_q816 AND symb_decoder(16#3b#)) OR
 					(reg_q816 AND symb_decoder(16#19#)) OR
 					(reg_q816 AND symb_decoder(16#9f#)) OR
 					(reg_q816 AND symb_decoder(16#91#)) OR
 					(reg_q816 AND symb_decoder(16#e7#)) OR
 					(reg_q816 AND symb_decoder(16#86#)) OR
 					(reg_q816 AND symb_decoder(16#4f#)) OR
 					(reg_q816 AND symb_decoder(16#65#)) OR
 					(reg_q816 AND symb_decoder(16#96#)) OR
 					(reg_q816 AND symb_decoder(16#ce#)) OR
 					(reg_q816 AND symb_decoder(16#1a#)) OR
 					(reg_q816 AND symb_decoder(16#9e#)) OR
 					(reg_q816 AND symb_decoder(16#ac#)) OR
 					(reg_q816 AND symb_decoder(16#9a#)) OR
 					(reg_q816 AND symb_decoder(16#b0#)) OR
 					(reg_q816 AND symb_decoder(16#cd#)) OR
 					(reg_q816 AND symb_decoder(16#6e#)) OR
 					(reg_q816 AND symb_decoder(16#64#)) OR
 					(reg_q816 AND symb_decoder(16#cc#)) OR
 					(reg_q816 AND symb_decoder(16#79#)) OR
 					(reg_q816 AND symb_decoder(16#d2#)) OR
 					(reg_q816 AND symb_decoder(16#e2#)) OR
 					(reg_q816 AND symb_decoder(16#dd#)) OR
 					(reg_q816 AND symb_decoder(16#2e#)) OR
 					(reg_q816 AND symb_decoder(16#35#)) OR
 					(reg_q816 AND symb_decoder(16#48#)) OR
 					(reg_q816 AND symb_decoder(16#5c#)) OR
 					(reg_q816 AND symb_decoder(16#4c#)) OR
 					(reg_q816 AND symb_decoder(16#c2#)) OR
 					(reg_q816 AND symb_decoder(16#95#)) OR
 					(reg_q816 AND symb_decoder(16#1c#)) OR
 					(reg_q816 AND symb_decoder(16#53#)) OR
 					(reg_q816 AND symb_decoder(16#6b#)) OR
 					(reg_q816 AND symb_decoder(16#d3#)) OR
 					(reg_q816 AND symb_decoder(16#c5#)) OR
 					(reg_q816 AND symb_decoder(16#b1#)) OR
 					(reg_q816 AND symb_decoder(16#58#)) OR
 					(reg_q816 AND symb_decoder(16#17#)) OR
 					(reg_q816 AND symb_decoder(16#f5#)) OR
 					(reg_q816 AND symb_decoder(16#bb#)) OR
 					(reg_q816 AND symb_decoder(16#ab#)) OR
 					(reg_q816 AND symb_decoder(16#fb#)) OR
 					(reg_q816 AND symb_decoder(16#88#)) OR
 					(reg_q816 AND symb_decoder(16#f7#)) OR
 					(reg_q816 AND symb_decoder(16#04#)) OR
 					(reg_q816 AND symb_decoder(16#9b#)) OR
 					(reg_q816 AND symb_decoder(16#5f#)) OR
 					(reg_q816 AND symb_decoder(16#b6#)) OR
 					(reg_q816 AND symb_decoder(16#b8#)) OR
 					(reg_q816 AND symb_decoder(16#fe#)) OR
 					(reg_q816 AND symb_decoder(16#8c#)) OR
 					(reg_q816 AND symb_decoder(16#db#)) OR
 					(reg_q816 AND symb_decoder(16#6c#)) OR
 					(reg_q816 AND symb_decoder(16#68#)) OR
 					(reg_q816 AND symb_decoder(16#1d#)) OR
 					(reg_q816 AND symb_decoder(16#11#)) OR
 					(reg_q816 AND symb_decoder(16#8a#)) OR
 					(reg_q816 AND symb_decoder(16#7c#)) OR
 					(reg_q816 AND symb_decoder(16#20#)) OR
 					(reg_q816 AND symb_decoder(16#44#)) OR
 					(reg_q816 AND symb_decoder(16#e8#)) OR
 					(reg_q816 AND symb_decoder(16#c9#)) OR
 					(reg_q816 AND symb_decoder(16#78#)) OR
 					(reg_q816 AND symb_decoder(16#83#)) OR
 					(reg_q816 AND symb_decoder(16#e6#)) OR
 					(reg_q816 AND symb_decoder(16#56#)) OR
 					(reg_q816 AND symb_decoder(16#73#)) OR
 					(reg_q816 AND symb_decoder(16#d9#)) OR
 					(reg_q816 AND symb_decoder(16#2c#)) OR
 					(reg_q816 AND symb_decoder(16#7e#)) OR
 					(reg_q816 AND symb_decoder(16#12#)) OR
 					(reg_q816 AND symb_decoder(16#69#)) OR
 					(reg_q816 AND symb_decoder(16#21#)) OR
 					(reg_q816 AND symb_decoder(16#84#)) OR
 					(reg_q816 AND symb_decoder(16#92#)) OR
 					(reg_q816 AND symb_decoder(16#1e#)) OR
 					(reg_q816 AND symb_decoder(16#ff#)) OR
 					(reg_q816 AND symb_decoder(16#ef#)) OR
 					(reg_q816 AND symb_decoder(16#43#)) OR
 					(reg_q816 AND symb_decoder(16#9c#)) OR
 					(reg_q816 AND symb_decoder(16#3e#)) OR
 					(reg_q816 AND symb_decoder(16#0b#)) OR
 					(reg_q816 AND symb_decoder(16#51#)) OR
 					(reg_q816 AND symb_decoder(16#0a#)) OR
 					(reg_q816 AND symb_decoder(16#f6#)) OR
 					(reg_q816 AND symb_decoder(16#ca#)) OR
 					(reg_q816 AND symb_decoder(16#41#)) OR
 					(reg_q816 AND symb_decoder(16#c0#)) OR
 					(reg_q816 AND symb_decoder(16#45#)) OR
 					(reg_q816 AND symb_decoder(16#a7#)) OR
 					(reg_q816 AND symb_decoder(16#9d#)) OR
 					(reg_q816 AND symb_decoder(16#f0#)) OR
 					(reg_q816 AND symb_decoder(16#f4#)) OR
 					(reg_q816 AND symb_decoder(16#07#)) OR
 					(reg_q816 AND symb_decoder(16#ba#)) OR
 					(reg_q816 AND symb_decoder(16#61#)) OR
 					(reg_q816 AND symb_decoder(16#ee#)) OR
 					(reg_q816 AND symb_decoder(16#89#)) OR
 					(reg_q816 AND symb_decoder(16#b2#)) OR
 					(reg_q816 AND symb_decoder(16#57#)) OR
 					(reg_q816 AND symb_decoder(16#2d#)) OR
 					(reg_q816 AND symb_decoder(16#df#)) OR
 					(reg_q816 AND symb_decoder(16#c1#)) OR
 					(reg_q816 AND symb_decoder(16#2b#)) OR
 					(reg_q816 AND symb_decoder(16#10#)) OR
 					(reg_q816 AND symb_decoder(16#77#)) OR
 					(reg_q816 AND symb_decoder(16#5e#)) OR
 					(reg_q816 AND symb_decoder(16#d8#)) OR
 					(reg_q816 AND symb_decoder(16#4a#)) OR
 					(reg_q816 AND symb_decoder(16#7a#)) OR
 					(reg_q816 AND symb_decoder(16#eb#)) OR
 					(reg_q816 AND symb_decoder(16#8f#)) OR
 					(reg_q816 AND symb_decoder(16#62#)) OR
 					(reg_q816 AND symb_decoder(16#60#)) OR
 					(reg_q816 AND symb_decoder(16#33#)) OR
 					(reg_q816 AND symb_decoder(16#54#)) OR
 					(reg_q816 AND symb_decoder(16#a4#)) OR
 					(reg_q816 AND symb_decoder(16#7d#)) OR
 					(reg_q816 AND symb_decoder(16#5a#)) OR
 					(reg_q816 AND symb_decoder(16#3d#)) OR
 					(reg_q816 AND symb_decoder(16#8e#)) OR
 					(reg_q816 AND symb_decoder(16#d6#)) OR
 					(reg_q816 AND symb_decoder(16#47#)) OR
 					(reg_q816 AND symb_decoder(16#15#)) OR
 					(reg_q816 AND symb_decoder(16#f2#)) OR
 					(reg_q816 AND symb_decoder(16#5b#)) OR
 					(reg_q816 AND symb_decoder(16#7f#)) OR
 					(reg_q816 AND symb_decoder(16#99#)) OR
 					(reg_q816 AND symb_decoder(16#e0#)) OR
 					(reg_q816 AND symb_decoder(16#36#)) OR
 					(reg_q816 AND symb_decoder(16#f1#)) OR
 					(reg_q816 AND symb_decoder(16#0c#)) OR
 					(reg_q816 AND symb_decoder(16#be#)) OR
 					(reg_q816 AND symb_decoder(16#bf#)) OR
 					(reg_q816 AND symb_decoder(16#94#)) OR
 					(reg_q816 AND symb_decoder(16#ec#)) OR
 					(reg_q816 AND symb_decoder(16#8b#)) OR
 					(reg_q816 AND symb_decoder(16#0d#)) OR
 					(reg_q816 AND symb_decoder(16#63#)) OR
 					(reg_q816 AND symb_decoder(16#e3#)) OR
 					(reg_q816 AND symb_decoder(16#03#)) OR
 					(reg_q816 AND symb_decoder(16#39#)) OR
 					(reg_q816 AND symb_decoder(16#ae#)) OR
 					(reg_q816 AND symb_decoder(16#b7#)) OR
 					(reg_q816 AND symb_decoder(16#18#)) OR
 					(reg_q816 AND symb_decoder(16#c4#)) OR
 					(reg_q816 AND symb_decoder(16#0f#)) OR
 					(reg_q816 AND symb_decoder(16#2a#)) OR
 					(reg_q816 AND symb_decoder(16#50#)) OR
 					(reg_q816 AND symb_decoder(16#c7#)) OR
 					(reg_q816 AND symb_decoder(16#00#)) OR
 					(reg_q816 AND symb_decoder(16#f3#)) OR
 					(reg_q816 AND symb_decoder(16#ad#)) OR
 					(reg_q816 AND symb_decoder(16#42#)) OR
 					(reg_q816 AND symb_decoder(16#6a#)) OR
 					(reg_q816 AND symb_decoder(16#3c#)) OR
 					(reg_q816 AND symb_decoder(16#b3#)) OR
 					(reg_q816 AND symb_decoder(16#59#)) OR
 					(reg_q816 AND symb_decoder(16#05#)) OR
 					(reg_q816 AND symb_decoder(16#01#)) OR
 					(reg_q816 AND symb_decoder(16#cf#)) OR
 					(reg_q816 AND symb_decoder(16#b5#)) OR
 					(reg_q816 AND symb_decoder(16#1b#)) OR
 					(reg_q816 AND symb_decoder(16#82#)) OR
 					(reg_q816 AND symb_decoder(16#fc#)) OR
 					(reg_q816 AND symb_decoder(16#4e#)) OR
 					(reg_q816 AND symb_decoder(16#90#)) OR
 					(reg_q816 AND symb_decoder(16#a8#)) OR
 					(reg_q816 AND symb_decoder(16#38#)) OR
 					(reg_q816 AND symb_decoder(16#22#)) OR
 					(reg_q816 AND symb_decoder(16#67#)) OR
 					(reg_q816 AND symb_decoder(16#f8#)) OR
 					(reg_q816 AND symb_decoder(16#b9#)) OR
 					(reg_q816 AND symb_decoder(16#d1#)) OR
 					(reg_q816 AND symb_decoder(16#85#)) OR
 					(reg_q816 AND symb_decoder(16#34#)) OR
 					(reg_q816 AND symb_decoder(16#af#)) OR
 					(reg_q816 AND symb_decoder(16#46#)) OR
 					(reg_q816 AND symb_decoder(16#c3#)) OR
 					(reg_q816 AND symb_decoder(16#c6#)) OR
 					(reg_q816 AND symb_decoder(16#93#)) OR
 					(reg_q816 AND symb_decoder(16#e4#)) OR
 					(reg_q816 AND symb_decoder(16#30#)) OR
 					(reg_q816 AND symb_decoder(16#13#)) OR
 					(reg_q816 AND symb_decoder(16#fa#)) OR
 					(reg_q816 AND symb_decoder(16#24#)) OR
 					(reg_q816 AND symb_decoder(16#02#)) OR
 					(reg_q816 AND symb_decoder(16#e5#)) OR
 					(reg_q816 AND symb_decoder(16#1f#)) OR
 					(reg_q816 AND symb_decoder(16#a0#)) OR
 					(reg_q816 AND symb_decoder(16#6f#)) OR
 					(reg_q816 AND symb_decoder(16#8d#)) OR
 					(reg_q816 AND symb_decoder(16#72#)) OR
 					(reg_q816 AND symb_decoder(16#55#)) OR
 					(reg_q816 AND symb_decoder(16#6d#)) OR
 					(reg_q816 AND symb_decoder(16#06#)) OR
 					(reg_q816 AND symb_decoder(16#4d#)) OR
 					(reg_q816 AND symb_decoder(16#0e#)) OR
 					(reg_q816 AND symb_decoder(16#25#)) OR
 					(reg_q816 AND symb_decoder(16#31#)) OR
 					(reg_q816 AND symb_decoder(16#de#)) OR
 					(reg_q816 AND symb_decoder(16#09#)) OR
 					(reg_q816 AND symb_decoder(16#e9#)) OR
 					(reg_q816 AND symb_decoder(16#29#)) OR
 					(reg_q816 AND symb_decoder(16#a5#)) OR
 					(reg_q816 AND symb_decoder(16#5d#)) OR
 					(reg_q816 AND symb_decoder(16#a9#)) OR
 					(reg_q816 AND symb_decoder(16#bd#)) OR
 					(reg_q816 AND symb_decoder(16#a1#)) OR
 					(reg_q816 AND symb_decoder(16#71#)) OR
 					(reg_q816 AND symb_decoder(16#4b#)) OR
 					(reg_q816 AND symb_decoder(16#76#)) OR
 					(reg_q816 AND symb_decoder(16#d0#)) OR
 					(reg_q816 AND symb_decoder(16#a6#)) OR
 					(reg_q816 AND symb_decoder(16#2f#)) OR
 					(reg_q816 AND symb_decoder(16#d4#)) OR
 					(reg_q816 AND symb_decoder(16#aa#)) OR
 					(reg_q816 AND symb_decoder(16#a3#)) OR
 					(reg_q816 AND symb_decoder(16#e1#)) OR
 					(reg_q816 AND symb_decoder(16#b4#)) OR
 					(reg_q816 AND symb_decoder(16#37#)) OR
 					(reg_q816 AND symb_decoder(16#c8#)) OR
 					(reg_q816 AND symb_decoder(16#75#)) OR
 					(reg_q816 AND symb_decoder(16#49#)) OR
 					(reg_q816 AND symb_decoder(16#40#)) OR
 					(reg_q816 AND symb_decoder(16#23#)) OR
 					(reg_q816 AND symb_decoder(16#3f#)) OR
 					(reg_q816 AND symb_decoder(16#cb#)) OR
 					(reg_q816 AND symb_decoder(16#da#)) OR
 					(reg_q816 AND symb_decoder(16#f9#)) OR
 					(reg_q816 AND symb_decoder(16#26#)) OR
 					(reg_q816 AND symb_decoder(16#ed#)) OR
 					(reg_q816 AND symb_decoder(16#97#)) OR
 					(reg_q816 AND symb_decoder(16#66#)) OR
 					(reg_q816 AND symb_decoder(16#52#)) OR
 					(reg_q816 AND symb_decoder(16#98#)) OR
 					(reg_q816 AND symb_decoder(16#3a#)) OR
 					(reg_q816 AND symb_decoder(16#16#)) OR
 					(reg_q816 AND symb_decoder(16#d5#)) OR
 					(reg_q816 AND symb_decoder(16#bc#));
reg_q816_init <= '0' ;
	p_reg_q816: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q816 <= reg_q816_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q816 <= reg_q816_init;
        else
          reg_q816 <= reg_q816_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1297_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1297 AND symb_decoder(16#bb#)) OR
 					(reg_q1297 AND symb_decoder(16#3b#)) OR
 					(reg_q1297 AND symb_decoder(16#61#)) OR
 					(reg_q1297 AND symb_decoder(16#6b#)) OR
 					(reg_q1297 AND symb_decoder(16#33#)) OR
 					(reg_q1297 AND symb_decoder(16#fc#)) OR
 					(reg_q1297 AND symb_decoder(16#a5#)) OR
 					(reg_q1297 AND symb_decoder(16#94#)) OR
 					(reg_q1297 AND symb_decoder(16#74#)) OR
 					(reg_q1297 AND symb_decoder(16#84#)) OR
 					(reg_q1297 AND symb_decoder(16#57#)) OR
 					(reg_q1297 AND symb_decoder(16#3d#)) OR
 					(reg_q1297 AND symb_decoder(16#77#)) OR
 					(reg_q1297 AND symb_decoder(16#72#)) OR
 					(reg_q1297 AND symb_decoder(16#4f#)) OR
 					(reg_q1297 AND symb_decoder(16#02#)) OR
 					(reg_q1297 AND symb_decoder(16#e5#)) OR
 					(reg_q1297 AND symb_decoder(16#a0#)) OR
 					(reg_q1297 AND symb_decoder(16#ef#)) OR
 					(reg_q1297 AND symb_decoder(16#18#)) OR
 					(reg_q1297 AND symb_decoder(16#b6#)) OR
 					(reg_q1297 AND symb_decoder(16#cd#)) OR
 					(reg_q1297 AND symb_decoder(16#59#)) OR
 					(reg_q1297 AND symb_decoder(16#cf#)) OR
 					(reg_q1297 AND symb_decoder(16#30#)) OR
 					(reg_q1297 AND symb_decoder(16#e1#)) OR
 					(reg_q1297 AND symb_decoder(16#07#)) OR
 					(reg_q1297 AND symb_decoder(16#c1#)) OR
 					(reg_q1297 AND symb_decoder(16#3f#)) OR
 					(reg_q1297 AND symb_decoder(16#39#)) OR
 					(reg_q1297 AND symb_decoder(16#55#)) OR
 					(reg_q1297 AND symb_decoder(16#6f#)) OR
 					(reg_q1297 AND symb_decoder(16#1e#)) OR
 					(reg_q1297 AND symb_decoder(16#f9#)) OR
 					(reg_q1297 AND symb_decoder(16#7e#)) OR
 					(reg_q1297 AND symb_decoder(16#38#)) OR
 					(reg_q1297 AND symb_decoder(16#09#)) OR
 					(reg_q1297 AND symb_decoder(16#f1#)) OR
 					(reg_q1297 AND symb_decoder(16#a1#)) OR
 					(reg_q1297 AND symb_decoder(16#5a#)) OR
 					(reg_q1297 AND symb_decoder(16#8e#)) OR
 					(reg_q1297 AND symb_decoder(16#52#)) OR
 					(reg_q1297 AND symb_decoder(16#bf#)) OR
 					(reg_q1297 AND symb_decoder(16#64#)) OR
 					(reg_q1297 AND symb_decoder(16#9c#)) OR
 					(reg_q1297 AND symb_decoder(16#86#)) OR
 					(reg_q1297 AND symb_decoder(16#cc#)) OR
 					(reg_q1297 AND symb_decoder(16#0d#)) OR
 					(reg_q1297 AND symb_decoder(16#85#)) OR
 					(reg_q1297 AND symb_decoder(16#67#)) OR
 					(reg_q1297 AND symb_decoder(16#4d#)) OR
 					(reg_q1297 AND symb_decoder(16#aa#)) OR
 					(reg_q1297 AND symb_decoder(16#ba#)) OR
 					(reg_q1297 AND symb_decoder(16#ff#)) OR
 					(reg_q1297 AND symb_decoder(16#34#)) OR
 					(reg_q1297 AND symb_decoder(16#c6#)) OR
 					(reg_q1297 AND symb_decoder(16#4c#)) OR
 					(reg_q1297 AND symb_decoder(16#d9#)) OR
 					(reg_q1297 AND symb_decoder(16#8b#)) OR
 					(reg_q1297 AND symb_decoder(16#a4#)) OR
 					(reg_q1297 AND symb_decoder(16#ce#)) OR
 					(reg_q1297 AND symb_decoder(16#d5#)) OR
 					(reg_q1297 AND symb_decoder(16#6d#)) OR
 					(reg_q1297 AND symb_decoder(16#5f#)) OR
 					(reg_q1297 AND symb_decoder(16#ea#)) OR
 					(reg_q1297 AND symb_decoder(16#56#)) OR
 					(reg_q1297 AND symb_decoder(16#0a#)) OR
 					(reg_q1297 AND symb_decoder(16#81#)) OR
 					(reg_q1297 AND symb_decoder(16#25#)) OR
 					(reg_q1297 AND symb_decoder(16#83#)) OR
 					(reg_q1297 AND symb_decoder(16#58#)) OR
 					(reg_q1297 AND symb_decoder(16#36#)) OR
 					(reg_q1297 AND symb_decoder(16#ad#)) OR
 					(reg_q1297 AND symb_decoder(16#ae#)) OR
 					(reg_q1297 AND symb_decoder(16#05#)) OR
 					(reg_q1297 AND symb_decoder(16#3e#)) OR
 					(reg_q1297 AND symb_decoder(16#b7#)) OR
 					(reg_q1297 AND symb_decoder(16#0e#)) OR
 					(reg_q1297 AND symb_decoder(16#23#)) OR
 					(reg_q1297 AND symb_decoder(16#96#)) OR
 					(reg_q1297 AND symb_decoder(16#51#)) OR
 					(reg_q1297 AND symb_decoder(16#73#)) OR
 					(reg_q1297 AND symb_decoder(16#ca#)) OR
 					(reg_q1297 AND symb_decoder(16#fa#)) OR
 					(reg_q1297 AND symb_decoder(16#d3#)) OR
 					(reg_q1297 AND symb_decoder(16#f5#)) OR
 					(reg_q1297 AND symb_decoder(16#b5#)) OR
 					(reg_q1297 AND symb_decoder(16#2b#)) OR
 					(reg_q1297 AND symb_decoder(16#6e#)) OR
 					(reg_q1297 AND symb_decoder(16#e9#)) OR
 					(reg_q1297 AND symb_decoder(16#15#)) OR
 					(reg_q1297 AND symb_decoder(16#7d#)) OR
 					(reg_q1297 AND symb_decoder(16#42#)) OR
 					(reg_q1297 AND symb_decoder(16#0b#)) OR
 					(reg_q1297 AND symb_decoder(16#2a#)) OR
 					(reg_q1297 AND symb_decoder(16#cb#)) OR
 					(reg_q1297 AND symb_decoder(16#14#)) OR
 					(reg_q1297 AND symb_decoder(16#3a#)) OR
 					(reg_q1297 AND symb_decoder(16#98#)) OR
 					(reg_q1297 AND symb_decoder(16#17#)) OR
 					(reg_q1297 AND symb_decoder(16#dc#)) OR
 					(reg_q1297 AND symb_decoder(16#9e#)) OR
 					(reg_q1297 AND symb_decoder(16#82#)) OR
 					(reg_q1297 AND symb_decoder(16#da#)) OR
 					(reg_q1297 AND symb_decoder(16#8f#)) OR
 					(reg_q1297 AND symb_decoder(16#45#)) OR
 					(reg_q1297 AND symb_decoder(16#9b#)) OR
 					(reg_q1297 AND symb_decoder(16#f0#)) OR
 					(reg_q1297 AND symb_decoder(16#21#)) OR
 					(reg_q1297 AND symb_decoder(16#35#)) OR
 					(reg_q1297 AND symb_decoder(16#a8#)) OR
 					(reg_q1297 AND symb_decoder(16#29#)) OR
 					(reg_q1297 AND symb_decoder(16#48#)) OR
 					(reg_q1297 AND symb_decoder(16#d1#)) OR
 					(reg_q1297 AND symb_decoder(16#d6#)) OR
 					(reg_q1297 AND symb_decoder(16#f2#)) OR
 					(reg_q1297 AND symb_decoder(16#f3#)) OR
 					(reg_q1297 AND symb_decoder(16#8a#)) OR
 					(reg_q1297 AND symb_decoder(16#90#)) OR
 					(reg_q1297 AND symb_decoder(16#3c#)) OR
 					(reg_q1297 AND symb_decoder(16#4b#)) OR
 					(reg_q1297 AND symb_decoder(16#60#)) OR
 					(reg_q1297 AND symb_decoder(16#db#)) OR
 					(reg_q1297 AND symb_decoder(16#b4#)) OR
 					(reg_q1297 AND symb_decoder(16#1d#)) OR
 					(reg_q1297 AND symb_decoder(16#5c#)) OR
 					(reg_q1297 AND symb_decoder(16#7a#)) OR
 					(reg_q1297 AND symb_decoder(16#d0#)) OR
 					(reg_q1297 AND symb_decoder(16#fb#)) OR
 					(reg_q1297 AND symb_decoder(16#0f#)) OR
 					(reg_q1297 AND symb_decoder(16#2d#)) OR
 					(reg_q1297 AND symb_decoder(16#03#)) OR
 					(reg_q1297 AND symb_decoder(16#27#)) OR
 					(reg_q1297 AND symb_decoder(16#49#)) OR
 					(reg_q1297 AND symb_decoder(16#de#)) OR
 					(reg_q1297 AND symb_decoder(16#7f#)) OR
 					(reg_q1297 AND symb_decoder(16#c9#)) OR
 					(reg_q1297 AND symb_decoder(16#04#)) OR
 					(reg_q1297 AND symb_decoder(16#e0#)) OR
 					(reg_q1297 AND symb_decoder(16#c4#)) OR
 					(reg_q1297 AND symb_decoder(16#a9#)) OR
 					(reg_q1297 AND symb_decoder(16#9f#)) OR
 					(reg_q1297 AND symb_decoder(16#65#)) OR
 					(reg_q1297 AND symb_decoder(16#2c#)) OR
 					(reg_q1297 AND symb_decoder(16#df#)) OR
 					(reg_q1297 AND symb_decoder(16#d7#)) OR
 					(reg_q1297 AND symb_decoder(16#46#)) OR
 					(reg_q1297 AND symb_decoder(16#47#)) OR
 					(reg_q1297 AND symb_decoder(16#5d#)) OR
 					(reg_q1297 AND symb_decoder(16#13#)) OR
 					(reg_q1297 AND symb_decoder(16#0c#)) OR
 					(reg_q1297 AND symb_decoder(16#eb#)) OR
 					(reg_q1297 AND symb_decoder(16#41#)) OR
 					(reg_q1297 AND symb_decoder(16#40#)) OR
 					(reg_q1297 AND symb_decoder(16#9d#)) OR
 					(reg_q1297 AND symb_decoder(16#c7#)) OR
 					(reg_q1297 AND symb_decoder(16#b8#)) OR
 					(reg_q1297 AND symb_decoder(16#66#)) OR
 					(reg_q1297 AND symb_decoder(16#f7#)) OR
 					(reg_q1297 AND symb_decoder(16#a7#)) OR
 					(reg_q1297 AND symb_decoder(16#ed#)) OR
 					(reg_q1297 AND symb_decoder(16#53#)) OR
 					(reg_q1297 AND symb_decoder(16#26#)) OR
 					(reg_q1297 AND symb_decoder(16#16#)) OR
 					(reg_q1297 AND symb_decoder(16#c8#)) OR
 					(reg_q1297 AND symb_decoder(16#62#)) OR
 					(reg_q1297 AND symb_decoder(16#1b#)) OR
 					(reg_q1297 AND symb_decoder(16#d2#)) OR
 					(reg_q1297 AND symb_decoder(16#69#)) OR
 					(reg_q1297 AND symb_decoder(16#e6#)) OR
 					(reg_q1297 AND symb_decoder(16#af#)) OR
 					(reg_q1297 AND symb_decoder(16#f8#)) OR
 					(reg_q1297 AND symb_decoder(16#bc#)) OR
 					(reg_q1297 AND symb_decoder(16#54#)) OR
 					(reg_q1297 AND symb_decoder(16#00#)) OR
 					(reg_q1297 AND symb_decoder(16#22#)) OR
 					(reg_q1297 AND symb_decoder(16#99#)) OR
 					(reg_q1297 AND symb_decoder(16#93#)) OR
 					(reg_q1297 AND symb_decoder(16#8c#)) OR
 					(reg_q1297 AND symb_decoder(16#68#)) OR
 					(reg_q1297 AND symb_decoder(16#2e#)) OR
 					(reg_q1297 AND symb_decoder(16#5e#)) OR
 					(reg_q1297 AND symb_decoder(16#4e#)) OR
 					(reg_q1297 AND symb_decoder(16#2f#)) OR
 					(reg_q1297 AND symb_decoder(16#70#)) OR
 					(reg_q1297 AND symb_decoder(16#9a#)) OR
 					(reg_q1297 AND symb_decoder(16#91#)) OR
 					(reg_q1297 AND symb_decoder(16#ac#)) OR
 					(reg_q1297 AND symb_decoder(16#1c#)) OR
 					(reg_q1297 AND symb_decoder(16#d8#)) OR
 					(reg_q1297 AND symb_decoder(16#75#)) OR
 					(reg_q1297 AND symb_decoder(16#a3#)) OR
 					(reg_q1297 AND symb_decoder(16#f6#)) OR
 					(reg_q1297 AND symb_decoder(16#a6#)) OR
 					(reg_q1297 AND symb_decoder(16#76#)) OR
 					(reg_q1297 AND symb_decoder(16#fd#)) OR
 					(reg_q1297 AND symb_decoder(16#4a#)) OR
 					(reg_q1297 AND symb_decoder(16#95#)) OR
 					(reg_q1297 AND symb_decoder(16#e2#)) OR
 					(reg_q1297 AND symb_decoder(16#97#)) OR
 					(reg_q1297 AND symb_decoder(16#b2#)) OR
 					(reg_q1297 AND symb_decoder(16#63#)) OR
 					(reg_q1297 AND symb_decoder(16#f4#)) OR
 					(reg_q1297 AND symb_decoder(16#19#)) OR
 					(reg_q1297 AND symb_decoder(16#6c#)) OR
 					(reg_q1297 AND symb_decoder(16#88#)) OR
 					(reg_q1297 AND symb_decoder(16#50#)) OR
 					(reg_q1297 AND symb_decoder(16#5b#)) OR
 					(reg_q1297 AND symb_decoder(16#06#)) OR
 					(reg_q1297 AND symb_decoder(16#43#)) OR
 					(reg_q1297 AND symb_decoder(16#b1#)) OR
 					(reg_q1297 AND symb_decoder(16#e8#)) OR
 					(reg_q1297 AND symb_decoder(16#28#)) OR
 					(reg_q1297 AND symb_decoder(16#ee#)) OR
 					(reg_q1297 AND symb_decoder(16#8d#)) OR
 					(reg_q1297 AND symb_decoder(16#1a#)) OR
 					(reg_q1297 AND symb_decoder(16#80#)) OR
 					(reg_q1297 AND symb_decoder(16#b9#)) OR
 					(reg_q1297 AND symb_decoder(16#e4#)) OR
 					(reg_q1297 AND symb_decoder(16#e7#)) OR
 					(reg_q1297 AND symb_decoder(16#fe#)) OR
 					(reg_q1297 AND symb_decoder(16#31#)) OR
 					(reg_q1297 AND symb_decoder(16#12#)) OR
 					(reg_q1297 AND symb_decoder(16#c5#)) OR
 					(reg_q1297 AND symb_decoder(16#11#)) OR
 					(reg_q1297 AND symb_decoder(16#6a#)) OR
 					(reg_q1297 AND symb_decoder(16#bd#)) OR
 					(reg_q1297 AND symb_decoder(16#1f#)) OR
 					(reg_q1297 AND symb_decoder(16#10#)) OR
 					(reg_q1297 AND symb_decoder(16#dd#)) OR
 					(reg_q1297 AND symb_decoder(16#c2#)) OR
 					(reg_q1297 AND symb_decoder(16#a2#)) OR
 					(reg_q1297 AND symb_decoder(16#71#)) OR
 					(reg_q1297 AND symb_decoder(16#c3#)) OR
 					(reg_q1297 AND symb_decoder(16#e3#)) OR
 					(reg_q1297 AND symb_decoder(16#7b#)) OR
 					(reg_q1297 AND symb_decoder(16#37#)) OR
 					(reg_q1297 AND symb_decoder(16#ec#)) OR
 					(reg_q1297 AND symb_decoder(16#d4#)) OR
 					(reg_q1297 AND symb_decoder(16#be#)) OR
 					(reg_q1297 AND symb_decoder(16#ab#)) OR
 					(reg_q1297 AND symb_decoder(16#01#)) OR
 					(reg_q1297 AND symb_decoder(16#20#)) OR
 					(reg_q1297 AND symb_decoder(16#89#)) OR
 					(reg_q1297 AND symb_decoder(16#87#)) OR
 					(reg_q1297 AND symb_decoder(16#c0#)) OR
 					(reg_q1297 AND symb_decoder(16#24#)) OR
 					(reg_q1297 AND symb_decoder(16#32#)) OR
 					(reg_q1297 AND symb_decoder(16#78#)) OR
 					(reg_q1297 AND symb_decoder(16#08#)) OR
 					(reg_q1297 AND symb_decoder(16#92#)) OR
 					(reg_q1297 AND symb_decoder(16#79#)) OR
 					(reg_q1297 AND symb_decoder(16#44#)) OR
 					(reg_q1297 AND symb_decoder(16#b3#)) OR
 					(reg_q1297 AND symb_decoder(16#b0#)) OR
 					(reg_q1297 AND symb_decoder(16#7c#));
reg_q1297_init <= '0' ;
	p_reg_q1297: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1297 <= reg_q1297_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1297 <= reg_q1297_init;
        else
          reg_q1297 <= reg_q1297_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2618_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2618 AND symb_decoder(16#0f#)) OR
 					(reg_q2618 AND symb_decoder(16#eb#)) OR
 					(reg_q2618 AND symb_decoder(16#48#)) OR
 					(reg_q2618 AND symb_decoder(16#d0#)) OR
 					(reg_q2618 AND symb_decoder(16#e0#)) OR
 					(reg_q2618 AND symb_decoder(16#9c#)) OR
 					(reg_q2618 AND symb_decoder(16#59#)) OR
 					(reg_q2618 AND symb_decoder(16#98#)) OR
 					(reg_q2618 AND symb_decoder(16#7d#)) OR
 					(reg_q2618 AND symb_decoder(16#67#)) OR
 					(reg_q2618 AND symb_decoder(16#1f#)) OR
 					(reg_q2618 AND symb_decoder(16#65#)) OR
 					(reg_q2618 AND symb_decoder(16#74#)) OR
 					(reg_q2618 AND symb_decoder(16#0a#)) OR
 					(reg_q2618 AND symb_decoder(16#83#)) OR
 					(reg_q2618 AND symb_decoder(16#f1#)) OR
 					(reg_q2618 AND symb_decoder(16#4e#)) OR
 					(reg_q2618 AND symb_decoder(16#99#)) OR
 					(reg_q2618 AND symb_decoder(16#55#)) OR
 					(reg_q2618 AND symb_decoder(16#8a#)) OR
 					(reg_q2618 AND symb_decoder(16#4c#)) OR
 					(reg_q2618 AND symb_decoder(16#49#)) OR
 					(reg_q2618 AND symb_decoder(16#5b#)) OR
 					(reg_q2618 AND symb_decoder(16#06#)) OR
 					(reg_q2618 AND symb_decoder(16#ca#)) OR
 					(reg_q2618 AND symb_decoder(16#8c#)) OR
 					(reg_q2618 AND symb_decoder(16#93#)) OR
 					(reg_q2618 AND symb_decoder(16#6d#)) OR
 					(reg_q2618 AND symb_decoder(16#14#)) OR
 					(reg_q2618 AND symb_decoder(16#62#)) OR
 					(reg_q2618 AND symb_decoder(16#1b#)) OR
 					(reg_q2618 AND symb_decoder(16#2d#)) OR
 					(reg_q2618 AND symb_decoder(16#78#)) OR
 					(reg_q2618 AND symb_decoder(16#6a#)) OR
 					(reg_q2618 AND symb_decoder(16#ee#)) OR
 					(reg_q2618 AND symb_decoder(16#d4#)) OR
 					(reg_q2618 AND symb_decoder(16#53#)) OR
 					(reg_q2618 AND symb_decoder(16#a1#)) OR
 					(reg_q2618 AND symb_decoder(16#07#)) OR
 					(reg_q2618 AND symb_decoder(16#3c#)) OR
 					(reg_q2618 AND symb_decoder(16#e4#)) OR
 					(reg_q2618 AND symb_decoder(16#f5#)) OR
 					(reg_q2618 AND symb_decoder(16#c4#)) OR
 					(reg_q2618 AND symb_decoder(16#5e#)) OR
 					(reg_q2618 AND symb_decoder(16#ae#)) OR
 					(reg_q2618 AND symb_decoder(16#08#)) OR
 					(reg_q2618 AND symb_decoder(16#40#)) OR
 					(reg_q2618 AND symb_decoder(16#c6#)) OR
 					(reg_q2618 AND symb_decoder(16#39#)) OR
 					(reg_q2618 AND symb_decoder(16#2e#)) OR
 					(reg_q2618 AND symb_decoder(16#ff#)) OR
 					(reg_q2618 AND symb_decoder(16#8d#)) OR
 					(reg_q2618 AND symb_decoder(16#51#)) OR
 					(reg_q2618 AND symb_decoder(16#c1#)) OR
 					(reg_q2618 AND symb_decoder(16#a2#)) OR
 					(reg_q2618 AND symb_decoder(16#ab#)) OR
 					(reg_q2618 AND symb_decoder(16#7a#)) OR
 					(reg_q2618 AND symb_decoder(16#ad#)) OR
 					(reg_q2618 AND symb_decoder(16#97#)) OR
 					(reg_q2618 AND symb_decoder(16#d3#)) OR
 					(reg_q2618 AND symb_decoder(16#03#)) OR
 					(reg_q2618 AND symb_decoder(16#7b#)) OR
 					(reg_q2618 AND symb_decoder(16#2f#)) OR
 					(reg_q2618 AND symb_decoder(16#2b#)) OR
 					(reg_q2618 AND symb_decoder(16#00#)) OR
 					(reg_q2618 AND symb_decoder(16#17#)) OR
 					(reg_q2618 AND symb_decoder(16#73#)) OR
 					(reg_q2618 AND symb_decoder(16#13#)) OR
 					(reg_q2618 AND symb_decoder(16#80#)) OR
 					(reg_q2618 AND symb_decoder(16#12#)) OR
 					(reg_q2618 AND symb_decoder(16#71#)) OR
 					(reg_q2618 AND symb_decoder(16#e8#)) OR
 					(reg_q2618 AND symb_decoder(16#b5#)) OR
 					(reg_q2618 AND symb_decoder(16#d6#)) OR
 					(reg_q2618 AND symb_decoder(16#d9#)) OR
 					(reg_q2618 AND symb_decoder(16#57#)) OR
 					(reg_q2618 AND symb_decoder(16#5a#)) OR
 					(reg_q2618 AND symb_decoder(16#c9#)) OR
 					(reg_q2618 AND symb_decoder(16#bd#)) OR
 					(reg_q2618 AND symb_decoder(16#dd#)) OR
 					(reg_q2618 AND symb_decoder(16#11#)) OR
 					(reg_q2618 AND symb_decoder(16#87#)) OR
 					(reg_q2618 AND symb_decoder(16#33#)) OR
 					(reg_q2618 AND symb_decoder(16#d2#)) OR
 					(reg_q2618 AND symb_decoder(16#54#)) OR
 					(reg_q2618 AND symb_decoder(16#4a#)) OR
 					(reg_q2618 AND symb_decoder(16#bb#)) OR
 					(reg_q2618 AND symb_decoder(16#af#)) OR
 					(reg_q2618 AND symb_decoder(16#b9#)) OR
 					(reg_q2618 AND symb_decoder(16#e9#)) OR
 					(reg_q2618 AND symb_decoder(16#1a#)) OR
 					(reg_q2618 AND symb_decoder(16#a4#)) OR
 					(reg_q2618 AND symb_decoder(16#92#)) OR
 					(reg_q2618 AND symb_decoder(16#7e#)) OR
 					(reg_q2618 AND symb_decoder(16#77#)) OR
 					(reg_q2618 AND symb_decoder(16#f8#)) OR
 					(reg_q2618 AND symb_decoder(16#cb#)) OR
 					(reg_q2618 AND symb_decoder(16#84#)) OR
 					(reg_q2618 AND symb_decoder(16#e2#)) OR
 					(reg_q2618 AND symb_decoder(16#b0#)) OR
 					(reg_q2618 AND symb_decoder(16#43#)) OR
 					(reg_q2618 AND symb_decoder(16#ea#)) OR
 					(reg_q2618 AND symb_decoder(16#be#)) OR
 					(reg_q2618 AND symb_decoder(16#c0#)) OR
 					(reg_q2618 AND symb_decoder(16#89#)) OR
 					(reg_q2618 AND symb_decoder(16#dc#)) OR
 					(reg_q2618 AND symb_decoder(16#b4#)) OR
 					(reg_q2618 AND symb_decoder(16#82#)) OR
 					(reg_q2618 AND symb_decoder(16#86#)) OR
 					(reg_q2618 AND symb_decoder(16#41#)) OR
 					(reg_q2618 AND symb_decoder(16#e3#)) OR
 					(reg_q2618 AND symb_decoder(16#8e#)) OR
 					(reg_q2618 AND symb_decoder(16#35#)) OR
 					(reg_q2618 AND symb_decoder(16#a8#)) OR
 					(reg_q2618 AND symb_decoder(16#3b#)) OR
 					(reg_q2618 AND symb_decoder(16#20#)) OR
 					(reg_q2618 AND symb_decoder(16#90#)) OR
 					(reg_q2618 AND symb_decoder(16#f0#)) OR
 					(reg_q2618 AND symb_decoder(16#26#)) OR
 					(reg_q2618 AND symb_decoder(16#d7#)) OR
 					(reg_q2618 AND symb_decoder(16#31#)) OR
 					(reg_q2618 AND symb_decoder(16#c5#)) OR
 					(reg_q2618 AND symb_decoder(16#36#)) OR
 					(reg_q2618 AND symb_decoder(16#47#)) OR
 					(reg_q2618 AND symb_decoder(16#01#)) OR
 					(reg_q2618 AND symb_decoder(16#79#)) OR
 					(reg_q2618 AND symb_decoder(16#c7#)) OR
 					(reg_q2618 AND symb_decoder(16#32#)) OR
 					(reg_q2618 AND symb_decoder(16#ed#)) OR
 					(reg_q2618 AND symb_decoder(16#16#)) OR
 					(reg_q2618 AND symb_decoder(16#75#)) OR
 					(reg_q2618 AND symb_decoder(16#0e#)) OR
 					(reg_q2618 AND symb_decoder(16#42#)) OR
 					(reg_q2618 AND symb_decoder(16#19#)) OR
 					(reg_q2618 AND symb_decoder(16#2a#)) OR
 					(reg_q2618 AND symb_decoder(16#c3#)) OR
 					(reg_q2618 AND symb_decoder(16#3f#)) OR
 					(reg_q2618 AND symb_decoder(16#69#)) OR
 					(reg_q2618 AND symb_decoder(16#0b#)) OR
 					(reg_q2618 AND symb_decoder(16#15#)) OR
 					(reg_q2618 AND symb_decoder(16#09#)) OR
 					(reg_q2618 AND symb_decoder(16#e7#)) OR
 					(reg_q2618 AND symb_decoder(16#04#)) OR
 					(reg_q2618 AND symb_decoder(16#05#)) OR
 					(reg_q2618 AND symb_decoder(16#7f#)) OR
 					(reg_q2618 AND symb_decoder(16#cd#)) OR
 					(reg_q2618 AND symb_decoder(16#18#)) OR
 					(reg_q2618 AND symb_decoder(16#f9#)) OR
 					(reg_q2618 AND symb_decoder(16#0d#)) OR
 					(reg_q2618 AND symb_decoder(16#da#)) OR
 					(reg_q2618 AND symb_decoder(16#64#)) OR
 					(reg_q2618 AND symb_decoder(16#9d#)) OR
 					(reg_q2618 AND symb_decoder(16#cf#)) OR
 					(reg_q2618 AND symb_decoder(16#a9#)) OR
 					(reg_q2618 AND symb_decoder(16#60#)) OR
 					(reg_q2618 AND symb_decoder(16#30#)) OR
 					(reg_q2618 AND symb_decoder(16#96#)) OR
 					(reg_q2618 AND symb_decoder(16#28#)) OR
 					(reg_q2618 AND symb_decoder(16#aa#)) OR
 					(reg_q2618 AND symb_decoder(16#f4#)) OR
 					(reg_q2618 AND symb_decoder(16#6f#)) OR
 					(reg_q2618 AND symb_decoder(16#10#)) OR
 					(reg_q2618 AND symb_decoder(16#3e#)) OR
 					(reg_q2618 AND symb_decoder(16#e5#)) OR
 					(reg_q2618 AND symb_decoder(16#a5#)) OR
 					(reg_q2618 AND symb_decoder(16#c8#)) OR
 					(reg_q2618 AND symb_decoder(16#df#)) OR
 					(reg_q2618 AND symb_decoder(16#6b#)) OR
 					(reg_q2618 AND symb_decoder(16#58#)) OR
 					(reg_q2618 AND symb_decoder(16#4f#)) OR
 					(reg_q2618 AND symb_decoder(16#34#)) OR
 					(reg_q2618 AND symb_decoder(16#f7#)) OR
 					(reg_q2618 AND symb_decoder(16#3d#)) OR
 					(reg_q2618 AND symb_decoder(16#24#)) OR
 					(reg_q2618 AND symb_decoder(16#46#)) OR
 					(reg_q2618 AND symb_decoder(16#de#)) OR
 					(reg_q2618 AND symb_decoder(16#9b#)) OR
 					(reg_q2618 AND symb_decoder(16#ef#)) OR
 					(reg_q2618 AND symb_decoder(16#37#)) OR
 					(reg_q2618 AND symb_decoder(16#c2#)) OR
 					(reg_q2618 AND symb_decoder(16#d5#)) OR
 					(reg_q2618 AND symb_decoder(16#5c#)) OR
 					(reg_q2618 AND symb_decoder(16#1c#)) OR
 					(reg_q2618 AND symb_decoder(16#e1#)) OR
 					(reg_q2618 AND symb_decoder(16#b7#)) OR
 					(reg_q2618 AND symb_decoder(16#70#)) OR
 					(reg_q2618 AND symb_decoder(16#76#)) OR
 					(reg_q2618 AND symb_decoder(16#23#)) OR
 					(reg_q2618 AND symb_decoder(16#bf#)) OR
 					(reg_q2618 AND symb_decoder(16#5f#)) OR
 					(reg_q2618 AND symb_decoder(16#d8#)) OR
 					(reg_q2618 AND symb_decoder(16#bc#)) OR
 					(reg_q2618 AND symb_decoder(16#21#)) OR
 					(reg_q2618 AND symb_decoder(16#6e#)) OR
 					(reg_q2618 AND symb_decoder(16#a7#)) OR
 					(reg_q2618 AND symb_decoder(16#50#)) OR
 					(reg_q2618 AND symb_decoder(16#a6#)) OR
 					(reg_q2618 AND symb_decoder(16#94#)) OR
 					(reg_q2618 AND symb_decoder(16#d1#)) OR
 					(reg_q2618 AND symb_decoder(16#45#)) OR
 					(reg_q2618 AND symb_decoder(16#b2#)) OR
 					(reg_q2618 AND symb_decoder(16#7c#)) OR
 					(reg_q2618 AND symb_decoder(16#ec#)) OR
 					(reg_q2618 AND symb_decoder(16#68#)) OR
 					(reg_q2618 AND symb_decoder(16#fb#)) OR
 					(reg_q2618 AND symb_decoder(16#f6#)) OR
 					(reg_q2618 AND symb_decoder(16#e6#)) OR
 					(reg_q2618 AND symb_decoder(16#29#)) OR
 					(reg_q2618 AND symb_decoder(16#91#)) OR
 					(reg_q2618 AND symb_decoder(16#ac#)) OR
 					(reg_q2618 AND symb_decoder(16#b1#)) OR
 					(reg_q2618 AND symb_decoder(16#85#)) OR
 					(reg_q2618 AND symb_decoder(16#f3#)) OR
 					(reg_q2618 AND symb_decoder(16#88#)) OR
 					(reg_q2618 AND symb_decoder(16#4d#)) OR
 					(reg_q2618 AND symb_decoder(16#63#)) OR
 					(reg_q2618 AND symb_decoder(16#9a#)) OR
 					(reg_q2618 AND symb_decoder(16#b6#)) OR
 					(reg_q2618 AND symb_decoder(16#fe#)) OR
 					(reg_q2618 AND symb_decoder(16#27#)) OR
 					(reg_q2618 AND symb_decoder(16#fa#)) OR
 					(reg_q2618 AND symb_decoder(16#02#)) OR
 					(reg_q2618 AND symb_decoder(16#6c#)) OR
 					(reg_q2618 AND symb_decoder(16#f2#)) OR
 					(reg_q2618 AND symb_decoder(16#db#)) OR
 					(reg_q2618 AND symb_decoder(16#52#)) OR
 					(reg_q2618 AND symb_decoder(16#ce#)) OR
 					(reg_q2618 AND symb_decoder(16#2c#)) OR
 					(reg_q2618 AND symb_decoder(16#a3#)) OR
 					(reg_q2618 AND symb_decoder(16#b3#)) OR
 					(reg_q2618 AND symb_decoder(16#9e#)) OR
 					(reg_q2618 AND symb_decoder(16#8b#)) OR
 					(reg_q2618 AND symb_decoder(16#81#)) OR
 					(reg_q2618 AND symb_decoder(16#cc#)) OR
 					(reg_q2618 AND symb_decoder(16#44#)) OR
 					(reg_q2618 AND symb_decoder(16#3a#)) OR
 					(reg_q2618 AND symb_decoder(16#95#)) OR
 					(reg_q2618 AND symb_decoder(16#61#)) OR
 					(reg_q2618 AND symb_decoder(16#25#)) OR
 					(reg_q2618 AND symb_decoder(16#1d#)) OR
 					(reg_q2618 AND symb_decoder(16#56#)) OR
 					(reg_q2618 AND symb_decoder(16#22#)) OR
 					(reg_q2618 AND symb_decoder(16#a0#)) OR
 					(reg_q2618 AND symb_decoder(16#b8#)) OR
 					(reg_q2618 AND symb_decoder(16#fd#)) OR
 					(reg_q2618 AND symb_decoder(16#72#)) OR
 					(reg_q2618 AND symb_decoder(16#5d#)) OR
 					(reg_q2618 AND symb_decoder(16#1e#)) OR
 					(reg_q2618 AND symb_decoder(16#fc#)) OR
 					(reg_q2618 AND symb_decoder(16#0c#)) OR
 					(reg_q2618 AND symb_decoder(16#9f#)) OR
 					(reg_q2618 AND symb_decoder(16#ba#)) OR
 					(reg_q2618 AND symb_decoder(16#38#)) OR
 					(reg_q2618 AND symb_decoder(16#66#)) OR
 					(reg_q2618 AND symb_decoder(16#4b#)) OR
 					(reg_q2618 AND symb_decoder(16#8f#));
reg_q2618_init <= '0' ;
	p_reg_q2618: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2618 <= reg_q2618_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2618 <= reg_q2618_init;
        else
          reg_q2618 <= reg_q2618_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q850_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q850 AND symb_decoder(16#20#)) OR
 					(reg_q850 AND symb_decoder(16#5e#)) OR
 					(reg_q850 AND symb_decoder(16#46#)) OR
 					(reg_q850 AND symb_decoder(16#d4#)) OR
 					(reg_q850 AND symb_decoder(16#e0#)) OR
 					(reg_q850 AND symb_decoder(16#2f#)) OR
 					(reg_q850 AND symb_decoder(16#0c#)) OR
 					(reg_q850 AND symb_decoder(16#6f#)) OR
 					(reg_q850 AND symb_decoder(16#7f#)) OR
 					(reg_q850 AND symb_decoder(16#10#)) OR
 					(reg_q850 AND symb_decoder(16#5f#)) OR
 					(reg_q850 AND symb_decoder(16#a6#)) OR
 					(reg_q850 AND symb_decoder(16#0a#)) OR
 					(reg_q850 AND symb_decoder(16#29#)) OR
 					(reg_q850 AND symb_decoder(16#c4#)) OR
 					(reg_q850 AND symb_decoder(16#fc#)) OR
 					(reg_q850 AND symb_decoder(16#76#)) OR
 					(reg_q850 AND symb_decoder(16#2c#)) OR
 					(reg_q850 AND symb_decoder(16#8c#)) OR
 					(reg_q850 AND symb_decoder(16#24#)) OR
 					(reg_q850 AND symb_decoder(16#c6#)) OR
 					(reg_q850 AND symb_decoder(16#0b#)) OR
 					(reg_q850 AND symb_decoder(16#12#)) OR
 					(reg_q850 AND symb_decoder(16#6c#)) OR
 					(reg_q850 AND symb_decoder(16#f5#)) OR
 					(reg_q850 AND symb_decoder(16#1c#)) OR
 					(reg_q850 AND symb_decoder(16#04#)) OR
 					(reg_q850 AND symb_decoder(16#48#)) OR
 					(reg_q850 AND symb_decoder(16#86#)) OR
 					(reg_q850 AND symb_decoder(16#81#)) OR
 					(reg_q850 AND symb_decoder(16#bb#)) OR
 					(reg_q850 AND symb_decoder(16#e3#)) OR
 					(reg_q850 AND symb_decoder(16#73#)) OR
 					(reg_q850 AND symb_decoder(16#5b#)) OR
 					(reg_q850 AND symb_decoder(16#83#)) OR
 					(reg_q850 AND symb_decoder(16#dd#)) OR
 					(reg_q850 AND symb_decoder(16#90#)) OR
 					(reg_q850 AND symb_decoder(16#19#)) OR
 					(reg_q850 AND symb_decoder(16#99#)) OR
 					(reg_q850 AND symb_decoder(16#bc#)) OR
 					(reg_q850 AND symb_decoder(16#b4#)) OR
 					(reg_q850 AND symb_decoder(16#9c#)) OR
 					(reg_q850 AND symb_decoder(16#41#)) OR
 					(reg_q850 AND symb_decoder(16#cb#)) OR
 					(reg_q850 AND symb_decoder(16#d0#)) OR
 					(reg_q850 AND symb_decoder(16#5c#)) OR
 					(reg_q850 AND symb_decoder(16#33#)) OR
 					(reg_q850 AND symb_decoder(16#e7#)) OR
 					(reg_q850 AND symb_decoder(16#74#)) OR
 					(reg_q850 AND symb_decoder(16#05#)) OR
 					(reg_q850 AND symb_decoder(16#0d#)) OR
 					(reg_q850 AND symb_decoder(16#17#)) OR
 					(reg_q850 AND symb_decoder(16#30#)) OR
 					(reg_q850 AND symb_decoder(16#4b#)) OR
 					(reg_q850 AND symb_decoder(16#36#)) OR
 					(reg_q850 AND symb_decoder(16#e4#)) OR
 					(reg_q850 AND symb_decoder(16#b8#)) OR
 					(reg_q850 AND symb_decoder(16#7d#)) OR
 					(reg_q850 AND symb_decoder(16#f8#)) OR
 					(reg_q850 AND symb_decoder(16#4f#)) OR
 					(reg_q850 AND symb_decoder(16#aa#)) OR
 					(reg_q850 AND symb_decoder(16#e2#)) OR
 					(reg_q850 AND symb_decoder(16#55#)) OR
 					(reg_q850 AND symb_decoder(16#58#)) OR
 					(reg_q850 AND symb_decoder(16#ec#)) OR
 					(reg_q850 AND symb_decoder(16#d7#)) OR
 					(reg_q850 AND symb_decoder(16#69#)) OR
 					(reg_q850 AND symb_decoder(16#d1#)) OR
 					(reg_q850 AND symb_decoder(16#ee#)) OR
 					(reg_q850 AND symb_decoder(16#34#)) OR
 					(reg_q850 AND symb_decoder(16#2e#)) OR
 					(reg_q850 AND symb_decoder(16#4a#)) OR
 					(reg_q850 AND symb_decoder(16#09#)) OR
 					(reg_q850 AND symb_decoder(16#32#)) OR
 					(reg_q850 AND symb_decoder(16#01#)) OR
 					(reg_q850 AND symb_decoder(16#28#)) OR
 					(reg_q850 AND symb_decoder(16#07#)) OR
 					(reg_q850 AND symb_decoder(16#22#)) OR
 					(reg_q850 AND symb_decoder(16#e9#)) OR
 					(reg_q850 AND symb_decoder(16#0f#)) OR
 					(reg_q850 AND symb_decoder(16#eb#)) OR
 					(reg_q850 AND symb_decoder(16#1b#)) OR
 					(reg_q850 AND symb_decoder(16#16#)) OR
 					(reg_q850 AND symb_decoder(16#72#)) OR
 					(reg_q850 AND symb_decoder(16#c7#)) OR
 					(reg_q850 AND symb_decoder(16#c0#)) OR
 					(reg_q850 AND symb_decoder(16#02#)) OR
 					(reg_q850 AND symb_decoder(16#d3#)) OR
 					(reg_q850 AND symb_decoder(16#3c#)) OR
 					(reg_q850 AND symb_decoder(16#47#)) OR
 					(reg_q850 AND symb_decoder(16#56#)) OR
 					(reg_q850 AND symb_decoder(16#a5#)) OR
 					(reg_q850 AND symb_decoder(16#31#)) OR
 					(reg_q850 AND symb_decoder(16#7a#)) OR
 					(reg_q850 AND symb_decoder(16#00#)) OR
 					(reg_q850 AND symb_decoder(16#b5#)) OR
 					(reg_q850 AND symb_decoder(16#8f#)) OR
 					(reg_q850 AND symb_decoder(16#bd#)) OR
 					(reg_q850 AND symb_decoder(16#4e#)) OR
 					(reg_q850 AND symb_decoder(16#23#)) OR
 					(reg_q850 AND symb_decoder(16#85#)) OR
 					(reg_q850 AND symb_decoder(16#5a#)) OR
 					(reg_q850 AND symb_decoder(16#03#)) OR
 					(reg_q850 AND symb_decoder(16#7e#)) OR
 					(reg_q850 AND symb_decoder(16#21#)) OR
 					(reg_q850 AND symb_decoder(16#18#)) OR
 					(reg_q850 AND symb_decoder(16#26#)) OR
 					(reg_q850 AND symb_decoder(16#b6#)) OR
 					(reg_q850 AND symb_decoder(16#b2#)) OR
 					(reg_q850 AND symb_decoder(16#37#)) OR
 					(reg_q850 AND symb_decoder(16#13#)) OR
 					(reg_q850 AND symb_decoder(16#b0#)) OR
 					(reg_q850 AND symb_decoder(16#9f#)) OR
 					(reg_q850 AND symb_decoder(16#8a#)) OR
 					(reg_q850 AND symb_decoder(16#cf#)) OR
 					(reg_q850 AND symb_decoder(16#f4#)) OR
 					(reg_q850 AND symb_decoder(16#a4#)) OR
 					(reg_q850 AND symb_decoder(16#80#)) OR
 					(reg_q850 AND symb_decoder(16#7b#)) OR
 					(reg_q850 AND symb_decoder(16#3f#)) OR
 					(reg_q850 AND symb_decoder(16#fb#)) OR
 					(reg_q850 AND symb_decoder(16#c2#)) OR
 					(reg_q850 AND symb_decoder(16#cd#)) OR
 					(reg_q850 AND symb_decoder(16#a1#)) OR
 					(reg_q850 AND symb_decoder(16#f9#)) OR
 					(reg_q850 AND symb_decoder(16#38#)) OR
 					(reg_q850 AND symb_decoder(16#54#)) OR
 					(reg_q850 AND symb_decoder(16#1a#)) OR
 					(reg_q850 AND symb_decoder(16#68#)) OR
 					(reg_q850 AND symb_decoder(16#51#)) OR
 					(reg_q850 AND symb_decoder(16#d2#)) OR
 					(reg_q850 AND symb_decoder(16#42#)) OR
 					(reg_q850 AND symb_decoder(16#77#)) OR
 					(reg_q850 AND symb_decoder(16#06#)) OR
 					(reg_q850 AND symb_decoder(16#89#)) OR
 					(reg_q850 AND symb_decoder(16#78#)) OR
 					(reg_q850 AND symb_decoder(16#3e#)) OR
 					(reg_q850 AND symb_decoder(16#67#)) OR
 					(reg_q850 AND symb_decoder(16#75#)) OR
 					(reg_q850 AND symb_decoder(16#d9#)) OR
 					(reg_q850 AND symb_decoder(16#ca#)) OR
 					(reg_q850 AND symb_decoder(16#c8#)) OR
 					(reg_q850 AND symb_decoder(16#79#)) OR
 					(reg_q850 AND symb_decoder(16#a3#)) OR
 					(reg_q850 AND symb_decoder(16#a2#)) OR
 					(reg_q850 AND symb_decoder(16#65#)) OR
 					(reg_q850 AND symb_decoder(16#0e#)) OR
 					(reg_q850 AND symb_decoder(16#94#)) OR
 					(reg_q850 AND symb_decoder(16#fa#)) OR
 					(reg_q850 AND symb_decoder(16#40#)) OR
 					(reg_q850 AND symb_decoder(16#6d#)) OR
 					(reg_q850 AND symb_decoder(16#84#)) OR
 					(reg_q850 AND symb_decoder(16#93#)) OR
 					(reg_q850 AND symb_decoder(16#64#)) OR
 					(reg_q850 AND symb_decoder(16#c5#)) OR
 					(reg_q850 AND symb_decoder(16#ac#)) OR
 					(reg_q850 AND symb_decoder(16#88#)) OR
 					(reg_q850 AND symb_decoder(16#cc#)) OR
 					(reg_q850 AND symb_decoder(16#60#)) OR
 					(reg_q850 AND symb_decoder(16#e1#)) OR
 					(reg_q850 AND symb_decoder(16#d8#)) OR
 					(reg_q850 AND symb_decoder(16#50#)) OR
 					(reg_q850 AND symb_decoder(16#a0#)) OR
 					(reg_q850 AND symb_decoder(16#3b#)) OR
 					(reg_q850 AND symb_decoder(16#91#)) OR
 					(reg_q850 AND symb_decoder(16#3a#)) OR
 					(reg_q850 AND symb_decoder(16#2d#)) OR
 					(reg_q850 AND symb_decoder(16#1d#)) OR
 					(reg_q850 AND symb_decoder(16#8d#)) OR
 					(reg_q850 AND symb_decoder(16#3d#)) OR
 					(reg_q850 AND symb_decoder(16#ae#)) OR
 					(reg_q850 AND symb_decoder(16#c1#)) OR
 					(reg_q850 AND symb_decoder(16#6b#)) OR
 					(reg_q850 AND symb_decoder(16#49#)) OR
 					(reg_q850 AND symb_decoder(16#08#)) OR
 					(reg_q850 AND symb_decoder(16#52#)) OR
 					(reg_q850 AND symb_decoder(16#be#)) OR
 					(reg_q850 AND symb_decoder(16#6e#)) OR
 					(reg_q850 AND symb_decoder(16#1f#)) OR
 					(reg_q850 AND symb_decoder(16#53#)) OR
 					(reg_q850 AND symb_decoder(16#8b#)) OR
 					(reg_q850 AND symb_decoder(16#af#)) OR
 					(reg_q850 AND symb_decoder(16#98#)) OR
 					(reg_q850 AND symb_decoder(16#2a#)) OR
 					(reg_q850 AND symb_decoder(16#ea#)) OR
 					(reg_q850 AND symb_decoder(16#82#)) OR
 					(reg_q850 AND symb_decoder(16#66#)) OR
 					(reg_q850 AND symb_decoder(16#bf#)) OR
 					(reg_q850 AND symb_decoder(16#fd#)) OR
 					(reg_q850 AND symb_decoder(16#fe#)) OR
 					(reg_q850 AND symb_decoder(16#27#)) OR
 					(reg_q850 AND symb_decoder(16#61#)) OR
 					(reg_q850 AND symb_decoder(16#b9#)) OR
 					(reg_q850 AND symb_decoder(16#db#)) OR
 					(reg_q850 AND symb_decoder(16#a9#)) OR
 					(reg_q850 AND symb_decoder(16#a7#)) OR
 					(reg_q850 AND symb_decoder(16#e6#)) OR
 					(reg_q850 AND symb_decoder(16#f2#)) OR
 					(reg_q850 AND symb_decoder(16#f0#)) OR
 					(reg_q850 AND symb_decoder(16#de#)) OR
 					(reg_q850 AND symb_decoder(16#15#)) OR
 					(reg_q850 AND symb_decoder(16#43#)) OR
 					(reg_q850 AND symb_decoder(16#45#)) OR
 					(reg_q850 AND symb_decoder(16#4c#)) OR
 					(reg_q850 AND symb_decoder(16#d5#)) OR
 					(reg_q850 AND symb_decoder(16#9e#)) OR
 					(reg_q850 AND symb_decoder(16#9b#)) OR
 					(reg_q850 AND symb_decoder(16#63#)) OR
 					(reg_q850 AND symb_decoder(16#ef#)) OR
 					(reg_q850 AND symb_decoder(16#ba#)) OR
 					(reg_q850 AND symb_decoder(16#a8#)) OR
 					(reg_q850 AND symb_decoder(16#d6#)) OR
 					(reg_q850 AND symb_decoder(16#62#)) OR
 					(reg_q850 AND symb_decoder(16#1e#)) OR
 					(reg_q850 AND symb_decoder(16#df#)) OR
 					(reg_q850 AND symb_decoder(16#c9#)) OR
 					(reg_q850 AND symb_decoder(16#35#)) OR
 					(reg_q850 AND symb_decoder(16#7c#)) OR
 					(reg_q850 AND symb_decoder(16#5d#)) OR
 					(reg_q850 AND symb_decoder(16#dc#)) OR
 					(reg_q850 AND symb_decoder(16#ff#)) OR
 					(reg_q850 AND symb_decoder(16#39#)) OR
 					(reg_q850 AND symb_decoder(16#14#)) OR
 					(reg_q850 AND symb_decoder(16#87#)) OR
 					(reg_q850 AND symb_decoder(16#ce#)) OR
 					(reg_q850 AND symb_decoder(16#f7#)) OR
 					(reg_q850 AND symb_decoder(16#59#)) OR
 					(reg_q850 AND symb_decoder(16#ed#)) OR
 					(reg_q850 AND symb_decoder(16#f1#)) OR
 					(reg_q850 AND symb_decoder(16#f3#)) OR
 					(reg_q850 AND symb_decoder(16#4d#)) OR
 					(reg_q850 AND symb_decoder(16#ad#)) OR
 					(reg_q850 AND symb_decoder(16#71#)) OR
 					(reg_q850 AND symb_decoder(16#e8#)) OR
 					(reg_q850 AND symb_decoder(16#11#)) OR
 					(reg_q850 AND symb_decoder(16#b7#)) OR
 					(reg_q850 AND symb_decoder(16#f6#)) OR
 					(reg_q850 AND symb_decoder(16#6a#)) OR
 					(reg_q850 AND symb_decoder(16#44#)) OR
 					(reg_q850 AND symb_decoder(16#97#)) OR
 					(reg_q850 AND symb_decoder(16#70#)) OR
 					(reg_q850 AND symb_decoder(16#b1#)) OR
 					(reg_q850 AND symb_decoder(16#ab#)) OR
 					(reg_q850 AND symb_decoder(16#96#)) OR
 					(reg_q850 AND symb_decoder(16#e5#)) OR
 					(reg_q850 AND symb_decoder(16#da#)) OR
 					(reg_q850 AND symb_decoder(16#92#)) OR
 					(reg_q850 AND symb_decoder(16#8e#)) OR
 					(reg_q850 AND symb_decoder(16#c3#)) OR
 					(reg_q850 AND symb_decoder(16#57#)) OR
 					(reg_q850 AND symb_decoder(16#b3#)) OR
 					(reg_q850 AND symb_decoder(16#9a#)) OR
 					(reg_q850 AND symb_decoder(16#9d#)) OR
 					(reg_q850 AND symb_decoder(16#2b#)) OR
 					(reg_q850 AND symb_decoder(16#95#)) OR
 					(reg_q850 AND symb_decoder(16#25#));
reg_q850_init <= '0' ;
	p_reg_q850: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q850 <= reg_q850_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q850 <= reg_q850_init;
        else
          reg_q850 <= reg_q850_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1224_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1224 AND symb_decoder(16#a5#)) OR
 					(reg_q1224 AND symb_decoder(16#89#)) OR
 					(reg_q1224 AND symb_decoder(16#b7#)) OR
 					(reg_q1224 AND symb_decoder(16#14#)) OR
 					(reg_q1224 AND symb_decoder(16#fb#)) OR
 					(reg_q1224 AND symb_decoder(16#0d#)) OR
 					(reg_q1224 AND symb_decoder(16#22#)) OR
 					(reg_q1224 AND symb_decoder(16#60#)) OR
 					(reg_q1224 AND symb_decoder(16#ad#)) OR
 					(reg_q1224 AND symb_decoder(16#8b#)) OR
 					(reg_q1224 AND symb_decoder(16#18#)) OR
 					(reg_q1224 AND symb_decoder(16#fe#)) OR
 					(reg_q1224 AND symb_decoder(16#10#)) OR
 					(reg_q1224 AND symb_decoder(16#c1#)) OR
 					(reg_q1224 AND symb_decoder(16#bb#)) OR
 					(reg_q1224 AND symb_decoder(16#cf#)) OR
 					(reg_q1224 AND symb_decoder(16#de#)) OR
 					(reg_q1224 AND symb_decoder(16#bf#)) OR
 					(reg_q1224 AND symb_decoder(16#6d#)) OR
 					(reg_q1224 AND symb_decoder(16#46#)) OR
 					(reg_q1224 AND symb_decoder(16#85#)) OR
 					(reg_q1224 AND symb_decoder(16#01#)) OR
 					(reg_q1224 AND symb_decoder(16#86#)) OR
 					(reg_q1224 AND symb_decoder(16#e2#)) OR
 					(reg_q1224 AND symb_decoder(16#bc#)) OR
 					(reg_q1224 AND symb_decoder(16#4e#)) OR
 					(reg_q1224 AND symb_decoder(16#e6#)) OR
 					(reg_q1224 AND symb_decoder(16#1a#)) OR
 					(reg_q1224 AND symb_decoder(16#2d#)) OR
 					(reg_q1224 AND symb_decoder(16#a6#)) OR
 					(reg_q1224 AND symb_decoder(16#1e#)) OR
 					(reg_q1224 AND symb_decoder(16#a7#)) OR
 					(reg_q1224 AND symb_decoder(16#44#)) OR
 					(reg_q1224 AND symb_decoder(16#5c#)) OR
 					(reg_q1224 AND symb_decoder(16#00#)) OR
 					(reg_q1224 AND symb_decoder(16#c4#)) OR
 					(reg_q1224 AND symb_decoder(16#6b#)) OR
 					(reg_q1224 AND symb_decoder(16#d5#)) OR
 					(reg_q1224 AND symb_decoder(16#3f#)) OR
 					(reg_q1224 AND symb_decoder(16#d4#)) OR
 					(reg_q1224 AND symb_decoder(16#08#)) OR
 					(reg_q1224 AND symb_decoder(16#24#)) OR
 					(reg_q1224 AND symb_decoder(16#23#)) OR
 					(reg_q1224 AND symb_decoder(16#32#)) OR
 					(reg_q1224 AND symb_decoder(16#8f#)) OR
 					(reg_q1224 AND symb_decoder(16#40#)) OR
 					(reg_q1224 AND symb_decoder(16#bd#)) OR
 					(reg_q1224 AND symb_decoder(16#97#)) OR
 					(reg_q1224 AND symb_decoder(16#a1#)) OR
 					(reg_q1224 AND symb_decoder(16#09#)) OR
 					(reg_q1224 AND symb_decoder(16#12#)) OR
 					(reg_q1224 AND symb_decoder(16#39#)) OR
 					(reg_q1224 AND symb_decoder(16#dd#)) OR
 					(reg_q1224 AND symb_decoder(16#7f#)) OR
 					(reg_q1224 AND symb_decoder(16#b3#)) OR
 					(reg_q1224 AND symb_decoder(16#3b#)) OR
 					(reg_q1224 AND symb_decoder(16#f7#)) OR
 					(reg_q1224 AND symb_decoder(16#5d#)) OR
 					(reg_q1224 AND symb_decoder(16#da#)) OR
 					(reg_q1224 AND symb_decoder(16#95#)) OR
 					(reg_q1224 AND symb_decoder(16#ed#)) OR
 					(reg_q1224 AND symb_decoder(16#fa#)) OR
 					(reg_q1224 AND symb_decoder(16#5a#)) OR
 					(reg_q1224 AND symb_decoder(16#9c#)) OR
 					(reg_q1224 AND symb_decoder(16#19#)) OR
 					(reg_q1224 AND symb_decoder(16#eb#)) OR
 					(reg_q1224 AND symb_decoder(16#98#)) OR
 					(reg_q1224 AND symb_decoder(16#73#)) OR
 					(reg_q1224 AND symb_decoder(16#1d#)) OR
 					(reg_q1224 AND symb_decoder(16#9d#)) OR
 					(reg_q1224 AND symb_decoder(16#16#)) OR
 					(reg_q1224 AND symb_decoder(16#5e#)) OR
 					(reg_q1224 AND symb_decoder(16#83#)) OR
 					(reg_q1224 AND symb_decoder(16#96#)) OR
 					(reg_q1224 AND symb_decoder(16#e8#)) OR
 					(reg_q1224 AND symb_decoder(16#c0#)) OR
 					(reg_q1224 AND symb_decoder(16#f8#)) OR
 					(reg_q1224 AND symb_decoder(16#c2#)) OR
 					(reg_q1224 AND symb_decoder(16#4c#)) OR
 					(reg_q1224 AND symb_decoder(16#45#)) OR
 					(reg_q1224 AND symb_decoder(16#0a#)) OR
 					(reg_q1224 AND symb_decoder(16#74#)) OR
 					(reg_q1224 AND symb_decoder(16#aa#)) OR
 					(reg_q1224 AND symb_decoder(16#a9#)) OR
 					(reg_q1224 AND symb_decoder(16#c9#)) OR
 					(reg_q1224 AND symb_decoder(16#9e#)) OR
 					(reg_q1224 AND symb_decoder(16#02#)) OR
 					(reg_q1224 AND symb_decoder(16#76#)) OR
 					(reg_q1224 AND symb_decoder(16#59#)) OR
 					(reg_q1224 AND symb_decoder(16#72#)) OR
 					(reg_q1224 AND symb_decoder(16#ab#)) OR
 					(reg_q1224 AND symb_decoder(16#3d#)) OR
 					(reg_q1224 AND symb_decoder(16#94#)) OR
 					(reg_q1224 AND symb_decoder(16#df#)) OR
 					(reg_q1224 AND symb_decoder(16#78#)) OR
 					(reg_q1224 AND symb_decoder(16#e0#)) OR
 					(reg_q1224 AND symb_decoder(16#e1#)) OR
 					(reg_q1224 AND symb_decoder(16#ca#)) OR
 					(reg_q1224 AND symb_decoder(16#fc#)) OR
 					(reg_q1224 AND symb_decoder(16#13#)) OR
 					(reg_q1224 AND symb_decoder(16#57#)) OR
 					(reg_q1224 AND symb_decoder(16#43#)) OR
 					(reg_q1224 AND symb_decoder(16#61#)) OR
 					(reg_q1224 AND symb_decoder(16#7d#)) OR
 					(reg_q1224 AND symb_decoder(16#0b#)) OR
 					(reg_q1224 AND symb_decoder(16#9f#)) OR
 					(reg_q1224 AND symb_decoder(16#30#)) OR
 					(reg_q1224 AND symb_decoder(16#03#)) OR
 					(reg_q1224 AND symb_decoder(16#77#)) OR
 					(reg_q1224 AND symb_decoder(16#50#)) OR
 					(reg_q1224 AND symb_decoder(16#e7#)) OR
 					(reg_q1224 AND symb_decoder(16#67#)) OR
 					(reg_q1224 AND symb_decoder(16#ec#)) OR
 					(reg_q1224 AND symb_decoder(16#68#)) OR
 					(reg_q1224 AND symb_decoder(16#c8#)) OR
 					(reg_q1224 AND symb_decoder(16#b4#)) OR
 					(reg_q1224 AND symb_decoder(16#79#)) OR
 					(reg_q1224 AND symb_decoder(16#fd#)) OR
 					(reg_q1224 AND symb_decoder(16#cd#)) OR
 					(reg_q1224 AND symb_decoder(16#0f#)) OR
 					(reg_q1224 AND symb_decoder(16#d6#)) OR
 					(reg_q1224 AND symb_decoder(16#31#)) OR
 					(reg_q1224 AND symb_decoder(16#4b#)) OR
 					(reg_q1224 AND symb_decoder(16#36#)) OR
 					(reg_q1224 AND symb_decoder(16#0e#)) OR
 					(reg_q1224 AND symb_decoder(16#ea#)) OR
 					(reg_q1224 AND symb_decoder(16#75#)) OR
 					(reg_q1224 AND symb_decoder(16#dc#)) OR
 					(reg_q1224 AND symb_decoder(16#e5#)) OR
 					(reg_q1224 AND symb_decoder(16#41#)) OR
 					(reg_q1224 AND symb_decoder(16#f1#)) OR
 					(reg_q1224 AND symb_decoder(16#4f#)) OR
 					(reg_q1224 AND symb_decoder(16#69#)) OR
 					(reg_q1224 AND symb_decoder(16#2f#)) OR
 					(reg_q1224 AND symb_decoder(16#a0#)) OR
 					(reg_q1224 AND symb_decoder(16#8e#)) OR
 					(reg_q1224 AND symb_decoder(16#21#)) OR
 					(reg_q1224 AND symb_decoder(16#6f#)) OR
 					(reg_q1224 AND symb_decoder(16#8d#)) OR
 					(reg_q1224 AND symb_decoder(16#4d#)) OR
 					(reg_q1224 AND symb_decoder(16#d0#)) OR
 					(reg_q1224 AND symb_decoder(16#7c#)) OR
 					(reg_q1224 AND symb_decoder(16#1b#)) OR
 					(reg_q1224 AND symb_decoder(16#62#)) OR
 					(reg_q1224 AND symb_decoder(16#9b#)) OR
 					(reg_q1224 AND symb_decoder(16#cc#)) OR
 					(reg_q1224 AND symb_decoder(16#f6#)) OR
 					(reg_q1224 AND symb_decoder(16#25#)) OR
 					(reg_q1224 AND symb_decoder(16#17#)) OR
 					(reg_q1224 AND symb_decoder(16#71#)) OR
 					(reg_q1224 AND symb_decoder(16#07#)) OR
 					(reg_q1224 AND symb_decoder(16#4a#)) OR
 					(reg_q1224 AND symb_decoder(16#91#)) OR
 					(reg_q1224 AND symb_decoder(16#d1#)) OR
 					(reg_q1224 AND symb_decoder(16#15#)) OR
 					(reg_q1224 AND symb_decoder(16#b6#)) OR
 					(reg_q1224 AND symb_decoder(16#b9#)) OR
 					(reg_q1224 AND symb_decoder(16#80#)) OR
 					(reg_q1224 AND symb_decoder(16#87#)) OR
 					(reg_q1224 AND symb_decoder(16#04#)) OR
 					(reg_q1224 AND symb_decoder(16#28#)) OR
 					(reg_q1224 AND symb_decoder(16#1c#)) OR
 					(reg_q1224 AND symb_decoder(16#2a#)) OR
 					(reg_q1224 AND symb_decoder(16#35#)) OR
 					(reg_q1224 AND symb_decoder(16#2b#)) OR
 					(reg_q1224 AND symb_decoder(16#53#)) OR
 					(reg_q1224 AND symb_decoder(16#cb#)) OR
 					(reg_q1224 AND symb_decoder(16#2e#)) OR
 					(reg_q1224 AND symb_decoder(16#c7#)) OR
 					(reg_q1224 AND symb_decoder(16#ae#)) OR
 					(reg_q1224 AND symb_decoder(16#51#)) OR
 					(reg_q1224 AND symb_decoder(16#d7#)) OR
 					(reg_q1224 AND symb_decoder(16#9a#)) OR
 					(reg_q1224 AND symb_decoder(16#63#)) OR
 					(reg_q1224 AND symb_decoder(16#58#)) OR
 					(reg_q1224 AND symb_decoder(16#33#)) OR
 					(reg_q1224 AND symb_decoder(16#be#)) OR
 					(reg_q1224 AND symb_decoder(16#b0#)) OR
 					(reg_q1224 AND symb_decoder(16#47#)) OR
 					(reg_q1224 AND symb_decoder(16#7e#)) OR
 					(reg_q1224 AND symb_decoder(16#29#)) OR
 					(reg_q1224 AND symb_decoder(16#f2#)) OR
 					(reg_q1224 AND symb_decoder(16#3c#)) OR
 					(reg_q1224 AND symb_decoder(16#82#)) OR
 					(reg_q1224 AND symb_decoder(16#ff#)) OR
 					(reg_q1224 AND symb_decoder(16#3a#)) OR
 					(reg_q1224 AND symb_decoder(16#af#)) OR
 					(reg_q1224 AND symb_decoder(16#b1#)) OR
 					(reg_q1224 AND symb_decoder(16#65#)) OR
 					(reg_q1224 AND symb_decoder(16#0c#)) OR
 					(reg_q1224 AND symb_decoder(16#f9#)) OR
 					(reg_q1224 AND symb_decoder(16#b8#)) OR
 					(reg_q1224 AND symb_decoder(16#7a#)) OR
 					(reg_q1224 AND symb_decoder(16#c3#)) OR
 					(reg_q1224 AND symb_decoder(16#6e#)) OR
 					(reg_q1224 AND symb_decoder(16#55#)) OR
 					(reg_q1224 AND symb_decoder(16#92#)) OR
 					(reg_q1224 AND symb_decoder(16#7b#)) OR
 					(reg_q1224 AND symb_decoder(16#70#)) OR
 					(reg_q1224 AND symb_decoder(16#ce#)) OR
 					(reg_q1224 AND symb_decoder(16#ef#)) OR
 					(reg_q1224 AND symb_decoder(16#b5#)) OR
 					(reg_q1224 AND symb_decoder(16#db#)) OR
 					(reg_q1224 AND symb_decoder(16#ac#)) OR
 					(reg_q1224 AND symb_decoder(16#20#)) OR
 					(reg_q1224 AND symb_decoder(16#f4#)) OR
 					(reg_q1224 AND symb_decoder(16#f5#)) OR
 					(reg_q1224 AND symb_decoder(16#a8#)) OR
 					(reg_q1224 AND symb_decoder(16#54#)) OR
 					(reg_q1224 AND symb_decoder(16#2c#)) OR
 					(reg_q1224 AND symb_decoder(16#c5#)) OR
 					(reg_q1224 AND symb_decoder(16#1f#)) OR
 					(reg_q1224 AND symb_decoder(16#c6#)) OR
 					(reg_q1224 AND symb_decoder(16#56#)) OR
 					(reg_q1224 AND symb_decoder(16#d8#)) OR
 					(reg_q1224 AND symb_decoder(16#81#)) OR
 					(reg_q1224 AND symb_decoder(16#34#)) OR
 					(reg_q1224 AND symb_decoder(16#06#)) OR
 					(reg_q1224 AND symb_decoder(16#d2#)) OR
 					(reg_q1224 AND symb_decoder(16#a3#)) OR
 					(reg_q1224 AND symb_decoder(16#e9#)) OR
 					(reg_q1224 AND symb_decoder(16#5f#)) OR
 					(reg_q1224 AND symb_decoder(16#64#)) OR
 					(reg_q1224 AND symb_decoder(16#ba#)) OR
 					(reg_q1224 AND symb_decoder(16#e4#)) OR
 					(reg_q1224 AND symb_decoder(16#8a#)) OR
 					(reg_q1224 AND symb_decoder(16#37#)) OR
 					(reg_q1224 AND symb_decoder(16#6c#)) OR
 					(reg_q1224 AND symb_decoder(16#49#)) OR
 					(reg_q1224 AND symb_decoder(16#26#)) OR
 					(reg_q1224 AND symb_decoder(16#f3#)) OR
 					(reg_q1224 AND symb_decoder(16#ee#)) OR
 					(reg_q1224 AND symb_decoder(16#99#)) OR
 					(reg_q1224 AND symb_decoder(16#f0#)) OR
 					(reg_q1224 AND symb_decoder(16#52#)) OR
 					(reg_q1224 AND symb_decoder(16#27#)) OR
 					(reg_q1224 AND symb_decoder(16#b2#)) OR
 					(reg_q1224 AND symb_decoder(16#e3#)) OR
 					(reg_q1224 AND symb_decoder(16#93#)) OR
 					(reg_q1224 AND symb_decoder(16#d3#)) OR
 					(reg_q1224 AND symb_decoder(16#48#)) OR
 					(reg_q1224 AND symb_decoder(16#5b#)) OR
 					(reg_q1224 AND symb_decoder(16#11#)) OR
 					(reg_q1224 AND symb_decoder(16#42#)) OR
 					(reg_q1224 AND symb_decoder(16#38#)) OR
 					(reg_q1224 AND symb_decoder(16#66#)) OR
 					(reg_q1224 AND symb_decoder(16#8c#)) OR
 					(reg_q1224 AND symb_decoder(16#a2#)) OR
 					(reg_q1224 AND symb_decoder(16#6a#)) OR
 					(reg_q1224 AND symb_decoder(16#05#)) OR
 					(reg_q1224 AND symb_decoder(16#88#)) OR
 					(reg_q1224 AND symb_decoder(16#d9#)) OR
 					(reg_q1224 AND symb_decoder(16#3e#)) OR
 					(reg_q1224 AND symb_decoder(16#90#)) OR
 					(reg_q1224 AND symb_decoder(16#a4#)) OR
 					(reg_q1224 AND symb_decoder(16#84#));
reg_q1224_init <= '0' ;
	p_reg_q1224: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1224 <= reg_q1224_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1224 <= reg_q1224_init;
        else
          reg_q1224 <= reg_q1224_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q813_in <= (reg_q813 AND symb_decoder(16#9f#)) OR
 					(reg_q813 AND symb_decoder(16#ef#)) OR
 					(reg_q813 AND symb_decoder(16#43#)) OR
 					(reg_q813 AND symb_decoder(16#aa#)) OR
 					(reg_q813 AND symb_decoder(16#e5#)) OR
 					(reg_q813 AND symb_decoder(16#15#)) OR
 					(reg_q813 AND symb_decoder(16#f2#)) OR
 					(reg_q813 AND symb_decoder(16#23#)) OR
 					(reg_q813 AND symb_decoder(16#fa#)) OR
 					(reg_q813 AND symb_decoder(16#e1#)) OR
 					(reg_q813 AND symb_decoder(16#2b#)) OR
 					(reg_q813 AND symb_decoder(16#81#)) OR
 					(reg_q813 AND symb_decoder(16#eb#)) OR
 					(reg_q813 AND symb_decoder(16#9d#)) OR
 					(reg_q813 AND symb_decoder(16#40#)) OR
 					(reg_q813 AND symb_decoder(16#83#)) OR
 					(reg_q813 AND symb_decoder(16#87#)) OR
 					(reg_q813 AND symb_decoder(16#ce#)) OR
 					(reg_q813 AND symb_decoder(16#84#)) OR
 					(reg_q813 AND symb_decoder(16#ea#)) OR
 					(reg_q813 AND symb_decoder(16#bb#)) OR
 					(reg_q813 AND symb_decoder(16#95#)) OR
 					(reg_q813 AND symb_decoder(16#62#)) OR
 					(reg_q813 AND symb_decoder(16#18#)) OR
 					(reg_q813 AND symb_decoder(16#6d#)) OR
 					(reg_q813 AND symb_decoder(16#c5#)) OR
 					(reg_q813 AND symb_decoder(16#6f#)) OR
 					(reg_q813 AND symb_decoder(16#c8#)) OR
 					(reg_q813 AND symb_decoder(16#98#)) OR
 					(reg_q813 AND symb_decoder(16#a9#)) OR
 					(reg_q813 AND symb_decoder(16#c2#)) OR
 					(reg_q813 AND symb_decoder(16#3b#)) OR
 					(reg_q813 AND symb_decoder(16#74#)) OR
 					(reg_q813 AND symb_decoder(16#58#)) OR
 					(reg_q813 AND symb_decoder(16#4c#)) OR
 					(reg_q813 AND symb_decoder(16#28#)) OR
 					(reg_q813 AND symb_decoder(16#0e#)) OR
 					(reg_q813 AND symb_decoder(16#1a#)) OR
 					(reg_q813 AND symb_decoder(16#05#)) OR
 					(reg_q813 AND symb_decoder(16#f6#)) OR
 					(reg_q813 AND symb_decoder(16#30#)) OR
 					(reg_q813 AND symb_decoder(16#53#)) OR
 					(reg_q813 AND symb_decoder(16#ca#)) OR
 					(reg_q813 AND symb_decoder(16#26#)) OR
 					(reg_q813 AND symb_decoder(16#ed#)) OR
 					(reg_q813 AND symb_decoder(16#37#)) OR
 					(reg_q813 AND symb_decoder(16#42#)) OR
 					(reg_q813 AND symb_decoder(16#7a#)) OR
 					(reg_q813 AND symb_decoder(16#27#)) OR
 					(reg_q813 AND symb_decoder(16#51#)) OR
 					(reg_q813 AND symb_decoder(16#1e#)) OR
 					(reg_q813 AND symb_decoder(16#2d#)) OR
 					(reg_q813 AND symb_decoder(16#24#)) OR
 					(reg_q813 AND symb_decoder(16#9c#)) OR
 					(reg_q813 AND symb_decoder(16#4a#)) OR
 					(reg_q813 AND symb_decoder(16#54#)) OR
 					(reg_q813 AND symb_decoder(16#72#)) OR
 					(reg_q813 AND symb_decoder(16#5e#)) OR
 					(reg_q813 AND symb_decoder(16#b1#)) OR
 					(reg_q813 AND symb_decoder(16#19#)) OR
 					(reg_q813 AND symb_decoder(16#1b#)) OR
 					(reg_q813 AND symb_decoder(16#2c#)) OR
 					(reg_q813 AND symb_decoder(16#b6#)) OR
 					(reg_q813 AND symb_decoder(16#97#)) OR
 					(reg_q813 AND symb_decoder(16#20#)) OR
 					(reg_q813 AND symb_decoder(16#e3#)) OR
 					(reg_q813 AND symb_decoder(16#5a#)) OR
 					(reg_q813 AND symb_decoder(16#cb#)) OR
 					(reg_q813 AND symb_decoder(16#bd#)) OR
 					(reg_q813 AND symb_decoder(16#08#)) OR
 					(reg_q813 AND symb_decoder(16#5f#)) OR
 					(reg_q813 AND symb_decoder(16#49#)) OR
 					(reg_q813 AND symb_decoder(16#96#)) OR
 					(reg_q813 AND symb_decoder(16#d5#)) OR
 					(reg_q813 AND symb_decoder(16#9e#)) OR
 					(reg_q813 AND symb_decoder(16#1d#)) OR
 					(reg_q813 AND symb_decoder(16#29#)) OR
 					(reg_q813 AND symb_decoder(16#7f#)) OR
 					(reg_q813 AND symb_decoder(16#d3#)) OR
 					(reg_q813 AND symb_decoder(16#c7#)) OR
 					(reg_q813 AND symb_decoder(16#70#)) OR
 					(reg_q813 AND symb_decoder(16#44#)) OR
 					(reg_q813 AND symb_decoder(16#47#)) OR
 					(reg_q813 AND symb_decoder(16#df#)) OR
 					(reg_q813 AND symb_decoder(16#c9#)) OR
 					(reg_q813 AND symb_decoder(16#a6#)) OR
 					(reg_q813 AND symb_decoder(16#f4#)) OR
 					(reg_q813 AND symb_decoder(16#6c#)) OR
 					(reg_q813 AND symb_decoder(16#5c#)) OR
 					(reg_q813 AND symb_decoder(16#bf#)) OR
 					(reg_q813 AND symb_decoder(16#cc#)) OR
 					(reg_q813 AND symb_decoder(16#f7#)) OR
 					(reg_q813 AND symb_decoder(16#85#)) OR
 					(reg_q813 AND symb_decoder(16#2a#)) OR
 					(reg_q813 AND symb_decoder(16#9b#)) OR
 					(reg_q813 AND symb_decoder(16#73#)) OR
 					(reg_q813 AND symb_decoder(16#a2#)) OR
 					(reg_q813 AND symb_decoder(16#5d#)) OR
 					(reg_q813 AND symb_decoder(16#65#)) OR
 					(reg_q813 AND symb_decoder(16#56#)) OR
 					(reg_q813 AND symb_decoder(16#21#)) OR
 					(reg_q813 AND symb_decoder(16#17#)) OR
 					(reg_q813 AND symb_decoder(16#68#)) OR
 					(reg_q813 AND symb_decoder(16#b9#)) OR
 					(reg_q813 AND symb_decoder(16#89#)) OR
 					(reg_q813 AND symb_decoder(16#db#)) OR
 					(reg_q813 AND symb_decoder(16#11#)) OR
 					(reg_q813 AND symb_decoder(16#bc#)) OR
 					(reg_q813 AND symb_decoder(16#80#)) OR
 					(reg_q813 AND symb_decoder(16#8a#)) OR
 					(reg_q813 AND symb_decoder(16#64#)) OR
 					(reg_q813 AND symb_decoder(16#07#)) OR
 					(reg_q813 AND symb_decoder(16#de#)) OR
 					(reg_q813 AND symb_decoder(16#f9#)) OR
 					(reg_q813 AND symb_decoder(16#79#)) OR
 					(reg_q813 AND symb_decoder(16#34#)) OR
 					(reg_q813 AND symb_decoder(16#76#)) OR
 					(reg_q813 AND symb_decoder(16#d9#)) OR
 					(reg_q813 AND symb_decoder(16#60#)) OR
 					(reg_q813 AND symb_decoder(16#75#)) OR
 					(reg_q813 AND symb_decoder(16#a3#)) OR
 					(reg_q813 AND symb_decoder(16#03#)) OR
 					(reg_q813 AND symb_decoder(16#d4#)) OR
 					(reg_q813 AND symb_decoder(16#b2#)) OR
 					(reg_q813 AND symb_decoder(16#02#)) OR
 					(reg_q813 AND symb_decoder(16#b4#)) OR
 					(reg_q813 AND symb_decoder(16#01#)) OR
 					(reg_q813 AND symb_decoder(16#0c#)) OR
 					(reg_q813 AND symb_decoder(16#93#)) OR
 					(reg_q813 AND symb_decoder(16#e6#)) OR
 					(reg_q813 AND symb_decoder(16#61#)) OR
 					(reg_q813 AND symb_decoder(16#e9#)) OR
 					(reg_q813 AND symb_decoder(16#86#)) OR
 					(reg_q813 AND symb_decoder(16#50#)) OR
 					(reg_q813 AND symb_decoder(16#e8#)) OR
 					(reg_q813 AND symb_decoder(16#22#)) OR
 					(reg_q813 AND symb_decoder(16#46#)) OR
 					(reg_q813 AND symb_decoder(16#f0#)) OR
 					(reg_q813 AND symb_decoder(16#e7#)) OR
 					(reg_q813 AND symb_decoder(16#1f#)) OR
 					(reg_q813 AND symb_decoder(16#4d#)) OR
 					(reg_q813 AND symb_decoder(16#3d#)) OR
 					(reg_q813 AND symb_decoder(16#88#)) OR
 					(reg_q813 AND symb_decoder(16#25#)) OR
 					(reg_q813 AND symb_decoder(16#3a#)) OR
 					(reg_q813 AND symb_decoder(16#69#)) OR
 					(reg_q813 AND symb_decoder(16#4f#)) OR
 					(reg_q813 AND symb_decoder(16#fb#)) OR
 					(reg_q813 AND symb_decoder(16#ba#)) OR
 					(reg_q813 AND symb_decoder(16#94#)) OR
 					(reg_q813 AND symb_decoder(16#ab#)) OR
 					(reg_q813 AND symb_decoder(16#52#)) OR
 					(reg_q813 AND symb_decoder(16#7d#)) OR
 					(reg_q813 AND symb_decoder(16#38#)) OR
 					(reg_q813 AND symb_decoder(16#6a#)) OR
 					(reg_q813 AND symb_decoder(16#77#)) OR
 					(reg_q813 AND symb_decoder(16#c1#)) OR
 					(reg_q813 AND symb_decoder(16#1c#)) OR
 					(reg_q813 AND symb_decoder(16#0f#)) OR
 					(reg_q813 AND symb_decoder(16#8f#)) OR
 					(reg_q813 AND symb_decoder(16#c6#)) OR
 					(reg_q813 AND symb_decoder(16#b7#)) OR
 					(reg_q813 AND symb_decoder(16#8c#)) OR
 					(reg_q813 AND symb_decoder(16#a5#)) OR
 					(reg_q813 AND symb_decoder(16#09#)) OR
 					(reg_q813 AND symb_decoder(16#71#)) OR
 					(reg_q813 AND symb_decoder(16#63#)) OR
 					(reg_q813 AND symb_decoder(16#af#)) OR
 					(reg_q813 AND symb_decoder(16#3e#)) OR
 					(reg_q813 AND symb_decoder(16#ec#)) OR
 					(reg_q813 AND symb_decoder(16#6b#)) OR
 					(reg_q813 AND symb_decoder(16#13#)) OR
 					(reg_q813 AND symb_decoder(16#39#)) OR
 					(reg_q813 AND symb_decoder(16#33#)) OR
 					(reg_q813 AND symb_decoder(16#90#)) OR
 					(reg_q813 AND symb_decoder(16#d6#)) OR
 					(reg_q813 AND symb_decoder(16#7c#)) OR
 					(reg_q813 AND symb_decoder(16#e4#)) OR
 					(reg_q813 AND symb_decoder(16#5b#)) OR
 					(reg_q813 AND symb_decoder(16#66#)) OR
 					(reg_q813 AND symb_decoder(16#ae#)) OR
 					(reg_q813 AND symb_decoder(16#41#)) OR
 					(reg_q813 AND symb_decoder(16#14#)) OR
 					(reg_q813 AND symb_decoder(16#ee#)) OR
 					(reg_q813 AND symb_decoder(16#d2#)) OR
 					(reg_q813 AND symb_decoder(16#f8#)) OR
 					(reg_q813 AND symb_decoder(16#91#)) OR
 					(reg_q813 AND symb_decoder(16#78#)) OR
 					(reg_q813 AND symb_decoder(16#ff#)) OR
 					(reg_q813 AND symb_decoder(16#10#)) OR
 					(reg_q813 AND symb_decoder(16#a4#)) OR
 					(reg_q813 AND symb_decoder(16#2f#)) OR
 					(reg_q813 AND symb_decoder(16#fe#)) OR
 					(reg_q813 AND symb_decoder(16#b8#)) OR
 					(reg_q813 AND symb_decoder(16#be#)) OR
 					(reg_q813 AND symb_decoder(16#99#)) OR
 					(reg_q813 AND symb_decoder(16#3c#)) OR
 					(reg_q813 AND symb_decoder(16#0b#)) OR
 					(reg_q813 AND symb_decoder(16#f3#)) OR
 					(reg_q813 AND symb_decoder(16#a1#)) OR
 					(reg_q813 AND symb_decoder(16#b0#)) OR
 					(reg_q813 AND symb_decoder(16#8d#)) OR
 					(reg_q813 AND symb_decoder(16#f5#)) OR
 					(reg_q813 AND symb_decoder(16#d8#)) OR
 					(reg_q813 AND symb_decoder(16#cf#)) OR
 					(reg_q813 AND symb_decoder(16#d0#)) OR
 					(reg_q813 AND symb_decoder(16#31#)) OR
 					(reg_q813 AND symb_decoder(16#c0#)) OR
 					(reg_q813 AND symb_decoder(16#dd#)) OR
 					(reg_q813 AND symb_decoder(16#a7#)) OR
 					(reg_q813 AND symb_decoder(16#a0#)) OR
 					(reg_q813 AND symb_decoder(16#c3#)) OR
 					(reg_q813 AND symb_decoder(16#7e#)) OR
 					(reg_q813 AND symb_decoder(16#12#)) OR
 					(reg_q813 AND symb_decoder(16#8b#)) OR
 					(reg_q813 AND symb_decoder(16#b5#)) OR
 					(reg_q813 AND symb_decoder(16#a8#)) OR
 					(reg_q813 AND symb_decoder(16#e2#)) OR
 					(reg_q813 AND symb_decoder(16#04#)) OR
 					(reg_q813 AND symb_decoder(16#67#)) OR
 					(reg_q813 AND symb_decoder(16#7b#)) OR
 					(reg_q813 AND symb_decoder(16#00#)) OR
 					(reg_q813 AND symb_decoder(16#36#)) OR
 					(reg_q813 AND symb_decoder(16#ad#)) OR
 					(reg_q813 AND symb_decoder(16#e0#)) OR
 					(reg_q813 AND symb_decoder(16#45#)) OR
 					(reg_q813 AND symb_decoder(16#16#)) OR
 					(reg_q813 AND symb_decoder(16#55#)) OR
 					(reg_q813 AND symb_decoder(16#da#)) OR
 					(reg_q813 AND symb_decoder(16#4b#)) OR
 					(reg_q813 AND symb_decoder(16#35#)) OR
 					(reg_q813 AND symb_decoder(16#3f#)) OR
 					(reg_q813 AND symb_decoder(16#fc#)) OR
 					(reg_q813 AND symb_decoder(16#48#)) OR
 					(reg_q813 AND symb_decoder(16#ac#)) OR
 					(reg_q813 AND symb_decoder(16#c4#)) OR
 					(reg_q813 AND symb_decoder(16#59#)) OR
 					(reg_q813 AND symb_decoder(16#d1#)) OR
 					(reg_q813 AND symb_decoder(16#32#)) OR
 					(reg_q813 AND symb_decoder(16#92#)) OR
 					(reg_q813 AND symb_decoder(16#06#)) OR
 					(reg_q813 AND symb_decoder(16#fd#)) OR
 					(reg_q813 AND symb_decoder(16#4e#)) OR
 					(reg_q813 AND symb_decoder(16#f1#)) OR
 					(reg_q813 AND symb_decoder(16#d7#)) OR
 					(reg_q813 AND symb_decoder(16#82#)) OR
 					(reg_q813 AND symb_decoder(16#b3#)) OR
 					(reg_q813 AND symb_decoder(16#6e#)) OR
 					(reg_q813 AND symb_decoder(16#57#)) OR
 					(reg_q813 AND symb_decoder(16#8e#)) OR
 					(reg_q813 AND symb_decoder(16#9a#)) OR
 					(reg_q813 AND symb_decoder(16#cd#)) OR
 					(reg_q813 AND symb_decoder(16#dc#)) OR
 					(reg_q813 AND symb_decoder(16#2e#)) OR
 					(reg_q791 AND symb_decoder(16#3f#)) OR
 					(reg_q791 AND symb_decoder(16#c4#)) OR
 					(reg_q791 AND symb_decoder(16#51#)) OR
 					(reg_q791 AND symb_decoder(16#f8#)) OR
 					(reg_q791 AND symb_decoder(16#46#)) OR
 					(reg_q791 AND symb_decoder(16#df#)) OR
 					(reg_q791 AND symb_decoder(16#1b#)) OR
 					(reg_q791 AND symb_decoder(16#85#)) OR
 					(reg_q791 AND symb_decoder(16#01#)) OR
 					(reg_q791 AND symb_decoder(16#62#)) OR
 					(reg_q791 AND symb_decoder(16#90#)) OR
 					(reg_q791 AND symb_decoder(16#94#)) OR
 					(reg_q791 AND symb_decoder(16#5f#)) OR
 					(reg_q791 AND symb_decoder(16#5c#)) OR
 					(reg_q791 AND symb_decoder(16#7a#)) OR
 					(reg_q791 AND symb_decoder(16#9d#)) OR
 					(reg_q791 AND symb_decoder(16#ef#)) OR
 					(reg_q791 AND symb_decoder(16#96#)) OR
 					(reg_q791 AND symb_decoder(16#bc#)) OR
 					(reg_q791 AND symb_decoder(16#ab#)) OR
 					(reg_q791 AND symb_decoder(16#3c#)) OR
 					(reg_q791 AND symb_decoder(16#fe#)) OR
 					(reg_q791 AND symb_decoder(16#07#)) OR
 					(reg_q791 AND symb_decoder(16#bd#)) OR
 					(reg_q791 AND symb_decoder(16#61#)) OR
 					(reg_q791 AND symb_decoder(16#8b#)) OR
 					(reg_q791 AND symb_decoder(16#f7#)) OR
 					(reg_q791 AND symb_decoder(16#37#)) OR
 					(reg_q791 AND symb_decoder(16#2d#)) OR
 					(reg_q791 AND symb_decoder(16#15#)) OR
 					(reg_q791 AND symb_decoder(16#7e#)) OR
 					(reg_q791 AND symb_decoder(16#1f#)) OR
 					(reg_q791 AND symb_decoder(16#59#)) OR
 					(reg_q791 AND symb_decoder(16#d2#)) OR
 					(reg_q791 AND symb_decoder(16#92#)) OR
 					(reg_q791 AND symb_decoder(16#28#)) OR
 					(reg_q791 AND symb_decoder(16#4e#)) OR
 					(reg_q791 AND symb_decoder(16#88#)) OR
 					(reg_q791 AND symb_decoder(16#6a#)) OR
 					(reg_q791 AND symb_decoder(16#78#)) OR
 					(reg_q791 AND symb_decoder(16#38#)) OR
 					(reg_q791 AND symb_decoder(16#5a#)) OR
 					(reg_q791 AND symb_decoder(16#3b#)) OR
 					(reg_q791 AND symb_decoder(16#7c#)) OR
 					(reg_q791 AND symb_decoder(16#d7#)) OR
 					(reg_q791 AND symb_decoder(16#4d#)) OR
 					(reg_q791 AND symb_decoder(16#e5#)) OR
 					(reg_q791 AND symb_decoder(16#06#)) OR
 					(reg_q791 AND symb_decoder(16#0e#)) OR
 					(reg_q791 AND symb_decoder(16#fa#)) OR
 					(reg_q791 AND symb_decoder(16#f1#)) OR
 					(reg_q791 AND symb_decoder(16#69#)) OR
 					(reg_q791 AND symb_decoder(16#4c#)) OR
 					(reg_q791 AND symb_decoder(16#f9#)) OR
 					(reg_q791 AND symb_decoder(16#54#)) OR
 					(reg_q791 AND symb_decoder(16#19#)) OR
 					(reg_q791 AND symb_decoder(16#7f#)) OR
 					(reg_q791 AND symb_decoder(16#f3#)) OR
 					(reg_q791 AND symb_decoder(16#00#)) OR
 					(reg_q791 AND symb_decoder(16#db#)) OR
 					(reg_q791 AND symb_decoder(16#10#)) OR
 					(reg_q791 AND symb_decoder(16#6f#)) OR
 					(reg_q791 AND symb_decoder(16#64#)) OR
 					(reg_q791 AND symb_decoder(16#af#)) OR
 					(reg_q791 AND symb_decoder(16#ec#)) OR
 					(reg_q791 AND symb_decoder(16#4a#)) OR
 					(reg_q791 AND symb_decoder(16#d3#)) OR
 					(reg_q791 AND symb_decoder(16#93#)) OR
 					(reg_q791 AND symb_decoder(16#a4#)) OR
 					(reg_q791 AND symb_decoder(16#30#)) OR
 					(reg_q791 AND symb_decoder(16#de#)) OR
 					(reg_q791 AND symb_decoder(16#14#)) OR
 					(reg_q791 AND symb_decoder(16#1e#)) OR
 					(reg_q791 AND symb_decoder(16#1a#)) OR
 					(reg_q791 AND symb_decoder(16#77#)) OR
 					(reg_q791 AND symb_decoder(16#d0#)) OR
 					(reg_q791 AND symb_decoder(16#20#)) OR
 					(reg_q791 AND symb_decoder(16#a7#)) OR
 					(reg_q791 AND symb_decoder(16#41#)) OR
 					(reg_q791 AND symb_decoder(16#68#)) OR
 					(reg_q791 AND symb_decoder(16#25#)) OR
 					(reg_q791 AND symb_decoder(16#57#)) OR
 					(reg_q791 AND symb_decoder(16#5b#)) OR
 					(reg_q791 AND symb_decoder(16#56#)) OR
 					(reg_q791 AND symb_decoder(16#ca#)) OR
 					(reg_q791 AND symb_decoder(16#2c#)) OR
 					(reg_q791 AND symb_decoder(16#03#)) OR
 					(reg_q791 AND symb_decoder(16#09#)) OR
 					(reg_q791 AND symb_decoder(16#2b#)) OR
 					(reg_q791 AND symb_decoder(16#67#)) OR
 					(reg_q791 AND symb_decoder(16#95#)) OR
 					(reg_q791 AND symb_decoder(16#c9#)) OR
 					(reg_q791 AND symb_decoder(16#e7#)) OR
 					(reg_q791 AND symb_decoder(16#97#)) OR
 					(reg_q791 AND symb_decoder(16#e0#)) OR
 					(reg_q791 AND symb_decoder(16#f0#)) OR
 					(reg_q791 AND symb_decoder(16#79#)) OR
 					(reg_q791 AND symb_decoder(16#11#)) OR
 					(reg_q791 AND symb_decoder(16#02#)) OR
 					(reg_q791 AND symb_decoder(16#0c#)) OR
 					(reg_q791 AND symb_decoder(16#39#)) OR
 					(reg_q791 AND symb_decoder(16#8a#)) OR
 					(reg_q791 AND symb_decoder(16#a1#)) OR
 					(reg_q791 AND symb_decoder(16#6e#)) OR
 					(reg_q791 AND symb_decoder(16#b2#)) OR
 					(reg_q791 AND symb_decoder(16#12#)) OR
 					(reg_q791 AND symb_decoder(16#b1#)) OR
 					(reg_q791 AND symb_decoder(16#74#)) OR
 					(reg_q791 AND symb_decoder(16#b5#)) OR
 					(reg_q791 AND symb_decoder(16#99#)) OR
 					(reg_q791 AND symb_decoder(16#ac#)) OR
 					(reg_q791 AND symb_decoder(16#24#)) OR
 					(reg_q791 AND symb_decoder(16#ae#)) OR
 					(reg_q791 AND symb_decoder(16#eb#)) OR
 					(reg_q791 AND symb_decoder(16#a8#)) OR
 					(reg_q791 AND symb_decoder(16#c0#)) OR
 					(reg_q791 AND symb_decoder(16#45#)) OR
 					(reg_q791 AND symb_decoder(16#13#)) OR
 					(reg_q791 AND symb_decoder(16#b0#)) OR
 					(reg_q791 AND symb_decoder(16#9c#)) OR
 					(reg_q791 AND symb_decoder(16#9f#)) OR
 					(reg_q791 AND symb_decoder(16#29#)) OR
 					(reg_q791 AND symb_decoder(16#cc#)) OR
 					(reg_q791 AND symb_decoder(16#5d#)) OR
 					(reg_q791 AND symb_decoder(16#aa#)) OR
 					(reg_q791 AND symb_decoder(16#ce#)) OR
 					(reg_q791 AND symb_decoder(16#42#)) OR
 					(reg_q791 AND symb_decoder(16#bb#)) OR
 					(reg_q791 AND symb_decoder(16#bf#)) OR
 					(reg_q791 AND symb_decoder(16#43#)) OR
 					(reg_q791 AND symb_decoder(16#cb#)) OR
 					(reg_q791 AND symb_decoder(16#8d#)) OR
 					(reg_q791 AND symb_decoder(16#5e#)) OR
 					(reg_q791 AND symb_decoder(16#c3#)) OR
 					(reg_q791 AND symb_decoder(16#80#)) OR
 					(reg_q791 AND symb_decoder(16#83#)) OR
 					(reg_q791 AND symb_decoder(16#f4#)) OR
 					(reg_q791 AND symb_decoder(16#b9#)) OR
 					(reg_q791 AND symb_decoder(16#c7#)) OR
 					(reg_q791 AND symb_decoder(16#c8#)) OR
 					(reg_q791 AND symb_decoder(16#d6#)) OR
 					(reg_q791 AND symb_decoder(16#be#)) OR
 					(reg_q791 AND symb_decoder(16#e4#)) OR
 					(reg_q791 AND symb_decoder(16#75#)) OR
 					(reg_q791 AND symb_decoder(16#87#)) OR
 					(reg_q791 AND symb_decoder(16#dd#)) OR
 					(reg_q791 AND symb_decoder(16#55#)) OR
 					(reg_q791 AND symb_decoder(16#cf#)) OR
 					(reg_q791 AND symb_decoder(16#b3#)) OR
 					(reg_q791 AND symb_decoder(16#7d#)) OR
 					(reg_q791 AND symb_decoder(16#86#)) OR
 					(reg_q791 AND symb_decoder(16#d8#)) OR
 					(reg_q791 AND symb_decoder(16#6d#)) OR
 					(reg_q791 AND symb_decoder(16#22#)) OR
 					(reg_q791 AND symb_decoder(16#27#)) OR
 					(reg_q791 AND symb_decoder(16#32#)) OR
 					(reg_q791 AND symb_decoder(16#9e#)) OR
 					(reg_q791 AND symb_decoder(16#7b#)) OR
 					(reg_q791 AND symb_decoder(16#21#)) OR
 					(reg_q791 AND symb_decoder(16#53#)) OR
 					(reg_q791 AND symb_decoder(16#08#)) OR
 					(reg_q791 AND symb_decoder(16#ea#)) OR
 					(reg_q791 AND symb_decoder(16#91#)) OR
 					(reg_q791 AND symb_decoder(16#d9#)) OR
 					(reg_q791 AND symb_decoder(16#2a#)) OR
 					(reg_q791 AND symb_decoder(16#c6#)) OR
 					(reg_q791 AND symb_decoder(16#81#)) OR
 					(reg_q791 AND symb_decoder(16#8e#)) OR
 					(reg_q791 AND symb_decoder(16#ff#)) OR
 					(reg_q791 AND symb_decoder(16#a5#)) OR
 					(reg_q791 AND symb_decoder(16#47#)) OR
 					(reg_q791 AND symb_decoder(16#44#)) OR
 					(reg_q791 AND symb_decoder(16#fb#)) OR
 					(reg_q791 AND symb_decoder(16#2f#)) OR
 					(reg_q791 AND symb_decoder(16#72#)) OR
 					(reg_q791 AND symb_decoder(16#c1#)) OR
 					(reg_q791 AND symb_decoder(16#ee#)) OR
 					(reg_q791 AND symb_decoder(16#17#)) OR
 					(reg_q791 AND symb_decoder(16#1c#)) OR
 					(reg_q791 AND symb_decoder(16#e1#)) OR
 					(reg_q791 AND symb_decoder(16#d4#)) OR
 					(reg_q791 AND symb_decoder(16#82#)) OR
 					(reg_q791 AND symb_decoder(16#04#)) OR
 					(reg_q791 AND symb_decoder(16#1d#)) OR
 					(reg_q791 AND symb_decoder(16#0f#)) OR
 					(reg_q791 AND symb_decoder(16#6c#)) OR
 					(reg_q791 AND symb_decoder(16#a6#)) OR
 					(reg_q791 AND symb_decoder(16#63#)) OR
 					(reg_q791 AND symb_decoder(16#b8#)) OR
 					(reg_q791 AND symb_decoder(16#70#)) OR
 					(reg_q791 AND symb_decoder(16#8c#)) OR
 					(reg_q791 AND symb_decoder(16#ba#)) OR
 					(reg_q791 AND symb_decoder(16#05#)) OR
 					(reg_q791 AND symb_decoder(16#34#)) OR
 					(reg_q791 AND symb_decoder(16#cd#)) OR
 					(reg_q791 AND symb_decoder(16#58#)) OR
 					(reg_q791 AND symb_decoder(16#e2#)) OR
 					(reg_q791 AND symb_decoder(16#52#)) OR
 					(reg_q791 AND symb_decoder(16#e8#)) OR
 					(reg_q791 AND symb_decoder(16#4b#)) OR
 					(reg_q791 AND symb_decoder(16#c5#)) OR
 					(reg_q791 AND symb_decoder(16#d5#)) OR
 					(reg_q791 AND symb_decoder(16#76#)) OR
 					(reg_q791 AND symb_decoder(16#35#)) OR
 					(reg_q791 AND symb_decoder(16#a2#)) OR
 					(reg_q791 AND symb_decoder(16#9a#)) OR
 					(reg_q791 AND symb_decoder(16#49#)) OR
 					(reg_q791 AND symb_decoder(16#60#)) OR
 					(reg_q791 AND symb_decoder(16#23#)) OR
 					(reg_q791 AND symb_decoder(16#b7#)) OR
 					(reg_q791 AND symb_decoder(16#dc#)) OR
 					(reg_q791 AND symb_decoder(16#89#)) OR
 					(reg_q791 AND symb_decoder(16#c2#)) OR
 					(reg_q791 AND symb_decoder(16#73#)) OR
 					(reg_q791 AND symb_decoder(16#3d#)) OR
 					(reg_q791 AND symb_decoder(16#16#)) OR
 					(reg_q791 AND symb_decoder(16#31#)) OR
 					(reg_q791 AND symb_decoder(16#e3#)) OR
 					(reg_q791 AND symb_decoder(16#a9#)) OR
 					(reg_q791 AND symb_decoder(16#e6#)) OR
 					(reg_q791 AND symb_decoder(16#e9#)) OR
 					(reg_q791 AND symb_decoder(16#36#)) OR
 					(reg_q791 AND symb_decoder(16#33#)) OR
 					(reg_q791 AND symb_decoder(16#fc#)) OR
 					(reg_q791 AND symb_decoder(16#2e#)) OR
 					(reg_q791 AND symb_decoder(16#8f#)) OR
 					(reg_q791 AND symb_decoder(16#ed#)) OR
 					(reg_q791 AND symb_decoder(16#ad#)) OR
 					(reg_q791 AND symb_decoder(16#f5#)) OR
 					(reg_q791 AND symb_decoder(16#3a#)) OR
 					(reg_q791 AND symb_decoder(16#84#)) OR
 					(reg_q791 AND symb_decoder(16#d1#)) OR
 					(reg_q791 AND symb_decoder(16#b4#)) OR
 					(reg_q791 AND symb_decoder(16#9b#)) OR
 					(reg_q791 AND symb_decoder(16#0b#)) OR
 					(reg_q791 AND symb_decoder(16#a0#)) OR
 					(reg_q791 AND symb_decoder(16#40#)) OR
 					(reg_q791 AND symb_decoder(16#4f#)) OR
 					(reg_q791 AND symb_decoder(16#48#)) OR
 					(reg_q791 AND symb_decoder(16#da#)) OR
 					(reg_q791 AND symb_decoder(16#66#)) OR
 					(reg_q791 AND symb_decoder(16#a3#)) OR
 					(reg_q791 AND symb_decoder(16#98#)) OR
 					(reg_q791 AND symb_decoder(16#fd#)) OR
 					(reg_q791 AND symb_decoder(16#f2#)) OR
 					(reg_q791 AND symb_decoder(16#3e#)) OR
 					(reg_q791 AND symb_decoder(16#18#)) OR
 					(reg_q791 AND symb_decoder(16#71#)) OR
 					(reg_q791 AND symb_decoder(16#f6#)) OR
 					(reg_q791 AND symb_decoder(16#6b#)) OR
 					(reg_q791 AND symb_decoder(16#b6#)) OR
 					(reg_q791 AND symb_decoder(16#50#)) OR
 					(reg_q791 AND symb_decoder(16#65#)) OR
 					(reg_q791 AND symb_decoder(16#26#));
reg_q813_init <= '0' ;
	p_reg_q813: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q813 <= reg_q813_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q813 <= reg_q813_init;
        else
          reg_q813 <= reg_q813_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2000_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2000 AND symb_decoder(16#e2#)) OR
 					(reg_q2000 AND symb_decoder(16#19#)) OR
 					(reg_q2000 AND symb_decoder(16#9b#)) OR
 					(reg_q2000 AND symb_decoder(16#56#)) OR
 					(reg_q2000 AND symb_decoder(16#9e#)) OR
 					(reg_q2000 AND symb_decoder(16#f4#)) OR
 					(reg_q2000 AND symb_decoder(16#e7#)) OR
 					(reg_q2000 AND symb_decoder(16#9f#)) OR
 					(reg_q2000 AND symb_decoder(16#ff#)) OR
 					(reg_q2000 AND symb_decoder(16#4a#)) OR
 					(reg_q2000 AND symb_decoder(16#0e#)) OR
 					(reg_q2000 AND symb_decoder(16#c0#)) OR
 					(reg_q2000 AND symb_decoder(16#70#)) OR
 					(reg_q2000 AND symb_decoder(16#e8#)) OR
 					(reg_q2000 AND symb_decoder(16#84#)) OR
 					(reg_q2000 AND symb_decoder(16#27#)) OR
 					(reg_q2000 AND symb_decoder(16#c1#)) OR
 					(reg_q2000 AND symb_decoder(16#09#)) OR
 					(reg_q2000 AND symb_decoder(16#e6#)) OR
 					(reg_q2000 AND symb_decoder(16#26#)) OR
 					(reg_q2000 AND symb_decoder(16#2f#)) OR
 					(reg_q2000 AND symb_decoder(16#63#)) OR
 					(reg_q2000 AND symb_decoder(16#6c#)) OR
 					(reg_q2000 AND symb_decoder(16#98#)) OR
 					(reg_q2000 AND symb_decoder(16#35#)) OR
 					(reg_q2000 AND symb_decoder(16#21#)) OR
 					(reg_q2000 AND symb_decoder(16#b5#)) OR
 					(reg_q2000 AND symb_decoder(16#d7#)) OR
 					(reg_q2000 AND symb_decoder(16#1d#)) OR
 					(reg_q2000 AND symb_decoder(16#a9#)) OR
 					(reg_q2000 AND symb_decoder(16#f6#)) OR
 					(reg_q2000 AND symb_decoder(16#5c#)) OR
 					(reg_q2000 AND symb_decoder(16#f1#)) OR
 					(reg_q2000 AND symb_decoder(16#53#)) OR
 					(reg_q2000 AND symb_decoder(16#fc#)) OR
 					(reg_q2000 AND symb_decoder(16#87#)) OR
 					(reg_q2000 AND symb_decoder(16#8f#)) OR
 					(reg_q2000 AND symb_decoder(16#78#)) OR
 					(reg_q2000 AND symb_decoder(16#69#)) OR
 					(reg_q2000 AND symb_decoder(16#7b#)) OR
 					(reg_q2000 AND symb_decoder(16#f2#)) OR
 					(reg_q2000 AND symb_decoder(16#ca#)) OR
 					(reg_q2000 AND symb_decoder(16#7e#)) OR
 					(reg_q2000 AND symb_decoder(16#01#)) OR
 					(reg_q2000 AND symb_decoder(16#82#)) OR
 					(reg_q2000 AND symb_decoder(16#ae#)) OR
 					(reg_q2000 AND symb_decoder(16#2d#)) OR
 					(reg_q2000 AND symb_decoder(16#77#)) OR
 					(reg_q2000 AND symb_decoder(16#72#)) OR
 					(reg_q2000 AND symb_decoder(16#e4#)) OR
 					(reg_q2000 AND symb_decoder(16#17#)) OR
 					(reg_q2000 AND symb_decoder(16#3b#)) OR
 					(reg_q2000 AND symb_decoder(16#fe#)) OR
 					(reg_q2000 AND symb_decoder(16#15#)) OR
 					(reg_q2000 AND symb_decoder(16#1c#)) OR
 					(reg_q2000 AND symb_decoder(16#23#)) OR
 					(reg_q2000 AND symb_decoder(16#20#)) OR
 					(reg_q2000 AND symb_decoder(16#11#)) OR
 					(reg_q2000 AND symb_decoder(16#de#)) OR
 					(reg_q2000 AND symb_decoder(16#7f#)) OR
 					(reg_q2000 AND symb_decoder(16#af#)) OR
 					(reg_q2000 AND symb_decoder(16#32#)) OR
 					(reg_q2000 AND symb_decoder(16#b0#)) OR
 					(reg_q2000 AND symb_decoder(16#57#)) OR
 					(reg_q2000 AND symb_decoder(16#7a#)) OR
 					(reg_q2000 AND symb_decoder(16#bb#)) OR
 					(reg_q2000 AND symb_decoder(16#0d#)) OR
 					(reg_q2000 AND symb_decoder(16#95#)) OR
 					(reg_q2000 AND symb_decoder(16#8d#)) OR
 					(reg_q2000 AND symb_decoder(16#48#)) OR
 					(reg_q2000 AND symb_decoder(16#06#)) OR
 					(reg_q2000 AND symb_decoder(16#07#)) OR
 					(reg_q2000 AND symb_decoder(16#2b#)) OR
 					(reg_q2000 AND symb_decoder(16#68#)) OR
 					(reg_q2000 AND symb_decoder(16#34#)) OR
 					(reg_q2000 AND symb_decoder(16#37#)) OR
 					(reg_q2000 AND symb_decoder(16#3c#)) OR
 					(reg_q2000 AND symb_decoder(16#6b#)) OR
 					(reg_q2000 AND symb_decoder(16#36#)) OR
 					(reg_q2000 AND symb_decoder(16#aa#)) OR
 					(reg_q2000 AND symb_decoder(16#66#)) OR
 					(reg_q2000 AND symb_decoder(16#59#)) OR
 					(reg_q2000 AND symb_decoder(16#6e#)) OR
 					(reg_q2000 AND symb_decoder(16#f0#)) OR
 					(reg_q2000 AND symb_decoder(16#ed#)) OR
 					(reg_q2000 AND symb_decoder(16#bf#)) OR
 					(reg_q2000 AND symb_decoder(16#ef#)) OR
 					(reg_q2000 AND symb_decoder(16#71#)) OR
 					(reg_q2000 AND symb_decoder(16#a6#)) OR
 					(reg_q2000 AND symb_decoder(16#a4#)) OR
 					(reg_q2000 AND symb_decoder(16#a2#)) OR
 					(reg_q2000 AND symb_decoder(16#61#)) OR
 					(reg_q2000 AND symb_decoder(16#3f#)) OR
 					(reg_q2000 AND symb_decoder(16#a3#)) OR
 					(reg_q2000 AND symb_decoder(16#ac#)) OR
 					(reg_q2000 AND symb_decoder(16#1f#)) OR
 					(reg_q2000 AND symb_decoder(16#c8#)) OR
 					(reg_q2000 AND symb_decoder(16#55#)) OR
 					(reg_q2000 AND symb_decoder(16#b7#)) OR
 					(reg_q2000 AND symb_decoder(16#46#)) OR
 					(reg_q2000 AND symb_decoder(16#f7#)) OR
 					(reg_q2000 AND symb_decoder(16#fd#)) OR
 					(reg_q2000 AND symb_decoder(16#ba#)) OR
 					(reg_q2000 AND symb_decoder(16#14#)) OR
 					(reg_q2000 AND symb_decoder(16#c4#)) OR
 					(reg_q2000 AND symb_decoder(16#41#)) OR
 					(reg_q2000 AND symb_decoder(16#6a#)) OR
 					(reg_q2000 AND symb_decoder(16#d6#)) OR
 					(reg_q2000 AND symb_decoder(16#00#)) OR
 					(reg_q2000 AND symb_decoder(16#4e#)) OR
 					(reg_q2000 AND symb_decoder(16#d9#)) OR
 					(reg_q2000 AND symb_decoder(16#d3#)) OR
 					(reg_q2000 AND symb_decoder(16#65#)) OR
 					(reg_q2000 AND symb_decoder(16#51#)) OR
 					(reg_q2000 AND symb_decoder(16#88#)) OR
 					(reg_q2000 AND symb_decoder(16#fa#)) OR
 					(reg_q2000 AND symb_decoder(16#c3#)) OR
 					(reg_q2000 AND symb_decoder(16#29#)) OR
 					(reg_q2000 AND symb_decoder(16#3a#)) OR
 					(reg_q2000 AND symb_decoder(16#a8#)) OR
 					(reg_q2000 AND symb_decoder(16#44#)) OR
 					(reg_q2000 AND symb_decoder(16#e5#)) OR
 					(reg_q2000 AND symb_decoder(16#13#)) OR
 					(reg_q2000 AND symb_decoder(16#ab#)) OR
 					(reg_q2000 AND symb_decoder(16#d5#)) OR
 					(reg_q2000 AND symb_decoder(16#33#)) OR
 					(reg_q2000 AND symb_decoder(16#94#)) OR
 					(reg_q2000 AND symb_decoder(16#02#)) OR
 					(reg_q2000 AND symb_decoder(16#40#)) OR
 					(reg_q2000 AND symb_decoder(16#b8#)) OR
 					(reg_q2000 AND symb_decoder(16#db#)) OR
 					(reg_q2000 AND symb_decoder(16#9c#)) OR
 					(reg_q2000 AND symb_decoder(16#75#)) OR
 					(reg_q2000 AND symb_decoder(16#a5#)) OR
 					(reg_q2000 AND symb_decoder(16#e0#)) OR
 					(reg_q2000 AND symb_decoder(16#54#)) OR
 					(reg_q2000 AND symb_decoder(16#f8#)) OR
 					(reg_q2000 AND symb_decoder(16#38#)) OR
 					(reg_q2000 AND symb_decoder(16#be#)) OR
 					(reg_q2000 AND symb_decoder(16#b4#)) OR
 					(reg_q2000 AND symb_decoder(16#c7#)) OR
 					(reg_q2000 AND symb_decoder(16#bd#)) OR
 					(reg_q2000 AND symb_decoder(16#47#)) OR
 					(reg_q2000 AND symb_decoder(16#50#)) OR
 					(reg_q2000 AND symb_decoder(16#18#)) OR
 					(reg_q2000 AND symb_decoder(16#ad#)) OR
 					(reg_q2000 AND symb_decoder(16#9d#)) OR
 					(reg_q2000 AND symb_decoder(16#1b#)) OR
 					(reg_q2000 AND symb_decoder(16#74#)) OR
 					(reg_q2000 AND symb_decoder(16#03#)) OR
 					(reg_q2000 AND symb_decoder(16#96#)) OR
 					(reg_q2000 AND symb_decoder(16#dd#)) OR
 					(reg_q2000 AND symb_decoder(16#1e#)) OR
 					(reg_q2000 AND symb_decoder(16#d0#)) OR
 					(reg_q2000 AND symb_decoder(16#a0#)) OR
 					(reg_q2000 AND symb_decoder(16#99#)) OR
 					(reg_q2000 AND symb_decoder(16#83#)) OR
 					(reg_q2000 AND symb_decoder(16#ea#)) OR
 					(reg_q2000 AND symb_decoder(16#67#)) OR
 					(reg_q2000 AND symb_decoder(16#5a#)) OR
 					(reg_q2000 AND symb_decoder(16#45#)) OR
 					(reg_q2000 AND symb_decoder(16#d1#)) OR
 					(reg_q2000 AND symb_decoder(16#cc#)) OR
 					(reg_q2000 AND symb_decoder(16#8a#)) OR
 					(reg_q2000 AND symb_decoder(16#5d#)) OR
 					(reg_q2000 AND symb_decoder(16#9a#)) OR
 					(reg_q2000 AND symb_decoder(16#da#)) OR
 					(reg_q2000 AND symb_decoder(16#52#)) OR
 					(reg_q2000 AND symb_decoder(16#2a#)) OR
 					(reg_q2000 AND symb_decoder(16#2e#)) OR
 					(reg_q2000 AND symb_decoder(16#91#)) OR
 					(reg_q2000 AND symb_decoder(16#cf#)) OR
 					(reg_q2000 AND symb_decoder(16#0f#)) OR
 					(reg_q2000 AND symb_decoder(16#df#)) OR
 					(reg_q2000 AND symb_decoder(16#43#)) OR
 					(reg_q2000 AND symb_decoder(16#d2#)) OR
 					(reg_q2000 AND symb_decoder(16#12#)) OR
 					(reg_q2000 AND symb_decoder(16#89#)) OR
 					(reg_q2000 AND symb_decoder(16#8e#)) OR
 					(reg_q2000 AND symb_decoder(16#49#)) OR
 					(reg_q2000 AND symb_decoder(16#64#)) OR
 					(reg_q2000 AND symb_decoder(16#4f#)) OR
 					(reg_q2000 AND symb_decoder(16#39#)) OR
 					(reg_q2000 AND symb_decoder(16#08#)) OR
 					(reg_q2000 AND symb_decoder(16#d4#)) OR
 					(reg_q2000 AND symb_decoder(16#73#)) OR
 					(reg_q2000 AND symb_decoder(16#24#)) OR
 					(reg_q2000 AND symb_decoder(16#e3#)) OR
 					(reg_q2000 AND symb_decoder(16#90#)) OR
 					(reg_q2000 AND symb_decoder(16#85#)) OR
 					(reg_q2000 AND symb_decoder(16#5b#)) OR
 					(reg_q2000 AND symb_decoder(16#0c#)) OR
 					(reg_q2000 AND symb_decoder(16#62#)) OR
 					(reg_q2000 AND symb_decoder(16#d8#)) OR
 					(reg_q2000 AND symb_decoder(16#c6#)) OR
 					(reg_q2000 AND symb_decoder(16#2c#)) OR
 					(reg_q2000 AND symb_decoder(16#b1#)) OR
 					(reg_q2000 AND symb_decoder(16#a7#)) OR
 					(reg_q2000 AND symb_decoder(16#6f#)) OR
 					(reg_q2000 AND symb_decoder(16#22#)) OR
 					(reg_q2000 AND symb_decoder(16#cd#)) OR
 					(reg_q2000 AND symb_decoder(16#6d#)) OR
 					(reg_q2000 AND symb_decoder(16#97#)) OR
 					(reg_q2000 AND symb_decoder(16#0a#)) OR
 					(reg_q2000 AND symb_decoder(16#f5#)) OR
 					(reg_q2000 AND symb_decoder(16#92#)) OR
 					(reg_q2000 AND symb_decoder(16#a1#)) OR
 					(reg_q2000 AND symb_decoder(16#bc#)) OR
 					(reg_q2000 AND symb_decoder(16#25#)) OR
 					(reg_q2000 AND symb_decoder(16#04#)) OR
 					(reg_q2000 AND symb_decoder(16#dc#)) OR
 					(reg_q2000 AND symb_decoder(16#7d#)) OR
 					(reg_q2000 AND symb_decoder(16#4c#)) OR
 					(reg_q2000 AND symb_decoder(16#79#)) OR
 					(reg_q2000 AND symb_decoder(16#ee#)) OR
 					(reg_q2000 AND symb_decoder(16#8b#)) OR
 					(reg_q2000 AND symb_decoder(16#10#)) OR
 					(reg_q2000 AND symb_decoder(16#60#)) OR
 					(reg_q2000 AND symb_decoder(16#8c#)) OR
 					(reg_q2000 AND symb_decoder(16#3d#)) OR
 					(reg_q2000 AND symb_decoder(16#b2#)) OR
 					(reg_q2000 AND symb_decoder(16#30#)) OR
 					(reg_q2000 AND symb_decoder(16#81#)) OR
 					(reg_q2000 AND symb_decoder(16#76#)) OR
 					(reg_q2000 AND symb_decoder(16#31#)) OR
 					(reg_q2000 AND symb_decoder(16#c2#)) OR
 					(reg_q2000 AND symb_decoder(16#eb#)) OR
 					(reg_q2000 AND symb_decoder(16#5e#)) OR
 					(reg_q2000 AND symb_decoder(16#42#)) OR
 					(reg_q2000 AND symb_decoder(16#b6#)) OR
 					(reg_q2000 AND symb_decoder(16#28#)) OR
 					(reg_q2000 AND symb_decoder(16#b9#)) OR
 					(reg_q2000 AND symb_decoder(16#f3#)) OR
 					(reg_q2000 AND symb_decoder(16#05#)) OR
 					(reg_q2000 AND symb_decoder(16#80#)) OR
 					(reg_q2000 AND symb_decoder(16#c5#)) OR
 					(reg_q2000 AND symb_decoder(16#86#)) OR
 					(reg_q2000 AND symb_decoder(16#b3#)) OR
 					(reg_q2000 AND symb_decoder(16#16#)) OR
 					(reg_q2000 AND symb_decoder(16#0b#)) OR
 					(reg_q2000 AND symb_decoder(16#3e#)) OR
 					(reg_q2000 AND symb_decoder(16#e9#)) OR
 					(reg_q2000 AND symb_decoder(16#ce#)) OR
 					(reg_q2000 AND symb_decoder(16#4b#)) OR
 					(reg_q2000 AND symb_decoder(16#e1#)) OR
 					(reg_q2000 AND symb_decoder(16#58#)) OR
 					(reg_q2000 AND symb_decoder(16#4d#)) OR
 					(reg_q2000 AND symb_decoder(16#93#)) OR
 					(reg_q2000 AND symb_decoder(16#c9#)) OR
 					(reg_q2000 AND symb_decoder(16#ec#)) OR
 					(reg_q2000 AND symb_decoder(16#fb#)) OR
 					(reg_q2000 AND symb_decoder(16#f9#)) OR
 					(reg_q2000 AND symb_decoder(16#cb#)) OR
 					(reg_q2000 AND symb_decoder(16#1a#)) OR
 					(reg_q2000 AND symb_decoder(16#7c#)) OR
 					(reg_q2000 AND symb_decoder(16#5f#));
reg_q2000_init <= '0' ;
	p_reg_q2000: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2000 <= reg_q2000_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2000 <= reg_q2000_init;
        else
          reg_q2000 <= reg_q2000_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q225_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q225 AND symb_decoder(16#d9#)) OR
 					(reg_q225 AND symb_decoder(16#09#)) OR
 					(reg_q225 AND symb_decoder(16#a9#)) OR
 					(reg_q225 AND symb_decoder(16#74#)) OR
 					(reg_q225 AND symb_decoder(16#15#)) OR
 					(reg_q225 AND symb_decoder(16#a5#)) OR
 					(reg_q225 AND symb_decoder(16#98#)) OR
 					(reg_q225 AND symb_decoder(16#e3#)) OR
 					(reg_q225 AND symb_decoder(16#78#)) OR
 					(reg_q225 AND symb_decoder(16#45#)) OR
 					(reg_q225 AND symb_decoder(16#92#)) OR
 					(reg_q225 AND symb_decoder(16#0a#)) OR
 					(reg_q225 AND symb_decoder(16#e9#)) OR
 					(reg_q225 AND symb_decoder(16#63#)) OR
 					(reg_q225 AND symb_decoder(16#ae#)) OR
 					(reg_q225 AND symb_decoder(16#d5#)) OR
 					(reg_q225 AND symb_decoder(16#f3#)) OR
 					(reg_q225 AND symb_decoder(16#96#)) OR
 					(reg_q225 AND symb_decoder(16#80#)) OR
 					(reg_q225 AND symb_decoder(16#7c#)) OR
 					(reg_q225 AND symb_decoder(16#39#)) OR
 					(reg_q225 AND symb_decoder(16#1d#)) OR
 					(reg_q225 AND symb_decoder(16#8f#)) OR
 					(reg_q225 AND symb_decoder(16#0d#)) OR
 					(reg_q225 AND symb_decoder(16#01#)) OR
 					(reg_q225 AND symb_decoder(16#cc#)) OR
 					(reg_q225 AND symb_decoder(16#d0#)) OR
 					(reg_q225 AND symb_decoder(16#68#)) OR
 					(reg_q225 AND symb_decoder(16#6f#)) OR
 					(reg_q225 AND symb_decoder(16#37#)) OR
 					(reg_q225 AND symb_decoder(16#ba#)) OR
 					(reg_q225 AND symb_decoder(16#1b#)) OR
 					(reg_q225 AND symb_decoder(16#cf#)) OR
 					(reg_q225 AND symb_decoder(16#d3#)) OR
 					(reg_q225 AND symb_decoder(16#12#)) OR
 					(reg_q225 AND symb_decoder(16#a0#)) OR
 					(reg_q225 AND symb_decoder(16#eb#)) OR
 					(reg_q225 AND symb_decoder(16#87#)) OR
 					(reg_q225 AND symb_decoder(16#29#)) OR
 					(reg_q225 AND symb_decoder(16#32#)) OR
 					(reg_q225 AND symb_decoder(16#6e#)) OR
 					(reg_q225 AND symb_decoder(16#3c#)) OR
 					(reg_q225 AND symb_decoder(16#b6#)) OR
 					(reg_q225 AND symb_decoder(16#86#)) OR
 					(reg_q225 AND symb_decoder(16#6c#)) OR
 					(reg_q225 AND symb_decoder(16#b8#)) OR
 					(reg_q225 AND symb_decoder(16#e7#)) OR
 					(reg_q225 AND symb_decoder(16#ca#)) OR
 					(reg_q225 AND symb_decoder(16#02#)) OR
 					(reg_q225 AND symb_decoder(16#51#)) OR
 					(reg_q225 AND symb_decoder(16#17#)) OR
 					(reg_q225 AND symb_decoder(16#2e#)) OR
 					(reg_q225 AND symb_decoder(16#f9#)) OR
 					(reg_q225 AND symb_decoder(16#5e#)) OR
 					(reg_q225 AND symb_decoder(16#76#)) OR
 					(reg_q225 AND symb_decoder(16#25#)) OR
 					(reg_q225 AND symb_decoder(16#30#)) OR
 					(reg_q225 AND symb_decoder(16#21#)) OR
 					(reg_q225 AND symb_decoder(16#55#)) OR
 					(reg_q225 AND symb_decoder(16#c1#)) OR
 					(reg_q225 AND symb_decoder(16#85#)) OR
 					(reg_q225 AND symb_decoder(16#7e#)) OR
 					(reg_q225 AND symb_decoder(16#f7#)) OR
 					(reg_q225 AND symb_decoder(16#82#)) OR
 					(reg_q225 AND symb_decoder(16#af#)) OR
 					(reg_q225 AND symb_decoder(16#7b#)) OR
 					(reg_q225 AND symb_decoder(16#b9#)) OR
 					(reg_q225 AND symb_decoder(16#08#)) OR
 					(reg_q225 AND symb_decoder(16#1c#)) OR
 					(reg_q225 AND symb_decoder(16#84#)) OR
 					(reg_q225 AND symb_decoder(16#3a#)) OR
 					(reg_q225 AND symb_decoder(16#4a#)) OR
 					(reg_q225 AND symb_decoder(16#58#)) OR
 					(reg_q225 AND symb_decoder(16#18#)) OR
 					(reg_q225 AND symb_decoder(16#9a#)) OR
 					(reg_q225 AND symb_decoder(16#8d#)) OR
 					(reg_q225 AND symb_decoder(16#e6#)) OR
 					(reg_q225 AND symb_decoder(16#db#)) OR
 					(reg_q225 AND symb_decoder(16#d4#)) OR
 					(reg_q225 AND symb_decoder(16#4d#)) OR
 					(reg_q225 AND symb_decoder(16#77#)) OR
 					(reg_q225 AND symb_decoder(16#06#)) OR
 					(reg_q225 AND symb_decoder(16#5a#)) OR
 					(reg_q225 AND symb_decoder(16#ec#)) OR
 					(reg_q225 AND symb_decoder(16#b0#)) OR
 					(reg_q225 AND symb_decoder(16#e5#)) OR
 					(reg_q225 AND symb_decoder(16#94#)) OR
 					(reg_q225 AND symb_decoder(16#4f#)) OR
 					(reg_q225 AND symb_decoder(16#cb#)) OR
 					(reg_q225 AND symb_decoder(16#19#)) OR
 					(reg_q225 AND symb_decoder(16#0b#)) OR
 					(reg_q225 AND symb_decoder(16#8b#)) OR
 					(reg_q225 AND symb_decoder(16#b4#)) OR
 					(reg_q225 AND symb_decoder(16#bc#)) OR
 					(reg_q225 AND symb_decoder(16#46#)) OR
 					(reg_q225 AND symb_decoder(16#c4#)) OR
 					(reg_q225 AND symb_decoder(16#05#)) OR
 					(reg_q225 AND symb_decoder(16#5d#)) OR
 					(reg_q225 AND symb_decoder(16#d1#)) OR
 					(reg_q225 AND symb_decoder(16#93#)) OR
 					(reg_q225 AND symb_decoder(16#24#)) OR
 					(reg_q225 AND symb_decoder(16#71#)) OR
 					(reg_q225 AND symb_decoder(16#c8#)) OR
 					(reg_q225 AND symb_decoder(16#95#)) OR
 					(reg_q225 AND symb_decoder(16#c3#)) OR
 					(reg_q225 AND symb_decoder(16#e1#)) OR
 					(reg_q225 AND symb_decoder(16#3d#)) OR
 					(reg_q225 AND symb_decoder(16#28#)) OR
 					(reg_q225 AND symb_decoder(16#d7#)) OR
 					(reg_q225 AND symb_decoder(16#fe#)) OR
 					(reg_q225 AND symb_decoder(16#ce#)) OR
 					(reg_q225 AND symb_decoder(16#2a#)) OR
 					(reg_q225 AND symb_decoder(16#e8#)) OR
 					(reg_q225 AND symb_decoder(16#83#)) OR
 					(reg_q225 AND symb_decoder(16#72#)) OR
 					(reg_q225 AND symb_decoder(16#ff#)) OR
 					(reg_q225 AND symb_decoder(16#f2#)) OR
 					(reg_q225 AND symb_decoder(16#88#)) OR
 					(reg_q225 AND symb_decoder(16#22#)) OR
 					(reg_q225 AND symb_decoder(16#43#)) OR
 					(reg_q225 AND symb_decoder(16#5f#)) OR
 					(reg_q225 AND symb_decoder(16#b7#)) OR
 					(reg_q225 AND symb_decoder(16#bd#)) OR
 					(reg_q225 AND symb_decoder(16#be#)) OR
 					(reg_q225 AND symb_decoder(16#59#)) OR
 					(reg_q225 AND symb_decoder(16#50#)) OR
 					(reg_q225 AND symb_decoder(16#0e#)) OR
 					(reg_q225 AND symb_decoder(16#8c#)) OR
 					(reg_q225 AND symb_decoder(16#60#)) OR
 					(reg_q225 AND symb_decoder(16#d8#)) OR
 					(reg_q225 AND symb_decoder(16#dc#)) OR
 					(reg_q225 AND symb_decoder(16#ef#)) OR
 					(reg_q225 AND symb_decoder(16#8e#)) OR
 					(reg_q225 AND symb_decoder(16#bb#)) OR
 					(reg_q225 AND symb_decoder(16#d2#)) OR
 					(reg_q225 AND symb_decoder(16#b5#)) OR
 					(reg_q225 AND symb_decoder(16#f4#)) OR
 					(reg_q225 AND symb_decoder(16#4c#)) OR
 					(reg_q225 AND symb_decoder(16#97#)) OR
 					(reg_q225 AND symb_decoder(16#27#)) OR
 					(reg_q225 AND symb_decoder(16#2b#)) OR
 					(reg_q225 AND symb_decoder(16#56#)) OR
 					(reg_q225 AND symb_decoder(16#62#)) OR
 					(reg_q225 AND symb_decoder(16#16#)) OR
 					(reg_q225 AND symb_decoder(16#9b#)) OR
 					(reg_q225 AND symb_decoder(16#91#)) OR
 					(reg_q225 AND symb_decoder(16#f0#)) OR
 					(reg_q225 AND symb_decoder(16#7f#)) OR
 					(reg_q225 AND symb_decoder(16#3e#)) OR
 					(reg_q225 AND symb_decoder(16#73#)) OR
 					(reg_q225 AND symb_decoder(16#c0#)) OR
 					(reg_q225 AND symb_decoder(16#81#)) OR
 					(reg_q225 AND symb_decoder(16#75#)) OR
 					(reg_q225 AND symb_decoder(16#a4#)) OR
 					(reg_q225 AND symb_decoder(16#9f#)) OR
 					(reg_q225 AND symb_decoder(16#52#)) OR
 					(reg_q225 AND symb_decoder(16#9e#)) OR
 					(reg_q225 AND symb_decoder(16#31#)) OR
 					(reg_q225 AND symb_decoder(16#41#)) OR
 					(reg_q225 AND symb_decoder(16#2d#)) OR
 					(reg_q225 AND symb_decoder(16#de#)) OR
 					(reg_q225 AND symb_decoder(16#fa#)) OR
 					(reg_q225 AND symb_decoder(16#5c#)) OR
 					(reg_q225 AND symb_decoder(16#5b#)) OR
 					(reg_q225 AND symb_decoder(16#a8#)) OR
 					(reg_q225 AND symb_decoder(16#da#)) OR
 					(reg_q225 AND symb_decoder(16#3b#)) OR
 					(reg_q225 AND symb_decoder(16#36#)) OR
 					(reg_q225 AND symb_decoder(16#89#)) OR
 					(reg_q225 AND symb_decoder(16#6b#)) OR
 					(reg_q225 AND symb_decoder(16#e4#)) OR
 					(reg_q225 AND symb_decoder(16#35#)) OR
 					(reg_q225 AND symb_decoder(16#14#)) OR
 					(reg_q225 AND symb_decoder(16#79#)) OR
 					(reg_q225 AND symb_decoder(16#48#)) OR
 					(reg_q225 AND symb_decoder(16#e2#)) OR
 					(reg_q225 AND symb_decoder(16#04#)) OR
 					(reg_q225 AND symb_decoder(16#c2#)) OR
 					(reg_q225 AND symb_decoder(16#a1#)) OR
 					(reg_q225 AND symb_decoder(16#90#)) OR
 					(reg_q225 AND symb_decoder(16#a7#)) OR
 					(reg_q225 AND symb_decoder(16#38#)) OR
 					(reg_q225 AND symb_decoder(16#99#)) OR
 					(reg_q225 AND symb_decoder(16#b3#)) OR
 					(reg_q225 AND symb_decoder(16#fc#)) OR
 					(reg_q225 AND symb_decoder(16#9d#)) OR
 					(reg_q225 AND symb_decoder(16#e0#)) OR
 					(reg_q225 AND symb_decoder(16#53#)) OR
 					(reg_q225 AND symb_decoder(16#70#)) OR
 					(reg_q225 AND symb_decoder(16#fb#)) OR
 					(reg_q225 AND symb_decoder(16#11#)) OR
 					(reg_q225 AND symb_decoder(16#a2#)) OR
 					(reg_q225 AND symb_decoder(16#00#)) OR
 					(reg_q225 AND symb_decoder(16#0c#)) OR
 					(reg_q225 AND symb_decoder(16#f1#)) OR
 					(reg_q225 AND symb_decoder(16#23#)) OR
 					(reg_q225 AND symb_decoder(16#c5#)) OR
 					(reg_q225 AND symb_decoder(16#ab#)) OR
 					(reg_q225 AND symb_decoder(16#2f#)) OR
 					(reg_q225 AND symb_decoder(16#f5#)) OR
 					(reg_q225 AND symb_decoder(16#dd#)) OR
 					(reg_q225 AND symb_decoder(16#8a#)) OR
 					(reg_q225 AND symb_decoder(16#4e#)) OR
 					(reg_q225 AND symb_decoder(16#ad#)) OR
 					(reg_q225 AND symb_decoder(16#9c#)) OR
 					(reg_q225 AND symb_decoder(16#10#)) OR
 					(reg_q225 AND symb_decoder(16#cd#)) OR
 					(reg_q225 AND symb_decoder(16#49#)) OR
 					(reg_q225 AND symb_decoder(16#b2#)) OR
 					(reg_q225 AND symb_decoder(16#b1#)) OR
 					(reg_q225 AND symb_decoder(16#69#)) OR
 					(reg_q225 AND symb_decoder(16#3f#)) OR
 					(reg_q225 AND symb_decoder(16#1f#)) OR
 					(reg_q225 AND symb_decoder(16#57#)) OR
 					(reg_q225 AND symb_decoder(16#ac#)) OR
 					(reg_q225 AND symb_decoder(16#6a#)) OR
 					(reg_q225 AND symb_decoder(16#26#)) OR
 					(reg_q225 AND symb_decoder(16#44#)) OR
 					(reg_q225 AND symb_decoder(16#34#)) OR
 					(reg_q225 AND symb_decoder(16#67#)) OR
 					(reg_q225 AND symb_decoder(16#64#)) OR
 					(reg_q225 AND symb_decoder(16#1e#)) OR
 					(reg_q225 AND symb_decoder(16#13#)) OR
 					(reg_q225 AND symb_decoder(16#c9#)) OR
 					(reg_q225 AND symb_decoder(16#4b#)) OR
 					(reg_q225 AND symb_decoder(16#2c#)) OR
 					(reg_q225 AND symb_decoder(16#df#)) OR
 					(reg_q225 AND symb_decoder(16#c6#)) OR
 					(reg_q225 AND symb_decoder(16#a6#)) OR
 					(reg_q225 AND symb_decoder(16#33#)) OR
 					(reg_q225 AND symb_decoder(16#f8#)) OR
 					(reg_q225 AND symb_decoder(16#66#)) OR
 					(reg_q225 AND symb_decoder(16#c7#)) OR
 					(reg_q225 AND symb_decoder(16#fd#)) OR
 					(reg_q225 AND symb_decoder(16#07#)) OR
 					(reg_q225 AND symb_decoder(16#aa#)) OR
 					(reg_q225 AND symb_decoder(16#20#)) OR
 					(reg_q225 AND symb_decoder(16#42#)) OR
 					(reg_q225 AND symb_decoder(16#ea#)) OR
 					(reg_q225 AND symb_decoder(16#7d#)) OR
 					(reg_q225 AND symb_decoder(16#a3#)) OR
 					(reg_q225 AND symb_decoder(16#0f#)) OR
 					(reg_q225 AND symb_decoder(16#47#)) OR
 					(reg_q225 AND symb_decoder(16#f6#)) OR
 					(reg_q225 AND symb_decoder(16#1a#)) OR
 					(reg_q225 AND symb_decoder(16#40#)) OR
 					(reg_q225 AND symb_decoder(16#ed#)) OR
 					(reg_q225 AND symb_decoder(16#bf#)) OR
 					(reg_q225 AND symb_decoder(16#d6#)) OR
 					(reg_q225 AND symb_decoder(16#61#)) OR
 					(reg_q225 AND symb_decoder(16#65#)) OR
 					(reg_q225 AND symb_decoder(16#03#)) OR
 					(reg_q225 AND symb_decoder(16#6d#)) OR
 					(reg_q225 AND symb_decoder(16#7a#)) OR
 					(reg_q225 AND symb_decoder(16#54#)) OR
 					(reg_q225 AND symb_decoder(16#ee#));
reg_q225_init <= '0' ;
	p_reg_q225: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q225 <= reg_q225_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q225 <= reg_q225_init;
        else
          reg_q225 <= reg_q225_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q899_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q899 AND symb_decoder(16#5d#)) OR
 					(reg_q899 AND symb_decoder(16#fd#)) OR
 					(reg_q899 AND symb_decoder(16#94#)) OR
 					(reg_q899 AND symb_decoder(16#7b#)) OR
 					(reg_q899 AND symb_decoder(16#b8#)) OR
 					(reg_q899 AND symb_decoder(16#2b#)) OR
 					(reg_q899 AND symb_decoder(16#1e#)) OR
 					(reg_q899 AND symb_decoder(16#7d#)) OR
 					(reg_q899 AND symb_decoder(16#e9#)) OR
 					(reg_q899 AND symb_decoder(16#4e#)) OR
 					(reg_q899 AND symb_decoder(16#48#)) OR
 					(reg_q899 AND symb_decoder(16#d0#)) OR
 					(reg_q899 AND symb_decoder(16#6c#)) OR
 					(reg_q899 AND symb_decoder(16#21#)) OR
 					(reg_q899 AND symb_decoder(16#59#)) OR
 					(reg_q899 AND symb_decoder(16#82#)) OR
 					(reg_q899 AND symb_decoder(16#5b#)) OR
 					(reg_q899 AND symb_decoder(16#99#)) OR
 					(reg_q899 AND symb_decoder(16#02#)) OR
 					(reg_q899 AND symb_decoder(16#74#)) OR
 					(reg_q899 AND symb_decoder(16#52#)) OR
 					(reg_q899 AND symb_decoder(16#bf#)) OR
 					(reg_q899 AND symb_decoder(16#35#)) OR
 					(reg_q899 AND symb_decoder(16#67#)) OR
 					(reg_q899 AND symb_decoder(16#51#)) OR
 					(reg_q899 AND symb_decoder(16#aa#)) OR
 					(reg_q899 AND symb_decoder(16#55#)) OR
 					(reg_q899 AND symb_decoder(16#62#)) OR
 					(reg_q899 AND symb_decoder(16#da#)) OR
 					(reg_q899 AND symb_decoder(16#4b#)) OR
 					(reg_q899 AND symb_decoder(16#12#)) OR
 					(reg_q899 AND symb_decoder(16#ac#)) OR
 					(reg_q899 AND symb_decoder(16#25#)) OR
 					(reg_q899 AND symb_decoder(16#38#)) OR
 					(reg_q899 AND symb_decoder(16#b0#)) OR
 					(reg_q899 AND symb_decoder(16#a9#)) OR
 					(reg_q899 AND symb_decoder(16#bb#)) OR
 					(reg_q899 AND symb_decoder(16#68#)) OR
 					(reg_q899 AND symb_decoder(16#60#)) OR
 					(reg_q899 AND symb_decoder(16#72#)) OR
 					(reg_q899 AND symb_decoder(16#b7#)) OR
 					(reg_q899 AND symb_decoder(16#c7#)) OR
 					(reg_q899 AND symb_decoder(16#c3#)) OR
 					(reg_q899 AND symb_decoder(16#a2#)) OR
 					(reg_q899 AND symb_decoder(16#71#)) OR
 					(reg_q899 AND symb_decoder(16#4f#)) OR
 					(reg_q899 AND symb_decoder(16#1c#)) OR
 					(reg_q899 AND symb_decoder(16#0c#)) OR
 					(reg_q899 AND symb_decoder(16#f9#)) OR
 					(reg_q899 AND symb_decoder(16#30#)) OR
 					(reg_q899 AND symb_decoder(16#07#)) OR
 					(reg_q899 AND symb_decoder(16#c9#)) OR
 					(reg_q899 AND symb_decoder(16#af#)) OR
 					(reg_q899 AND symb_decoder(16#e8#)) OR
 					(reg_q899 AND symb_decoder(16#6a#)) OR
 					(reg_q899 AND symb_decoder(16#ff#)) OR
 					(reg_q899 AND symb_decoder(16#2c#)) OR
 					(reg_q899 AND symb_decoder(16#6e#)) OR
 					(reg_q899 AND symb_decoder(16#3d#)) OR
 					(reg_q899 AND symb_decoder(16#d2#)) OR
 					(reg_q899 AND symb_decoder(16#93#)) OR
 					(reg_q899 AND symb_decoder(16#9a#)) OR
 					(reg_q899 AND symb_decoder(16#5c#)) OR
 					(reg_q899 AND symb_decoder(16#d7#)) OR
 					(reg_q899 AND symb_decoder(16#e6#)) OR
 					(reg_q899 AND symb_decoder(16#96#)) OR
 					(reg_q899 AND symb_decoder(16#c2#)) OR
 					(reg_q899 AND symb_decoder(16#c1#)) OR
 					(reg_q899 AND symb_decoder(16#ab#)) OR
 					(reg_q899 AND symb_decoder(16#73#)) OR
 					(reg_q899 AND symb_decoder(16#19#)) OR
 					(reg_q899 AND symb_decoder(16#56#)) OR
 					(reg_q899 AND symb_decoder(16#40#)) OR
 					(reg_q899 AND symb_decoder(16#01#)) OR
 					(reg_q899 AND symb_decoder(16#ef#)) OR
 					(reg_q899 AND symb_decoder(16#43#)) OR
 					(reg_q899 AND symb_decoder(16#b3#)) OR
 					(reg_q899 AND symb_decoder(16#2e#)) OR
 					(reg_q899 AND symb_decoder(16#fe#)) OR
 					(reg_q899 AND symb_decoder(16#cc#)) OR
 					(reg_q899 AND symb_decoder(16#f6#)) OR
 					(reg_q899 AND symb_decoder(16#8c#)) OR
 					(reg_q899 AND symb_decoder(16#29#)) OR
 					(reg_q899 AND symb_decoder(16#57#)) OR
 					(reg_q899 AND symb_decoder(16#76#)) OR
 					(reg_q899 AND symb_decoder(16#13#)) OR
 					(reg_q899 AND symb_decoder(16#eb#)) OR
 					(reg_q899 AND symb_decoder(16#c5#)) OR
 					(reg_q899 AND symb_decoder(16#7e#)) OR
 					(reg_q899 AND symb_decoder(16#9c#)) OR
 					(reg_q899 AND symb_decoder(16#34#)) OR
 					(reg_q899 AND symb_decoder(16#86#)) OR
 					(reg_q899 AND symb_decoder(16#1f#)) OR
 					(reg_q899 AND symb_decoder(16#5e#)) OR
 					(reg_q899 AND symb_decoder(16#e5#)) OR
 					(reg_q899 AND symb_decoder(16#70#)) OR
 					(reg_q899 AND symb_decoder(16#ba#)) OR
 					(reg_q899 AND symb_decoder(16#8e#)) OR
 					(reg_q899 AND symb_decoder(16#49#)) OR
 					(reg_q899 AND symb_decoder(16#79#)) OR
 					(reg_q899 AND symb_decoder(16#d5#)) OR
 					(reg_q899 AND symb_decoder(16#00#)) OR
 					(reg_q899 AND symb_decoder(16#d3#)) OR
 					(reg_q899 AND symb_decoder(16#cd#)) OR
 					(reg_q899 AND symb_decoder(16#cb#)) OR
 					(reg_q899 AND symb_decoder(16#65#)) OR
 					(reg_q899 AND symb_decoder(16#a1#)) OR
 					(reg_q899 AND symb_decoder(16#4d#)) OR
 					(reg_q899 AND symb_decoder(16#d1#)) OR
 					(reg_q899 AND symb_decoder(16#e4#)) OR
 					(reg_q899 AND symb_decoder(16#28#)) OR
 					(reg_q899 AND symb_decoder(16#91#)) OR
 					(reg_q899 AND symb_decoder(16#41#)) OR
 					(reg_q899 AND symb_decoder(16#9f#)) OR
 					(reg_q899 AND symb_decoder(16#ea#)) OR
 					(reg_q899 AND symb_decoder(16#3e#)) OR
 					(reg_q899 AND symb_decoder(16#fb#)) OR
 					(reg_q899 AND symb_decoder(16#e2#)) OR
 					(reg_q899 AND symb_decoder(16#6b#)) OR
 					(reg_q899 AND symb_decoder(16#08#)) OR
 					(reg_q899 AND symb_decoder(16#78#)) OR
 					(reg_q899 AND symb_decoder(16#7a#)) OR
 					(reg_q899 AND symb_decoder(16#85#)) OR
 					(reg_q899 AND symb_decoder(16#5f#)) OR
 					(reg_q899 AND symb_decoder(16#a0#)) OR
 					(reg_q899 AND symb_decoder(16#8f#)) OR
 					(reg_q899 AND symb_decoder(16#a3#)) OR
 					(reg_q899 AND symb_decoder(16#f4#)) OR
 					(reg_q899 AND symb_decoder(16#b9#)) OR
 					(reg_q899 AND symb_decoder(16#0a#)) OR
 					(reg_q899 AND symb_decoder(16#10#)) OR
 					(reg_q899 AND symb_decoder(16#63#)) OR
 					(reg_q899 AND symb_decoder(16#7c#)) OR
 					(reg_q899 AND symb_decoder(16#11#)) OR
 					(reg_q899 AND symb_decoder(16#f7#)) OR
 					(reg_q899 AND symb_decoder(16#84#)) OR
 					(reg_q899 AND symb_decoder(16#6d#)) OR
 					(reg_q899 AND symb_decoder(16#33#)) OR
 					(reg_q899 AND symb_decoder(16#89#)) OR
 					(reg_q899 AND symb_decoder(16#a4#)) OR
 					(reg_q899 AND symb_decoder(16#61#)) OR
 					(reg_q899 AND symb_decoder(16#9e#)) OR
 					(reg_q899 AND symb_decoder(16#98#)) OR
 					(reg_q899 AND symb_decoder(16#37#)) OR
 					(reg_q899 AND symb_decoder(16#0d#)) OR
 					(reg_q899 AND symb_decoder(16#69#)) OR
 					(reg_q899 AND symb_decoder(16#83#)) OR
 					(reg_q899 AND symb_decoder(16#9d#)) OR
 					(reg_q899 AND symb_decoder(16#7f#)) OR
 					(reg_q899 AND symb_decoder(16#58#)) OR
 					(reg_q899 AND symb_decoder(16#36#)) OR
 					(reg_q899 AND symb_decoder(16#1a#)) OR
 					(reg_q899 AND symb_decoder(16#bc#)) OR
 					(reg_q899 AND symb_decoder(16#dc#)) OR
 					(reg_q899 AND symb_decoder(16#ce#)) OR
 					(reg_q899 AND symb_decoder(16#1d#)) OR
 					(reg_q899 AND symb_decoder(16#0f#)) OR
 					(reg_q899 AND symb_decoder(16#80#)) OR
 					(reg_q899 AND symb_decoder(16#23#)) OR
 					(reg_q899 AND symb_decoder(16#ec#)) OR
 					(reg_q899 AND symb_decoder(16#18#)) OR
 					(reg_q899 AND symb_decoder(16#54#)) OR
 					(reg_q899 AND symb_decoder(16#c8#)) OR
 					(reg_q899 AND symb_decoder(16#3f#)) OR
 					(reg_q899 AND symb_decoder(16#c6#)) OR
 					(reg_q899 AND symb_decoder(16#42#)) OR
 					(reg_q899 AND symb_decoder(16#d4#)) OR
 					(reg_q899 AND symb_decoder(16#87#)) OR
 					(reg_q899 AND symb_decoder(16#a8#)) OR
 					(reg_q899 AND symb_decoder(16#15#)) OR
 					(reg_q899 AND symb_decoder(16#e1#)) OR
 					(reg_q899 AND symb_decoder(16#e3#)) OR
 					(reg_q899 AND symb_decoder(16#d9#)) OR
 					(reg_q899 AND symb_decoder(16#17#)) OR
 					(reg_q899 AND symb_decoder(16#14#)) OR
 					(reg_q899 AND symb_decoder(16#f0#)) OR
 					(reg_q899 AND symb_decoder(16#4c#)) OR
 					(reg_q899 AND symb_decoder(16#81#)) OR
 					(reg_q899 AND symb_decoder(16#2d#)) OR
 					(reg_q899 AND symb_decoder(16#df#)) OR
 					(reg_q899 AND symb_decoder(16#de#)) OR
 					(reg_q899 AND symb_decoder(16#fc#)) OR
 					(reg_q899 AND symb_decoder(16#db#)) OR
 					(reg_q899 AND symb_decoder(16#0e#)) OR
 					(reg_q899 AND symb_decoder(16#f8#)) OR
 					(reg_q899 AND symb_decoder(16#39#)) OR
 					(reg_q899 AND symb_decoder(16#fa#)) OR
 					(reg_q899 AND symb_decoder(16#31#)) OR
 					(reg_q899 AND symb_decoder(16#3a#)) OR
 					(reg_q899 AND symb_decoder(16#dd#)) OR
 					(reg_q899 AND symb_decoder(16#44#)) OR
 					(reg_q899 AND symb_decoder(16#6f#)) OR
 					(reg_q899 AND symb_decoder(16#05#)) OR
 					(reg_q899 AND symb_decoder(16#03#)) OR
 					(reg_q899 AND symb_decoder(16#88#)) OR
 					(reg_q899 AND symb_decoder(16#a6#)) OR
 					(reg_q899 AND symb_decoder(16#c4#)) OR
 					(reg_q899 AND symb_decoder(16#46#)) OR
 					(reg_q899 AND symb_decoder(16#20#)) OR
 					(reg_q899 AND symb_decoder(16#8a#)) OR
 					(reg_q899 AND symb_decoder(16#90#)) OR
 					(reg_q899 AND symb_decoder(16#be#)) OR
 					(reg_q899 AND symb_decoder(16#77#)) OR
 					(reg_q899 AND symb_decoder(16#3c#)) OR
 					(reg_q899 AND symb_decoder(16#9b#)) OR
 					(reg_q899 AND symb_decoder(16#64#)) OR
 					(reg_q899 AND symb_decoder(16#95#)) OR
 					(reg_q899 AND symb_decoder(16#ae#)) OR
 					(reg_q899 AND symb_decoder(16#04#)) OR
 					(reg_q899 AND symb_decoder(16#0b#)) OR
 					(reg_q899 AND symb_decoder(16#06#)) OR
 					(reg_q899 AND symb_decoder(16#4a#)) OR
 					(reg_q899 AND symb_decoder(16#ee#)) OR
 					(reg_q899 AND symb_decoder(16#ad#)) OR
 					(reg_q899 AND symb_decoder(16#a5#)) OR
 					(reg_q899 AND symb_decoder(16#3b#)) OR
 					(reg_q899 AND symb_decoder(16#ca#)) OR
 					(reg_q899 AND symb_decoder(16#d6#)) OR
 					(reg_q899 AND symb_decoder(16#2f#)) OR
 					(reg_q899 AND symb_decoder(16#50#)) OR
 					(reg_q899 AND symb_decoder(16#22#)) OR
 					(reg_q899 AND symb_decoder(16#e7#)) OR
 					(reg_q899 AND symb_decoder(16#97#)) OR
 					(reg_q899 AND symb_decoder(16#92#)) OR
 					(reg_q899 AND symb_decoder(16#f1#)) OR
 					(reg_q899 AND symb_decoder(16#75#)) OR
 					(reg_q899 AND symb_decoder(16#cf#)) OR
 					(reg_q899 AND symb_decoder(16#26#)) OR
 					(reg_q899 AND symb_decoder(16#b5#)) OR
 					(reg_q899 AND symb_decoder(16#b2#)) OR
 					(reg_q899 AND symb_decoder(16#8b#)) OR
 					(reg_q899 AND symb_decoder(16#24#)) OR
 					(reg_q899 AND symb_decoder(16#8d#)) OR
 					(reg_q899 AND symb_decoder(16#f2#)) OR
 					(reg_q899 AND symb_decoder(16#b4#)) OR
 					(reg_q899 AND symb_decoder(16#47#)) OR
 					(reg_q899 AND symb_decoder(16#a7#)) OR
 					(reg_q899 AND symb_decoder(16#b6#)) OR
 					(reg_q899 AND symb_decoder(16#16#)) OR
 					(reg_q899 AND symb_decoder(16#1b#)) OR
 					(reg_q899 AND symb_decoder(16#27#)) OR
 					(reg_q899 AND symb_decoder(16#c0#)) OR
 					(reg_q899 AND symb_decoder(16#53#)) OR
 					(reg_q899 AND symb_decoder(16#b1#)) OR
 					(reg_q899 AND symb_decoder(16#2a#)) OR
 					(reg_q899 AND symb_decoder(16#ed#)) OR
 					(reg_q899 AND symb_decoder(16#5a#)) OR
 					(reg_q899 AND symb_decoder(16#f3#)) OR
 					(reg_q899 AND symb_decoder(16#66#)) OR
 					(reg_q899 AND symb_decoder(16#e0#)) OR
 					(reg_q899 AND symb_decoder(16#bd#)) OR
 					(reg_q899 AND symb_decoder(16#32#)) OR
 					(reg_q899 AND symb_decoder(16#f5#)) OR
 					(reg_q899 AND symb_decoder(16#09#)) OR
 					(reg_q899 AND symb_decoder(16#d8#)) OR
 					(reg_q899 AND symb_decoder(16#45#));
reg_q899_init <= '0' ;
	p_reg_q899: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q899 <= reg_q899_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q899 <= reg_q899_init;
        else
          reg_q899 <= reg_q899_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1826_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1826 AND symb_decoder(16#5a#)) OR
 					(reg_q1826 AND symb_decoder(16#dd#)) OR
 					(reg_q1826 AND symb_decoder(16#73#)) OR
 					(reg_q1826 AND symb_decoder(16#07#)) OR
 					(reg_q1826 AND symb_decoder(16#11#)) OR
 					(reg_q1826 AND symb_decoder(16#49#)) OR
 					(reg_q1826 AND symb_decoder(16#bd#)) OR
 					(reg_q1826 AND symb_decoder(16#91#)) OR
 					(reg_q1826 AND symb_decoder(16#c2#)) OR
 					(reg_q1826 AND symb_decoder(16#d3#)) OR
 					(reg_q1826 AND symb_decoder(16#88#)) OR
 					(reg_q1826 AND symb_decoder(16#f7#)) OR
 					(reg_q1826 AND symb_decoder(16#16#)) OR
 					(reg_q1826 AND symb_decoder(16#1f#)) OR
 					(reg_q1826 AND symb_decoder(16#b8#)) OR
 					(reg_q1826 AND symb_decoder(16#cc#)) OR
 					(reg_q1826 AND symb_decoder(16#e7#)) OR
 					(reg_q1826 AND symb_decoder(16#6a#)) OR
 					(reg_q1826 AND symb_decoder(16#75#)) OR
 					(reg_q1826 AND symb_decoder(16#25#)) OR
 					(reg_q1826 AND symb_decoder(16#56#)) OR
 					(reg_q1826 AND symb_decoder(16#12#)) OR
 					(reg_q1826 AND symb_decoder(16#79#)) OR
 					(reg_q1826 AND symb_decoder(16#52#)) OR
 					(reg_q1826 AND symb_decoder(16#2a#)) OR
 					(reg_q1826 AND symb_decoder(16#fb#)) OR
 					(reg_q1826 AND symb_decoder(16#3f#)) OR
 					(reg_q1826 AND symb_decoder(16#37#)) OR
 					(reg_q1826 AND symb_decoder(16#d6#)) OR
 					(reg_q1826 AND symb_decoder(16#6b#)) OR
 					(reg_q1826 AND symb_decoder(16#13#)) OR
 					(reg_q1826 AND symb_decoder(16#df#)) OR
 					(reg_q1826 AND symb_decoder(16#fe#)) OR
 					(reg_q1826 AND symb_decoder(16#9d#)) OR
 					(reg_q1826 AND symb_decoder(16#4e#)) OR
 					(reg_q1826 AND symb_decoder(16#89#)) OR
 					(reg_q1826 AND symb_decoder(16#33#)) OR
 					(reg_q1826 AND symb_decoder(16#99#)) OR
 					(reg_q1826 AND symb_decoder(16#e3#)) OR
 					(reg_q1826 AND symb_decoder(16#7c#)) OR
 					(reg_q1826 AND symb_decoder(16#30#)) OR
 					(reg_q1826 AND symb_decoder(16#35#)) OR
 					(reg_q1826 AND symb_decoder(16#17#)) OR
 					(reg_q1826 AND symb_decoder(16#db#)) OR
 					(reg_q1826 AND symb_decoder(16#ce#)) OR
 					(reg_q1826 AND symb_decoder(16#96#)) OR
 					(reg_q1826 AND symb_decoder(16#c8#)) OR
 					(reg_q1826 AND symb_decoder(16#45#)) OR
 					(reg_q1826 AND symb_decoder(16#ac#)) OR
 					(reg_q1826 AND symb_decoder(16#e4#)) OR
 					(reg_q1826 AND symb_decoder(16#de#)) OR
 					(reg_q1826 AND symb_decoder(16#cd#)) OR
 					(reg_q1826 AND symb_decoder(16#90#)) OR
 					(reg_q1826 AND symb_decoder(16#60#)) OR
 					(reg_q1826 AND symb_decoder(16#b5#)) OR
 					(reg_q1826 AND symb_decoder(16#53#)) OR
 					(reg_q1826 AND symb_decoder(16#8a#)) OR
 					(reg_q1826 AND symb_decoder(16#3d#)) OR
 					(reg_q1826 AND symb_decoder(16#f4#)) OR
 					(reg_q1826 AND symb_decoder(16#c7#)) OR
 					(reg_q1826 AND symb_decoder(16#c5#)) OR
 					(reg_q1826 AND symb_decoder(16#85#)) OR
 					(reg_q1826 AND symb_decoder(16#dc#)) OR
 					(reg_q1826 AND symb_decoder(16#94#)) OR
 					(reg_q1826 AND symb_decoder(16#a3#)) OR
 					(reg_q1826 AND symb_decoder(16#7e#)) OR
 					(reg_q1826 AND symb_decoder(16#40#)) OR
 					(reg_q1826 AND symb_decoder(16#ea#)) OR
 					(reg_q1826 AND symb_decoder(16#f1#)) OR
 					(reg_q1826 AND symb_decoder(16#4a#)) OR
 					(reg_q1826 AND symb_decoder(16#86#)) OR
 					(reg_q1826 AND symb_decoder(16#29#)) OR
 					(reg_q1826 AND symb_decoder(16#39#)) OR
 					(reg_q1826 AND symb_decoder(16#70#)) OR
 					(reg_q1826 AND symb_decoder(16#fd#)) OR
 					(reg_q1826 AND symb_decoder(16#0a#)) OR
 					(reg_q1826 AND symb_decoder(16#ca#)) OR
 					(reg_q1826 AND symb_decoder(16#d2#)) OR
 					(reg_q1826 AND symb_decoder(16#b7#)) OR
 					(reg_q1826 AND symb_decoder(16#a2#)) OR
 					(reg_q1826 AND symb_decoder(16#be#)) OR
 					(reg_q1826 AND symb_decoder(16#15#)) OR
 					(reg_q1826 AND symb_decoder(16#22#)) OR
 					(reg_q1826 AND symb_decoder(16#05#)) OR
 					(reg_q1826 AND symb_decoder(16#4b#)) OR
 					(reg_q1826 AND symb_decoder(16#c9#)) OR
 					(reg_q1826 AND symb_decoder(16#27#)) OR
 					(reg_q1826 AND symb_decoder(16#da#)) OR
 					(reg_q1826 AND symb_decoder(16#b0#)) OR
 					(reg_q1826 AND symb_decoder(16#9f#)) OR
 					(reg_q1826 AND symb_decoder(16#2e#)) OR
 					(reg_q1826 AND symb_decoder(16#69#)) OR
 					(reg_q1826 AND symb_decoder(16#f0#)) OR
 					(reg_q1826 AND symb_decoder(16#8e#)) OR
 					(reg_q1826 AND symb_decoder(16#a1#)) OR
 					(reg_q1826 AND symb_decoder(16#51#)) OR
 					(reg_q1826 AND symb_decoder(16#ed#)) OR
 					(reg_q1826 AND symb_decoder(16#50#)) OR
 					(reg_q1826 AND symb_decoder(16#fa#)) OR
 					(reg_q1826 AND symb_decoder(16#98#)) OR
 					(reg_q1826 AND symb_decoder(16#b2#)) OR
 					(reg_q1826 AND symb_decoder(16#18#)) OR
 					(reg_q1826 AND symb_decoder(16#e2#)) OR
 					(reg_q1826 AND symb_decoder(16#2d#)) OR
 					(reg_q1826 AND symb_decoder(16#78#)) OR
 					(reg_q1826 AND symb_decoder(16#f6#)) OR
 					(reg_q1826 AND symb_decoder(16#a7#)) OR
 					(reg_q1826 AND symb_decoder(16#8c#)) OR
 					(reg_q1826 AND symb_decoder(16#9a#)) OR
 					(reg_q1826 AND symb_decoder(16#0c#)) OR
 					(reg_q1826 AND symb_decoder(16#26#)) OR
 					(reg_q1826 AND symb_decoder(16#ab#)) OR
 					(reg_q1826 AND symb_decoder(16#f9#)) OR
 					(reg_q1826 AND symb_decoder(16#a4#)) OR
 					(reg_q1826 AND symb_decoder(16#03#)) OR
 					(reg_q1826 AND symb_decoder(16#84#)) OR
 					(reg_q1826 AND symb_decoder(16#4c#)) OR
 					(reg_q1826 AND symb_decoder(16#0b#)) OR
 					(reg_q1826 AND symb_decoder(16#f5#)) OR
 					(reg_q1826 AND symb_decoder(16#06#)) OR
 					(reg_q1826 AND symb_decoder(16#5b#)) OR
 					(reg_q1826 AND symb_decoder(16#b4#)) OR
 					(reg_q1826 AND symb_decoder(16#77#)) OR
 					(reg_q1826 AND symb_decoder(16#d9#)) OR
 					(reg_q1826 AND symb_decoder(16#10#)) OR
 					(reg_q1826 AND symb_decoder(16#ef#)) OR
 					(reg_q1826 AND symb_decoder(16#d7#)) OR
 					(reg_q1826 AND symb_decoder(16#58#)) OR
 					(reg_q1826 AND symb_decoder(16#0f#)) OR
 					(reg_q1826 AND symb_decoder(16#eb#)) OR
 					(reg_q1826 AND symb_decoder(16#2f#)) OR
 					(reg_q1826 AND symb_decoder(16#72#)) OR
 					(reg_q1826 AND symb_decoder(16#6c#)) OR
 					(reg_q1826 AND symb_decoder(16#f3#)) OR
 					(reg_q1826 AND symb_decoder(16#8b#)) OR
 					(reg_q1826 AND symb_decoder(16#0e#)) OR
 					(reg_q1826 AND symb_decoder(16#ba#)) OR
 					(reg_q1826 AND symb_decoder(16#92#)) OR
 					(reg_q1826 AND symb_decoder(16#43#)) OR
 					(reg_q1826 AND symb_decoder(16#bf#)) OR
 					(reg_q1826 AND symb_decoder(16#36#)) OR
 					(reg_q1826 AND symb_decoder(16#55#)) OR
 					(reg_q1826 AND symb_decoder(16#8d#)) OR
 					(reg_q1826 AND symb_decoder(16#21#)) OR
 					(reg_q1826 AND symb_decoder(16#04#)) OR
 					(reg_q1826 AND symb_decoder(16#af#)) OR
 					(reg_q1826 AND symb_decoder(16#46#)) OR
 					(reg_q1826 AND symb_decoder(16#c0#)) OR
 					(reg_q1826 AND symb_decoder(16#41#)) OR
 					(reg_q1826 AND symb_decoder(16#e8#)) OR
 					(reg_q1826 AND symb_decoder(16#42#)) OR
 					(reg_q1826 AND symb_decoder(16#f8#)) OR
 					(reg_q1826 AND symb_decoder(16#a8#)) OR
 					(reg_q1826 AND symb_decoder(16#14#)) OR
 					(reg_q1826 AND symb_decoder(16#ad#)) OR
 					(reg_q1826 AND symb_decoder(16#66#)) OR
 					(reg_q1826 AND symb_decoder(16#bb#)) OR
 					(reg_q1826 AND symb_decoder(16#83#)) OR
 					(reg_q1826 AND symb_decoder(16#68#)) OR
 					(reg_q1826 AND symb_decoder(16#ae#)) OR
 					(reg_q1826 AND symb_decoder(16#28#)) OR
 					(reg_q1826 AND symb_decoder(16#bc#)) OR
 					(reg_q1826 AND symb_decoder(16#00#)) OR
 					(reg_q1826 AND symb_decoder(16#4d#)) OR
 					(reg_q1826 AND symb_decoder(16#34#)) OR
 					(reg_q1826 AND symb_decoder(16#e5#)) OR
 					(reg_q1826 AND symb_decoder(16#74#)) OR
 					(reg_q1826 AND symb_decoder(16#57#)) OR
 					(reg_q1826 AND symb_decoder(16#7d#)) OR
 					(reg_q1826 AND symb_decoder(16#4f#)) OR
 					(reg_q1826 AND symb_decoder(16#1e#)) OR
 					(reg_q1826 AND symb_decoder(16#1d#)) OR
 					(reg_q1826 AND symb_decoder(16#6f#)) OR
 					(reg_q1826 AND symb_decoder(16#a0#)) OR
 					(reg_q1826 AND symb_decoder(16#09#)) OR
 					(reg_q1826 AND symb_decoder(16#61#)) OR
 					(reg_q1826 AND symb_decoder(16#d1#)) OR
 					(reg_q1826 AND symb_decoder(16#97#)) OR
 					(reg_q1826 AND symb_decoder(16#b1#)) OR
 					(reg_q1826 AND symb_decoder(16#9e#)) OR
 					(reg_q1826 AND symb_decoder(16#ec#)) OR
 					(reg_q1826 AND symb_decoder(16#2b#)) OR
 					(reg_q1826 AND symb_decoder(16#62#)) OR
 					(reg_q1826 AND symb_decoder(16#6e#)) OR
 					(reg_q1826 AND symb_decoder(16#d0#)) OR
 					(reg_q1826 AND symb_decoder(16#1a#)) OR
 					(reg_q1826 AND symb_decoder(16#02#)) OR
 					(reg_q1826 AND symb_decoder(16#19#)) OR
 					(reg_q1826 AND symb_decoder(16#d4#)) OR
 					(reg_q1826 AND symb_decoder(16#67#)) OR
 					(reg_q1826 AND symb_decoder(16#32#)) OR
 					(reg_q1826 AND symb_decoder(16#ff#)) OR
 					(reg_q1826 AND symb_decoder(16#cb#)) OR
 					(reg_q1826 AND symb_decoder(16#23#)) OR
 					(reg_q1826 AND symb_decoder(16#08#)) OR
 					(reg_q1826 AND symb_decoder(16#aa#)) OR
 					(reg_q1826 AND symb_decoder(16#3a#)) OR
 					(reg_q1826 AND symb_decoder(16#82#)) OR
 					(reg_q1826 AND symb_decoder(16#31#)) OR
 					(reg_q1826 AND symb_decoder(16#3e#)) OR
 					(reg_q1826 AND symb_decoder(16#5f#)) OR
 					(reg_q1826 AND symb_decoder(16#a5#)) OR
 					(reg_q1826 AND symb_decoder(16#a6#)) OR
 					(reg_q1826 AND symb_decoder(16#d5#)) OR
 					(reg_q1826 AND symb_decoder(16#f2#)) OR
 					(reg_q1826 AND symb_decoder(16#d8#)) OR
 					(reg_q1826 AND symb_decoder(16#71#)) OR
 					(reg_q1826 AND symb_decoder(16#65#)) OR
 					(reg_q1826 AND symb_decoder(16#1c#)) OR
 					(reg_q1826 AND symb_decoder(16#a9#)) OR
 					(reg_q1826 AND symb_decoder(16#e1#)) OR
 					(reg_q1826 AND symb_decoder(16#81#)) OR
 					(reg_q1826 AND symb_decoder(16#e9#)) OR
 					(reg_q1826 AND symb_decoder(16#47#)) OR
 					(reg_q1826 AND symb_decoder(16#9b#)) OR
 					(reg_q1826 AND symb_decoder(16#c3#)) OR
 					(reg_q1826 AND symb_decoder(16#5c#)) OR
 					(reg_q1826 AND symb_decoder(16#7b#)) OR
 					(reg_q1826 AND symb_decoder(16#2c#)) OR
 					(reg_q1826 AND symb_decoder(16#ee#)) OR
 					(reg_q1826 AND symb_decoder(16#5d#)) OR
 					(reg_q1826 AND symb_decoder(16#44#)) OR
 					(reg_q1826 AND symb_decoder(16#63#)) OR
 					(reg_q1826 AND symb_decoder(16#95#)) OR
 					(reg_q1826 AND symb_decoder(16#e0#)) OR
 					(reg_q1826 AND symb_decoder(16#6d#)) OR
 					(reg_q1826 AND symb_decoder(16#20#)) OR
 					(reg_q1826 AND symb_decoder(16#48#)) OR
 					(reg_q1826 AND symb_decoder(16#87#)) OR
 					(reg_q1826 AND symb_decoder(16#1b#)) OR
 					(reg_q1826 AND symb_decoder(16#01#)) OR
 					(reg_q1826 AND symb_decoder(16#3c#)) OR
 					(reg_q1826 AND symb_decoder(16#8f#)) OR
 					(reg_q1826 AND symb_decoder(16#38#)) OR
 					(reg_q1826 AND symb_decoder(16#b3#)) OR
 					(reg_q1826 AND symb_decoder(16#c1#)) OR
 					(reg_q1826 AND symb_decoder(16#7f#)) OR
 					(reg_q1826 AND symb_decoder(16#64#)) OR
 					(reg_q1826 AND symb_decoder(16#5e#)) OR
 					(reg_q1826 AND symb_decoder(16#b9#)) OR
 					(reg_q1826 AND symb_decoder(16#0d#)) OR
 					(reg_q1826 AND symb_decoder(16#c4#)) OR
 					(reg_q1826 AND symb_decoder(16#7a#)) OR
 					(reg_q1826 AND symb_decoder(16#3b#)) OR
 					(reg_q1826 AND symb_decoder(16#b6#)) OR
 					(reg_q1826 AND symb_decoder(16#e6#)) OR
 					(reg_q1826 AND symb_decoder(16#80#)) OR
 					(reg_q1826 AND symb_decoder(16#93#)) OR
 					(reg_q1826 AND symb_decoder(16#c6#)) OR
 					(reg_q1826 AND symb_decoder(16#76#)) OR
 					(reg_q1826 AND symb_decoder(16#54#)) OR
 					(reg_q1826 AND symb_decoder(16#24#)) OR
 					(reg_q1826 AND symb_decoder(16#fc#)) OR
 					(reg_q1826 AND symb_decoder(16#59#)) OR
 					(reg_q1826 AND symb_decoder(16#cf#)) OR
 					(reg_q1826 AND symb_decoder(16#9c#));
reg_q1826_init <= '0' ;
	p_reg_q1826: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1826 <= reg_q1826_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1826 <= reg_q1826_init;
        else
          reg_q1826 <= reg_q1826_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1452_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1452 AND symb_decoder(16#6d#)) OR
 					(reg_q1452 AND symb_decoder(16#55#)) OR
 					(reg_q1452 AND symb_decoder(16#ff#)) OR
 					(reg_q1452 AND symb_decoder(16#47#)) OR
 					(reg_q1452 AND symb_decoder(16#5f#)) OR
 					(reg_q1452 AND symb_decoder(16#6e#)) OR
 					(reg_q1452 AND symb_decoder(16#4a#)) OR
 					(reg_q1452 AND symb_decoder(16#5e#)) OR
 					(reg_q1452 AND symb_decoder(16#03#)) OR
 					(reg_q1452 AND symb_decoder(16#38#)) OR
 					(reg_q1452 AND symb_decoder(16#34#)) OR
 					(reg_q1452 AND symb_decoder(16#aa#)) OR
 					(reg_q1452 AND symb_decoder(16#5d#)) OR
 					(reg_q1452 AND symb_decoder(16#8b#)) OR
 					(reg_q1452 AND symb_decoder(16#0d#)) OR
 					(reg_q1452 AND symb_decoder(16#17#)) OR
 					(reg_q1452 AND symb_decoder(16#b9#)) OR
 					(reg_q1452 AND symb_decoder(16#0e#)) OR
 					(reg_q1452 AND symb_decoder(16#06#)) OR
 					(reg_q1452 AND symb_decoder(16#f7#)) OR
 					(reg_q1452 AND symb_decoder(16#59#)) OR
 					(reg_q1452 AND symb_decoder(16#c1#)) OR
 					(reg_q1452 AND symb_decoder(16#9d#)) OR
 					(reg_q1452 AND symb_decoder(16#3a#)) OR
 					(reg_q1452 AND symb_decoder(16#ab#)) OR
 					(reg_q1452 AND symb_decoder(16#79#)) OR
 					(reg_q1452 AND symb_decoder(16#a7#)) OR
 					(reg_q1452 AND symb_decoder(16#66#)) OR
 					(reg_q1452 AND symb_decoder(16#25#)) OR
 					(reg_q1452 AND symb_decoder(16#5a#)) OR
 					(reg_q1452 AND symb_decoder(16#b8#)) OR
 					(reg_q1452 AND symb_decoder(16#ef#)) OR
 					(reg_q1452 AND symb_decoder(16#84#)) OR
 					(reg_q1452 AND symb_decoder(16#de#)) OR
 					(reg_q1452 AND symb_decoder(16#02#)) OR
 					(reg_q1452 AND symb_decoder(16#86#)) OR
 					(reg_q1452 AND symb_decoder(16#f4#)) OR
 					(reg_q1452 AND symb_decoder(16#cc#)) OR
 					(reg_q1452 AND symb_decoder(16#35#)) OR
 					(reg_q1452 AND symb_decoder(16#ee#)) OR
 					(reg_q1452 AND symb_decoder(16#6c#)) OR
 					(reg_q1452 AND symb_decoder(16#ac#)) OR
 					(reg_q1452 AND symb_decoder(16#a5#)) OR
 					(reg_q1452 AND symb_decoder(16#39#)) OR
 					(reg_q1452 AND symb_decoder(16#73#)) OR
 					(reg_q1452 AND symb_decoder(16#4d#)) OR
 					(reg_q1452 AND symb_decoder(16#1c#)) OR
 					(reg_q1452 AND symb_decoder(16#1e#)) OR
 					(reg_q1452 AND symb_decoder(16#e0#)) OR
 					(reg_q1452 AND symb_decoder(16#83#)) OR
 					(reg_q1452 AND symb_decoder(16#cd#)) OR
 					(reg_q1452 AND symb_decoder(16#fa#)) OR
 					(reg_q1452 AND symb_decoder(16#da#)) OR
 					(reg_q1452 AND symb_decoder(16#30#)) OR
 					(reg_q1452 AND symb_decoder(16#fe#)) OR
 					(reg_q1452 AND symb_decoder(16#27#)) OR
 					(reg_q1452 AND symb_decoder(16#97#)) OR
 					(reg_q1452 AND symb_decoder(16#24#)) OR
 					(reg_q1452 AND symb_decoder(16#e4#)) OR
 					(reg_q1452 AND symb_decoder(16#bb#)) OR
 					(reg_q1452 AND symb_decoder(16#85#)) OR
 					(reg_q1452 AND symb_decoder(16#42#)) OR
 					(reg_q1452 AND symb_decoder(16#92#)) OR
 					(reg_q1452 AND symb_decoder(16#3c#)) OR
 					(reg_q1452 AND symb_decoder(16#a9#)) OR
 					(reg_q1452 AND symb_decoder(16#d0#)) OR
 					(reg_q1452 AND symb_decoder(16#6b#)) OR
 					(reg_q1452 AND symb_decoder(16#81#)) OR
 					(reg_q1452 AND symb_decoder(16#3d#)) OR
 					(reg_q1452 AND symb_decoder(16#a1#)) OR
 					(reg_q1452 AND symb_decoder(16#3b#)) OR
 					(reg_q1452 AND symb_decoder(16#7c#)) OR
 					(reg_q1452 AND symb_decoder(16#28#)) OR
 					(reg_q1452 AND symb_decoder(16#2e#)) OR
 					(reg_q1452 AND symb_decoder(16#b1#)) OR
 					(reg_q1452 AND symb_decoder(16#a0#)) OR
 					(reg_q1452 AND symb_decoder(16#2c#)) OR
 					(reg_q1452 AND symb_decoder(16#ba#)) OR
 					(reg_q1452 AND symb_decoder(16#3e#)) OR
 					(reg_q1452 AND symb_decoder(16#68#)) OR
 					(reg_q1452 AND symb_decoder(16#9b#)) OR
 					(reg_q1452 AND symb_decoder(16#c2#)) OR
 					(reg_q1452 AND symb_decoder(16#ae#)) OR
 					(reg_q1452 AND symb_decoder(16#0a#)) OR
 					(reg_q1452 AND symb_decoder(16#71#)) OR
 					(reg_q1452 AND symb_decoder(16#2b#)) OR
 					(reg_q1452 AND symb_decoder(16#df#)) OR
 					(reg_q1452 AND symb_decoder(16#00#)) OR
 					(reg_q1452 AND symb_decoder(16#07#)) OR
 					(reg_q1452 AND symb_decoder(16#8e#)) OR
 					(reg_q1452 AND symb_decoder(16#12#)) OR
 					(reg_q1452 AND symb_decoder(16#09#)) OR
 					(reg_q1452 AND symb_decoder(16#ec#)) OR
 					(reg_q1452 AND symb_decoder(16#82#)) OR
 					(reg_q1452 AND symb_decoder(16#c5#)) OR
 					(reg_q1452 AND symb_decoder(16#65#)) OR
 					(reg_q1452 AND symb_decoder(16#f1#)) OR
 					(reg_q1452 AND symb_decoder(16#2a#)) OR
 					(reg_q1452 AND symb_decoder(16#16#)) OR
 					(reg_q1452 AND symb_decoder(16#dc#)) OR
 					(reg_q1452 AND symb_decoder(16#e1#)) OR
 					(reg_q1452 AND symb_decoder(16#ad#)) OR
 					(reg_q1452 AND symb_decoder(16#60#)) OR
 					(reg_q1452 AND symb_decoder(16#14#)) OR
 					(reg_q1452 AND symb_decoder(16#56#)) OR
 					(reg_q1452 AND symb_decoder(16#04#)) OR
 					(reg_q1452 AND symb_decoder(16#b2#)) OR
 					(reg_q1452 AND symb_decoder(16#20#)) OR
 					(reg_q1452 AND symb_decoder(16#b3#)) OR
 					(reg_q1452 AND symb_decoder(16#f2#)) OR
 					(reg_q1452 AND symb_decoder(16#b7#)) OR
 					(reg_q1452 AND symb_decoder(16#c7#)) OR
 					(reg_q1452 AND symb_decoder(16#78#)) OR
 					(reg_q1452 AND symb_decoder(16#31#)) OR
 					(reg_q1452 AND symb_decoder(16#9c#)) OR
 					(reg_q1452 AND symb_decoder(16#63#)) OR
 					(reg_q1452 AND symb_decoder(16#f8#)) OR
 					(reg_q1452 AND symb_decoder(16#44#)) OR
 					(reg_q1452 AND symb_decoder(16#db#)) OR
 					(reg_q1452 AND symb_decoder(16#62#)) OR
 					(reg_q1452 AND symb_decoder(16#70#)) OR
 					(reg_q1452 AND symb_decoder(16#45#)) OR
 					(reg_q1452 AND symb_decoder(16#08#)) OR
 					(reg_q1452 AND symb_decoder(16#72#)) OR
 					(reg_q1452 AND symb_decoder(16#d9#)) OR
 					(reg_q1452 AND symb_decoder(16#e8#)) OR
 					(reg_q1452 AND symb_decoder(16#51#)) OR
 					(reg_q1452 AND symb_decoder(16#48#)) OR
 					(reg_q1452 AND symb_decoder(16#e5#)) OR
 					(reg_q1452 AND symb_decoder(16#f0#)) OR
 					(reg_q1452 AND symb_decoder(16#95#)) OR
 					(reg_q1452 AND symb_decoder(16#8f#)) OR
 					(reg_q1452 AND symb_decoder(16#01#)) OR
 					(reg_q1452 AND symb_decoder(16#2f#)) OR
 					(reg_q1452 AND symb_decoder(16#96#)) OR
 					(reg_q1452 AND symb_decoder(16#7d#)) OR
 					(reg_q1452 AND symb_decoder(16#cf#)) OR
 					(reg_q1452 AND symb_decoder(16#15#)) OR
 					(reg_q1452 AND symb_decoder(16#c3#)) OR
 					(reg_q1452 AND symb_decoder(16#a4#)) OR
 					(reg_q1452 AND symb_decoder(16#57#)) OR
 					(reg_q1452 AND symb_decoder(16#29#)) OR
 					(reg_q1452 AND symb_decoder(16#ea#)) OR
 					(reg_q1452 AND symb_decoder(16#c4#)) OR
 					(reg_q1452 AND symb_decoder(16#9a#)) OR
 					(reg_q1452 AND symb_decoder(16#c6#)) OR
 					(reg_q1452 AND symb_decoder(16#41#)) OR
 					(reg_q1452 AND symb_decoder(16#69#)) OR
 					(reg_q1452 AND symb_decoder(16#4c#)) OR
 					(reg_q1452 AND symb_decoder(16#4f#)) OR
 					(reg_q1452 AND symb_decoder(16#10#)) OR
 					(reg_q1452 AND symb_decoder(16#2d#)) OR
 					(reg_q1452 AND symb_decoder(16#32#)) OR
 					(reg_q1452 AND symb_decoder(16#26#)) OR
 					(reg_q1452 AND symb_decoder(16#94#)) OR
 					(reg_q1452 AND symb_decoder(16#50#)) OR
 					(reg_q1452 AND symb_decoder(16#d2#)) OR
 					(reg_q1452 AND symb_decoder(16#80#)) OR
 					(reg_q1452 AND symb_decoder(16#11#)) OR
 					(reg_q1452 AND symb_decoder(16#89#)) OR
 					(reg_q1452 AND symb_decoder(16#61#)) OR
 					(reg_q1452 AND symb_decoder(16#75#)) OR
 					(reg_q1452 AND symb_decoder(16#d6#)) OR
 					(reg_q1452 AND symb_decoder(16#d8#)) OR
 					(reg_q1452 AND symb_decoder(16#76#)) OR
 					(reg_q1452 AND symb_decoder(16#ca#)) OR
 					(reg_q1452 AND symb_decoder(16#88#)) OR
 					(reg_q1452 AND symb_decoder(16#22#)) OR
 					(reg_q1452 AND symb_decoder(16#cb#)) OR
 					(reg_q1452 AND symb_decoder(16#4b#)) OR
 					(reg_q1452 AND symb_decoder(16#52#)) OR
 					(reg_q1452 AND symb_decoder(16#e6#)) OR
 					(reg_q1452 AND symb_decoder(16#a2#)) OR
 					(reg_q1452 AND symb_decoder(16#0b#)) OR
 					(reg_q1452 AND symb_decoder(16#f6#)) OR
 					(reg_q1452 AND symb_decoder(16#46#)) OR
 					(reg_q1452 AND symb_decoder(16#90#)) OR
 					(reg_q1452 AND symb_decoder(16#f3#)) OR
 					(reg_q1452 AND symb_decoder(16#99#)) OR
 					(reg_q1452 AND symb_decoder(16#be#)) OR
 					(reg_q1452 AND symb_decoder(16#98#)) OR
 					(reg_q1452 AND symb_decoder(16#13#)) OR
 					(reg_q1452 AND symb_decoder(16#c8#)) OR
 					(reg_q1452 AND symb_decoder(16#8d#)) OR
 					(reg_q1452 AND symb_decoder(16#67#)) OR
 					(reg_q1452 AND symb_decoder(16#d4#)) OR
 					(reg_q1452 AND symb_decoder(16#e2#)) OR
 					(reg_q1452 AND symb_decoder(16#21#)) OR
 					(reg_q1452 AND symb_decoder(16#43#)) OR
 					(reg_q1452 AND symb_decoder(16#87#)) OR
 					(reg_q1452 AND symb_decoder(16#7b#)) OR
 					(reg_q1452 AND symb_decoder(16#7a#)) OR
 					(reg_q1452 AND symb_decoder(16#a3#)) OR
 					(reg_q1452 AND symb_decoder(16#58#)) OR
 					(reg_q1452 AND symb_decoder(16#05#)) OR
 					(reg_q1452 AND symb_decoder(16#4e#)) OR
 					(reg_q1452 AND symb_decoder(16#eb#)) OR
 					(reg_q1452 AND symb_decoder(16#9f#)) OR
 					(reg_q1452 AND symb_decoder(16#53#)) OR
 					(reg_q1452 AND symb_decoder(16#8a#)) OR
 					(reg_q1452 AND symb_decoder(16#93#)) OR
 					(reg_q1452 AND symb_decoder(16#37#)) OR
 					(reg_q1452 AND symb_decoder(16#a6#)) OR
 					(reg_q1452 AND symb_decoder(16#fb#)) OR
 					(reg_q1452 AND symb_decoder(16#d7#)) OR
 					(reg_q1452 AND symb_decoder(16#f9#)) OR
 					(reg_q1452 AND symb_decoder(16#74#)) OR
 					(reg_q1452 AND symb_decoder(16#b0#)) OR
 					(reg_q1452 AND symb_decoder(16#6f#)) OR
 					(reg_q1452 AND symb_decoder(16#b4#)) OR
 					(reg_q1452 AND symb_decoder(16#64#)) OR
 					(reg_q1452 AND symb_decoder(16#bf#)) OR
 					(reg_q1452 AND symb_decoder(16#b6#)) OR
 					(reg_q1452 AND symb_decoder(16#8c#)) OR
 					(reg_q1452 AND symb_decoder(16#33#)) OR
 					(reg_q1452 AND symb_decoder(16#77#)) OR
 					(reg_q1452 AND symb_decoder(16#c0#)) OR
 					(reg_q1452 AND symb_decoder(16#fd#)) OR
 					(reg_q1452 AND symb_decoder(16#1d#)) OR
 					(reg_q1452 AND symb_decoder(16#6a#)) OR
 					(reg_q1452 AND symb_decoder(16#c9#)) OR
 					(reg_q1452 AND symb_decoder(16#ed#)) OR
 					(reg_q1452 AND symb_decoder(16#d3#)) OR
 					(reg_q1452 AND symb_decoder(16#23#)) OR
 					(reg_q1452 AND symb_decoder(16#40#)) OR
 					(reg_q1452 AND symb_decoder(16#bc#)) OR
 					(reg_q1452 AND symb_decoder(16#1b#)) OR
 					(reg_q1452 AND symb_decoder(16#36#)) OR
 					(reg_q1452 AND symb_decoder(16#5c#)) OR
 					(reg_q1452 AND symb_decoder(16#91#)) OR
 					(reg_q1452 AND symb_decoder(16#e9#)) OR
 					(reg_q1452 AND symb_decoder(16#d1#)) OR
 					(reg_q1452 AND symb_decoder(16#dd#)) OR
 					(reg_q1452 AND symb_decoder(16#0f#)) OR
 					(reg_q1452 AND symb_decoder(16#5b#)) OR
 					(reg_q1452 AND symb_decoder(16#b5#)) OR
 					(reg_q1452 AND symb_decoder(16#7e#)) OR
 					(reg_q1452 AND symb_decoder(16#9e#)) OR
 					(reg_q1452 AND symb_decoder(16#ce#)) OR
 					(reg_q1452 AND symb_decoder(16#af#)) OR
 					(reg_q1452 AND symb_decoder(16#d5#)) OR
 					(reg_q1452 AND symb_decoder(16#49#)) OR
 					(reg_q1452 AND symb_decoder(16#1f#)) OR
 					(reg_q1452 AND symb_decoder(16#0c#)) OR
 					(reg_q1452 AND symb_decoder(16#bd#)) OR
 					(reg_q1452 AND symb_decoder(16#a8#)) OR
 					(reg_q1452 AND symb_decoder(16#54#)) OR
 					(reg_q1452 AND symb_decoder(16#e7#)) OR
 					(reg_q1452 AND symb_decoder(16#f5#)) OR
 					(reg_q1452 AND symb_decoder(16#19#)) OR
 					(reg_q1452 AND symb_decoder(16#e3#)) OR
 					(reg_q1452 AND symb_decoder(16#7f#)) OR
 					(reg_q1452 AND symb_decoder(16#1a#)) OR
 					(reg_q1452 AND symb_decoder(16#18#)) OR
 					(reg_q1452 AND symb_decoder(16#fc#)) OR
 					(reg_q1452 AND symb_decoder(16#3f#));
reg_q1452_init <= '0' ;
	p_reg_q1452: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1452 <= reg_q1452_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1452 <= reg_q1452_init;
        else
          reg_q1452 <= reg_q1452_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q958_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q958 AND symb_decoder(16#46#)) OR
 					(reg_q958 AND symb_decoder(16#18#)) OR
 					(reg_q958 AND symb_decoder(16#01#)) OR
 					(reg_q958 AND symb_decoder(16#86#)) OR
 					(reg_q958 AND symb_decoder(16#61#)) OR
 					(reg_q958 AND symb_decoder(16#c9#)) OR
 					(reg_q958 AND symb_decoder(16#9a#)) OR
 					(reg_q958 AND symb_decoder(16#76#)) OR
 					(reg_q958 AND symb_decoder(16#36#)) OR
 					(reg_q958 AND symb_decoder(16#e3#)) OR
 					(reg_q958 AND symb_decoder(16#95#)) OR
 					(reg_q958 AND symb_decoder(16#ba#)) OR
 					(reg_q958 AND symb_decoder(16#13#)) OR
 					(reg_q958 AND symb_decoder(16#f3#)) OR
 					(reg_q958 AND symb_decoder(16#e5#)) OR
 					(reg_q958 AND symb_decoder(16#07#)) OR
 					(reg_q958 AND symb_decoder(16#91#)) OR
 					(reg_q958 AND symb_decoder(16#a6#)) OR
 					(reg_q958 AND symb_decoder(16#39#)) OR
 					(reg_q958 AND symb_decoder(16#02#)) OR
 					(reg_q958 AND symb_decoder(16#d8#)) OR
 					(reg_q958 AND symb_decoder(16#70#)) OR
 					(reg_q958 AND symb_decoder(16#5b#)) OR
 					(reg_q958 AND symb_decoder(16#92#)) OR
 					(reg_q958 AND symb_decoder(16#1c#)) OR
 					(reg_q958 AND symb_decoder(16#f6#)) OR
 					(reg_q958 AND symb_decoder(16#a5#)) OR
 					(reg_q958 AND symb_decoder(16#b7#)) OR
 					(reg_q958 AND symb_decoder(16#03#)) OR
 					(reg_q958 AND symb_decoder(16#52#)) OR
 					(reg_q958 AND symb_decoder(16#3e#)) OR
 					(reg_q958 AND symb_decoder(16#b8#)) OR
 					(reg_q958 AND symb_decoder(16#40#)) OR
 					(reg_q958 AND symb_decoder(16#45#)) OR
 					(reg_q958 AND symb_decoder(16#51#)) OR
 					(reg_q958 AND symb_decoder(16#1b#)) OR
 					(reg_q958 AND symb_decoder(16#e2#)) OR
 					(reg_q958 AND symb_decoder(16#da#)) OR
 					(reg_q958 AND symb_decoder(16#fc#)) OR
 					(reg_q958 AND symb_decoder(16#33#)) OR
 					(reg_q958 AND symb_decoder(16#f4#)) OR
 					(reg_q958 AND symb_decoder(16#78#)) OR
 					(reg_q958 AND symb_decoder(16#96#)) OR
 					(reg_q958 AND symb_decoder(16#e4#)) OR
 					(reg_q958 AND symb_decoder(16#42#)) OR
 					(reg_q958 AND symb_decoder(16#62#)) OR
 					(reg_q958 AND symb_decoder(16#c4#)) OR
 					(reg_q958 AND symb_decoder(16#04#)) OR
 					(reg_q958 AND symb_decoder(16#b6#)) OR
 					(reg_q958 AND symb_decoder(16#db#)) OR
 					(reg_q958 AND symb_decoder(16#23#)) OR
 					(reg_q958 AND symb_decoder(16#fa#)) OR
 					(reg_q958 AND symb_decoder(16#19#)) OR
 					(reg_q958 AND symb_decoder(16#6b#)) OR
 					(reg_q958 AND symb_decoder(16#67#)) OR
 					(reg_q958 AND symb_decoder(16#d1#)) OR
 					(reg_q958 AND symb_decoder(16#0d#)) OR
 					(reg_q958 AND symb_decoder(16#fb#)) OR
 					(reg_q958 AND symb_decoder(16#5f#)) OR
 					(reg_q958 AND symb_decoder(16#c2#)) OR
 					(reg_q958 AND symb_decoder(16#4c#)) OR
 					(reg_q958 AND symb_decoder(16#6a#)) OR
 					(reg_q958 AND symb_decoder(16#d6#)) OR
 					(reg_q958 AND symb_decoder(16#26#)) OR
 					(reg_q958 AND symb_decoder(16#5d#)) OR
 					(reg_q958 AND symb_decoder(16#09#)) OR
 					(reg_q958 AND symb_decoder(16#9c#)) OR
 					(reg_q958 AND symb_decoder(16#c0#)) OR
 					(reg_q958 AND symb_decoder(16#ef#)) OR
 					(reg_q958 AND symb_decoder(16#11#)) OR
 					(reg_q958 AND symb_decoder(16#af#)) OR
 					(reg_q958 AND symb_decoder(16#f7#)) OR
 					(reg_q958 AND symb_decoder(16#57#)) OR
 					(reg_q958 AND symb_decoder(16#2c#)) OR
 					(reg_q958 AND symb_decoder(16#aa#)) OR
 					(reg_q958 AND symb_decoder(16#be#)) OR
 					(reg_q958 AND symb_decoder(16#71#)) OR
 					(reg_q958 AND symb_decoder(16#06#)) OR
 					(reg_q958 AND symb_decoder(16#d7#)) OR
 					(reg_q958 AND symb_decoder(16#94#)) OR
 					(reg_q958 AND symb_decoder(16#8b#)) OR
 					(reg_q958 AND symb_decoder(16#1f#)) OR
 					(reg_q958 AND symb_decoder(16#0b#)) OR
 					(reg_q958 AND symb_decoder(16#3f#)) OR
 					(reg_q958 AND symb_decoder(16#d0#)) OR
 					(reg_q958 AND symb_decoder(16#34#)) OR
 					(reg_q958 AND symb_decoder(16#f8#)) OR
 					(reg_q958 AND symb_decoder(16#14#)) OR
 					(reg_q958 AND symb_decoder(16#8d#)) OR
 					(reg_q958 AND symb_decoder(16#ca#)) OR
 					(reg_q958 AND symb_decoder(16#5a#)) OR
 					(reg_q958 AND symb_decoder(16#69#)) OR
 					(reg_q958 AND symb_decoder(16#64#)) OR
 					(reg_q958 AND symb_decoder(16#97#)) OR
 					(reg_q958 AND symb_decoder(16#e9#)) OR
 					(reg_q958 AND symb_decoder(16#dc#)) OR
 					(reg_q958 AND symb_decoder(16#c6#)) OR
 					(reg_q958 AND symb_decoder(16#fe#)) OR
 					(reg_q958 AND symb_decoder(16#53#)) OR
 					(reg_q958 AND symb_decoder(16#7c#)) OR
 					(reg_q958 AND symb_decoder(16#a7#)) OR
 					(reg_q958 AND symb_decoder(16#47#)) OR
 					(reg_q958 AND symb_decoder(16#4b#)) OR
 					(reg_q958 AND symb_decoder(16#15#)) OR
 					(reg_q958 AND symb_decoder(16#c8#)) OR
 					(reg_q958 AND symb_decoder(16#f2#)) OR
 					(reg_q958 AND symb_decoder(16#ad#)) OR
 					(reg_q958 AND symb_decoder(16#4a#)) OR
 					(reg_q958 AND symb_decoder(16#9f#)) OR
 					(reg_q958 AND symb_decoder(16#bd#)) OR
 					(reg_q958 AND symb_decoder(16#7b#)) OR
 					(reg_q958 AND symb_decoder(16#ae#)) OR
 					(reg_q958 AND symb_decoder(16#b4#)) OR
 					(reg_q958 AND symb_decoder(16#37#)) OR
 					(reg_q958 AND symb_decoder(16#28#)) OR
 					(reg_q958 AND symb_decoder(16#d3#)) OR
 					(reg_q958 AND symb_decoder(16#ab#)) OR
 					(reg_q958 AND symb_decoder(16#b0#)) OR
 					(reg_q958 AND symb_decoder(16#b3#)) OR
 					(reg_q958 AND symb_decoder(16#a4#)) OR
 					(reg_q958 AND symb_decoder(16#8a#)) OR
 					(reg_q958 AND symb_decoder(16#79#)) OR
 					(reg_q958 AND symb_decoder(16#50#)) OR
 					(reg_q958 AND symb_decoder(16#1e#)) OR
 					(reg_q958 AND symb_decoder(16#5e#)) OR
 					(reg_q958 AND symb_decoder(16#12#)) OR
 					(reg_q958 AND symb_decoder(16#2b#)) OR
 					(reg_q958 AND symb_decoder(16#a0#)) OR
 					(reg_q958 AND symb_decoder(16#16#)) OR
 					(reg_q958 AND symb_decoder(16#41#)) OR
 					(reg_q958 AND symb_decoder(16#63#)) OR
 					(reg_q958 AND symb_decoder(16#83#)) OR
 					(reg_q958 AND symb_decoder(16#30#)) OR
 					(reg_q958 AND symb_decoder(16#e8#)) OR
 					(reg_q958 AND symb_decoder(16#a1#)) OR
 					(reg_q958 AND symb_decoder(16#84#)) OR
 					(reg_q958 AND symb_decoder(16#ea#)) OR
 					(reg_q958 AND symb_decoder(16#d2#)) OR
 					(reg_q958 AND symb_decoder(16#54#)) OR
 					(reg_q958 AND symb_decoder(16#f5#)) OR
 					(reg_q958 AND symb_decoder(16#a8#)) OR
 					(reg_q958 AND symb_decoder(16#29#)) OR
 					(reg_q958 AND symb_decoder(16#c5#)) OR
 					(reg_q958 AND symb_decoder(16#74#)) OR
 					(reg_q958 AND symb_decoder(16#e0#)) OR
 					(reg_q958 AND symb_decoder(16#7a#)) OR
 					(reg_q958 AND symb_decoder(16#0a#)) OR
 					(reg_q958 AND symb_decoder(16#6e#)) OR
 					(reg_q958 AND symb_decoder(16#2d#)) OR
 					(reg_q958 AND symb_decoder(16#65#)) OR
 					(reg_q958 AND symb_decoder(16#3c#)) OR
 					(reg_q958 AND symb_decoder(16#c7#)) OR
 					(reg_q958 AND symb_decoder(16#e6#)) OR
 					(reg_q958 AND symb_decoder(16#56#)) OR
 					(reg_q958 AND symb_decoder(16#8e#)) OR
 					(reg_q958 AND symb_decoder(16#25#)) OR
 					(reg_q958 AND symb_decoder(16#38#)) OR
 					(reg_q958 AND symb_decoder(16#eb#)) OR
 					(reg_q958 AND symb_decoder(16#9d#)) OR
 					(reg_q958 AND symb_decoder(16#f0#)) OR
 					(reg_q958 AND symb_decoder(16#cc#)) OR
 					(reg_q958 AND symb_decoder(16#0e#)) OR
 					(reg_q958 AND symb_decoder(16#a9#)) OR
 					(reg_q958 AND symb_decoder(16#87#)) OR
 					(reg_q958 AND symb_decoder(16#81#)) OR
 					(reg_q958 AND symb_decoder(16#df#)) OR
 					(reg_q958 AND symb_decoder(16#ff#)) OR
 					(reg_q958 AND symb_decoder(16#21#)) OR
 					(reg_q958 AND symb_decoder(16#d5#)) OR
 					(reg_q958 AND symb_decoder(16#dd#)) OR
 					(reg_q958 AND symb_decoder(16#59#)) OR
 					(reg_q958 AND symb_decoder(16#e1#)) OR
 					(reg_q958 AND symb_decoder(16#7e#)) OR
 					(reg_q958 AND symb_decoder(16#17#)) OR
 					(reg_q958 AND symb_decoder(16#2f#)) OR
 					(reg_q958 AND symb_decoder(16#60#)) OR
 					(reg_q958 AND symb_decoder(16#6c#)) OR
 					(reg_q958 AND symb_decoder(16#05#)) OR
 					(reg_q958 AND symb_decoder(16#a3#)) OR
 					(reg_q958 AND symb_decoder(16#7d#)) OR
 					(reg_q958 AND symb_decoder(16#80#)) OR
 					(reg_q958 AND symb_decoder(16#1a#)) OR
 					(reg_q958 AND symb_decoder(16#77#)) OR
 					(reg_q958 AND symb_decoder(16#a2#)) OR
 					(reg_q958 AND symb_decoder(16#72#)) OR
 					(reg_q958 AND symb_decoder(16#85#)) OR
 					(reg_q958 AND symb_decoder(16#88#)) OR
 					(reg_q958 AND symb_decoder(16#98#)) OR
 					(reg_q958 AND symb_decoder(16#8c#)) OR
 					(reg_q958 AND symb_decoder(16#ee#)) OR
 					(reg_q958 AND symb_decoder(16#1d#)) OR
 					(reg_q958 AND symb_decoder(16#b2#)) OR
 					(reg_q958 AND symb_decoder(16#f9#)) OR
 					(reg_q958 AND symb_decoder(16#75#)) OR
 					(reg_q958 AND symb_decoder(16#89#)) OR
 					(reg_q958 AND symb_decoder(16#c1#)) OR
 					(reg_q958 AND symb_decoder(16#fd#)) OR
 					(reg_q958 AND symb_decoder(16#35#)) OR
 					(reg_q958 AND symb_decoder(16#9e#)) OR
 					(reg_q958 AND symb_decoder(16#ec#)) OR
 					(reg_q958 AND symb_decoder(16#27#)) OR
 					(reg_q958 AND symb_decoder(16#32#)) OR
 					(reg_q958 AND symb_decoder(16#cf#)) OR
 					(reg_q958 AND symb_decoder(16#44#)) OR
 					(reg_q958 AND symb_decoder(16#7f#)) OR
 					(reg_q958 AND symb_decoder(16#0c#)) OR
 					(reg_q958 AND symb_decoder(16#08#)) OR
 					(reg_q958 AND symb_decoder(16#d4#)) OR
 					(reg_q958 AND symb_decoder(16#d9#)) OR
 					(reg_q958 AND symb_decoder(16#68#)) OR
 					(reg_q958 AND symb_decoder(16#43#)) OR
 					(reg_q958 AND symb_decoder(16#cd#)) OR
 					(reg_q958 AND symb_decoder(16#0f#)) OR
 					(reg_q958 AND symb_decoder(16#8f#)) OR
 					(reg_q958 AND symb_decoder(16#bf#)) OR
 					(reg_q958 AND symb_decoder(16#3d#)) OR
 					(reg_q958 AND symb_decoder(16#82#)) OR
 					(reg_q958 AND symb_decoder(16#9b#)) OR
 					(reg_q958 AND symb_decoder(16#f1#)) OR
 					(reg_q958 AND symb_decoder(16#20#)) OR
 					(reg_q958 AND symb_decoder(16#2e#)) OR
 					(reg_q958 AND symb_decoder(16#3b#)) OR
 					(reg_q958 AND symb_decoder(16#6d#)) OR
 					(reg_q958 AND symb_decoder(16#93#)) OR
 					(reg_q958 AND symb_decoder(16#ce#)) OR
 					(reg_q958 AND symb_decoder(16#90#)) OR
 					(reg_q958 AND symb_decoder(16#b9#)) OR
 					(reg_q958 AND symb_decoder(16#31#)) OR
 					(reg_q958 AND symb_decoder(16#4e#)) OR
 					(reg_q958 AND symb_decoder(16#ac#)) OR
 					(reg_q958 AND symb_decoder(16#48#)) OR
 					(reg_q958 AND symb_decoder(16#cb#)) OR
 					(reg_q958 AND symb_decoder(16#bb#)) OR
 					(reg_q958 AND symb_decoder(16#49#)) OR
 					(reg_q958 AND symb_decoder(16#3a#)) OR
 					(reg_q958 AND symb_decoder(16#00#)) OR
 					(reg_q958 AND symb_decoder(16#73#)) OR
 					(reg_q958 AND symb_decoder(16#c3#)) OR
 					(reg_q958 AND symb_decoder(16#ed#)) OR
 					(reg_q958 AND symb_decoder(16#22#)) OR
 					(reg_q958 AND symb_decoder(16#6f#)) OR
 					(reg_q958 AND symb_decoder(16#4d#)) OR
 					(reg_q958 AND symb_decoder(16#2a#)) OR
 					(reg_q958 AND symb_decoder(16#10#)) OR
 					(reg_q958 AND symb_decoder(16#24#)) OR
 					(reg_q958 AND symb_decoder(16#58#)) OR
 					(reg_q958 AND symb_decoder(16#99#)) OR
 					(reg_q958 AND symb_decoder(16#b5#)) OR
 					(reg_q958 AND symb_decoder(16#b1#)) OR
 					(reg_q958 AND symb_decoder(16#55#)) OR
 					(reg_q958 AND symb_decoder(16#66#)) OR
 					(reg_q958 AND symb_decoder(16#de#)) OR
 					(reg_q958 AND symb_decoder(16#bc#)) OR
 					(reg_q958 AND symb_decoder(16#4f#)) OR
 					(reg_q958 AND symb_decoder(16#e7#)) OR
 					(reg_q958 AND symb_decoder(16#5c#));
reg_q958_init <= '0' ;
	p_reg_q958: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q958 <= reg_q958_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q958 <= reg_q958_init;
        else
          reg_q958 <= reg_q958_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2211_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2211 AND symb_decoder(16#43#)) OR
 					(reg_q2211 AND symb_decoder(16#18#)) OR
 					(reg_q2211 AND symb_decoder(16#a8#)) OR
 					(reg_q2211 AND symb_decoder(16#8d#)) OR
 					(reg_q2211 AND symb_decoder(16#d7#)) OR
 					(reg_q2211 AND symb_decoder(16#6b#)) OR
 					(reg_q2211 AND symb_decoder(16#93#)) OR
 					(reg_q2211 AND symb_decoder(16#a7#)) OR
 					(reg_q2211 AND symb_decoder(16#ce#)) OR
 					(reg_q2211 AND symb_decoder(16#d4#)) OR
 					(reg_q2211 AND symb_decoder(16#f1#)) OR
 					(reg_q2211 AND symb_decoder(16#85#)) OR
 					(reg_q2211 AND symb_decoder(16#ec#)) OR
 					(reg_q2211 AND symb_decoder(16#b9#)) OR
 					(reg_q2211 AND symb_decoder(16#df#)) OR
 					(reg_q2211 AND symb_decoder(16#ed#)) OR
 					(reg_q2211 AND symb_decoder(16#f3#)) OR
 					(reg_q2211 AND symb_decoder(16#4b#)) OR
 					(reg_q2211 AND symb_decoder(16#ae#)) OR
 					(reg_q2211 AND symb_decoder(16#8c#)) OR
 					(reg_q2211 AND symb_decoder(16#3b#)) OR
 					(reg_q2211 AND symb_decoder(16#3e#)) OR
 					(reg_q2211 AND symb_decoder(16#8e#)) OR
 					(reg_q2211 AND symb_decoder(16#31#)) OR
 					(reg_q2211 AND symb_decoder(16#2b#)) OR
 					(reg_q2211 AND symb_decoder(16#2e#)) OR
 					(reg_q2211 AND symb_decoder(16#84#)) OR
 					(reg_q2211 AND symb_decoder(16#20#)) OR
 					(reg_q2211 AND symb_decoder(16#92#)) OR
 					(reg_q2211 AND symb_decoder(16#7f#)) OR
 					(reg_q2211 AND symb_decoder(16#1b#)) OR
 					(reg_q2211 AND symb_decoder(16#d6#)) OR
 					(reg_q2211 AND symb_decoder(16#88#)) OR
 					(reg_q2211 AND symb_decoder(16#be#)) OR
 					(reg_q2211 AND symb_decoder(16#2a#)) OR
 					(reg_q2211 AND symb_decoder(16#1c#)) OR
 					(reg_q2211 AND symb_decoder(16#61#)) OR
 					(reg_q2211 AND symb_decoder(16#a1#)) OR
 					(reg_q2211 AND symb_decoder(16#53#)) OR
 					(reg_q2211 AND symb_decoder(16#d5#)) OR
 					(reg_q2211 AND symb_decoder(16#23#)) OR
 					(reg_q2211 AND symb_decoder(16#4d#)) OR
 					(reg_q2211 AND symb_decoder(16#f8#)) OR
 					(reg_q2211 AND symb_decoder(16#f5#)) OR
 					(reg_q2211 AND symb_decoder(16#e2#)) OR
 					(reg_q2211 AND symb_decoder(16#9a#)) OR
 					(reg_q2211 AND symb_decoder(16#65#)) OR
 					(reg_q2211 AND symb_decoder(16#c9#)) OR
 					(reg_q2211 AND symb_decoder(16#75#)) OR
 					(reg_q2211 AND symb_decoder(16#9b#)) OR
 					(reg_q2211 AND symb_decoder(16#8f#)) OR
 					(reg_q2211 AND symb_decoder(16#09#)) OR
 					(reg_q2211 AND symb_decoder(16#d2#)) OR
 					(reg_q2211 AND symb_decoder(16#dc#)) OR
 					(reg_q2211 AND symb_decoder(16#41#)) OR
 					(reg_q2211 AND symb_decoder(16#3c#)) OR
 					(reg_q2211 AND symb_decoder(16#24#)) OR
 					(reg_q2211 AND symb_decoder(16#6f#)) OR
 					(reg_q2211 AND symb_decoder(16#c4#)) OR
 					(reg_q2211 AND symb_decoder(16#81#)) OR
 					(reg_q2211 AND symb_decoder(16#b0#)) OR
 					(reg_q2211 AND symb_decoder(16#b7#)) OR
 					(reg_q2211 AND symb_decoder(16#9f#)) OR
 					(reg_q2211 AND symb_decoder(16#91#)) OR
 					(reg_q2211 AND symb_decoder(16#c5#)) OR
 					(reg_q2211 AND symb_decoder(16#48#)) OR
 					(reg_q2211 AND symb_decoder(16#7e#)) OR
 					(reg_q2211 AND symb_decoder(16#15#)) OR
 					(reg_q2211 AND symb_decoder(16#00#)) OR
 					(reg_q2211 AND symb_decoder(16#2d#)) OR
 					(reg_q2211 AND symb_decoder(16#5e#)) OR
 					(reg_q2211 AND symb_decoder(16#05#)) OR
 					(reg_q2211 AND symb_decoder(16#42#)) OR
 					(reg_q2211 AND symb_decoder(16#db#)) OR
 					(reg_q2211 AND symb_decoder(16#a9#)) OR
 					(reg_q2211 AND symb_decoder(16#4f#)) OR
 					(reg_q2211 AND symb_decoder(16#72#)) OR
 					(reg_q2211 AND symb_decoder(16#30#)) OR
 					(reg_q2211 AND symb_decoder(16#59#)) OR
 					(reg_q2211 AND symb_decoder(16#e9#)) OR
 					(reg_q2211 AND symb_decoder(16#ea#)) OR
 					(reg_q2211 AND symb_decoder(16#08#)) OR
 					(reg_q2211 AND symb_decoder(16#b2#)) OR
 					(reg_q2211 AND symb_decoder(16#57#)) OR
 					(reg_q2211 AND symb_decoder(16#9c#)) OR
 					(reg_q2211 AND symb_decoder(16#07#)) OR
 					(reg_q2211 AND symb_decoder(16#b3#)) OR
 					(reg_q2211 AND symb_decoder(16#32#)) OR
 					(reg_q2211 AND symb_decoder(16#ad#)) OR
 					(reg_q2211 AND symb_decoder(16#ee#)) OR
 					(reg_q2211 AND symb_decoder(16#35#)) OR
 					(reg_q2211 AND symb_decoder(16#0e#)) OR
 					(reg_q2211 AND symb_decoder(16#45#)) OR
 					(reg_q2211 AND symb_decoder(16#36#)) OR
 					(reg_q2211 AND symb_decoder(16#95#)) OR
 					(reg_q2211 AND symb_decoder(16#02#)) OR
 					(reg_q2211 AND symb_decoder(16#9d#)) OR
 					(reg_q2211 AND symb_decoder(16#0b#)) OR
 					(reg_q2211 AND symb_decoder(16#b1#)) OR
 					(reg_q2211 AND symb_decoder(16#27#)) OR
 					(reg_q2211 AND symb_decoder(16#d0#)) OR
 					(reg_q2211 AND symb_decoder(16#e5#)) OR
 					(reg_q2211 AND symb_decoder(16#51#)) OR
 					(reg_q2211 AND symb_decoder(16#c3#)) OR
 					(reg_q2211 AND symb_decoder(16#0a#)) OR
 					(reg_q2211 AND symb_decoder(16#11#)) OR
 					(reg_q2211 AND symb_decoder(16#2f#)) OR
 					(reg_q2211 AND symb_decoder(16#01#)) OR
 					(reg_q2211 AND symb_decoder(16#3d#)) OR
 					(reg_q2211 AND symb_decoder(16#82#)) OR
 					(reg_q2211 AND symb_decoder(16#4e#)) OR
 					(reg_q2211 AND symb_decoder(16#99#)) OR
 					(reg_q2211 AND symb_decoder(16#fb#)) OR
 					(reg_q2211 AND symb_decoder(16#5a#)) OR
 					(reg_q2211 AND symb_decoder(16#83#)) OR
 					(reg_q2211 AND symb_decoder(16#58#)) OR
 					(reg_q2211 AND symb_decoder(16#64#)) OR
 					(reg_q2211 AND symb_decoder(16#a3#)) OR
 					(reg_q2211 AND symb_decoder(16#bd#)) OR
 					(reg_q2211 AND symb_decoder(16#5d#)) OR
 					(reg_q2211 AND symb_decoder(16#d9#)) OR
 					(reg_q2211 AND symb_decoder(16#03#)) OR
 					(reg_q2211 AND symb_decoder(16#d1#)) OR
 					(reg_q2211 AND symb_decoder(16#d3#)) OR
 					(reg_q2211 AND symb_decoder(16#5b#)) OR
 					(reg_q2211 AND symb_decoder(16#bf#)) OR
 					(reg_q2211 AND symb_decoder(16#c1#)) OR
 					(reg_q2211 AND symb_decoder(16#f9#)) OR
 					(reg_q2211 AND symb_decoder(16#67#)) OR
 					(reg_q2211 AND symb_decoder(16#80#)) OR
 					(reg_q2211 AND symb_decoder(16#6e#)) OR
 					(reg_q2211 AND symb_decoder(16#7a#)) OR
 					(reg_q2211 AND symb_decoder(16#a0#)) OR
 					(reg_q2211 AND symb_decoder(16#90#)) OR
 					(reg_q2211 AND symb_decoder(16#66#)) OR
 					(reg_q2211 AND symb_decoder(16#fc#)) OR
 					(reg_q2211 AND symb_decoder(16#60#)) OR
 					(reg_q2211 AND symb_decoder(16#21#)) OR
 					(reg_q2211 AND symb_decoder(16#49#)) OR
 					(reg_q2211 AND symb_decoder(16#29#)) OR
 					(reg_q2211 AND symb_decoder(16#af#)) OR
 					(reg_q2211 AND symb_decoder(16#a6#)) OR
 					(reg_q2211 AND symb_decoder(16#5f#)) OR
 					(reg_q2211 AND symb_decoder(16#ef#)) OR
 					(reg_q2211 AND symb_decoder(16#b6#)) OR
 					(reg_q2211 AND symb_decoder(16#f4#)) OR
 					(reg_q2211 AND symb_decoder(16#46#)) OR
 					(reg_q2211 AND symb_decoder(16#71#)) OR
 					(reg_q2211 AND symb_decoder(16#89#)) OR
 					(reg_q2211 AND symb_decoder(16#f0#)) OR
 					(reg_q2211 AND symb_decoder(16#5c#)) OR
 					(reg_q2211 AND symb_decoder(16#26#)) OR
 					(reg_q2211 AND symb_decoder(16#e0#)) OR
 					(reg_q2211 AND symb_decoder(16#56#)) OR
 					(reg_q2211 AND symb_decoder(16#55#)) OR
 					(reg_q2211 AND symb_decoder(16#4c#)) OR
 					(reg_q2211 AND symb_decoder(16#06#)) OR
 					(reg_q2211 AND symb_decoder(16#b5#)) OR
 					(reg_q2211 AND symb_decoder(16#f7#)) OR
 					(reg_q2211 AND symb_decoder(16#78#)) OR
 					(reg_q2211 AND symb_decoder(16#12#)) OR
 					(reg_q2211 AND symb_decoder(16#a2#)) OR
 					(reg_q2211 AND symb_decoder(16#eb#)) OR
 					(reg_q2211 AND symb_decoder(16#6c#)) OR
 					(reg_q2211 AND symb_decoder(16#50#)) OR
 					(reg_q2211 AND symb_decoder(16#39#)) OR
 					(reg_q2211 AND symb_decoder(16#25#)) OR
 					(reg_q2211 AND symb_decoder(16#ff#)) OR
 					(reg_q2211 AND symb_decoder(16#1f#)) OR
 					(reg_q2211 AND symb_decoder(16#de#)) OR
 					(reg_q2211 AND symb_decoder(16#e7#)) OR
 					(reg_q2211 AND symb_decoder(16#62#)) OR
 					(reg_q2211 AND symb_decoder(16#40#)) OR
 					(reg_q2211 AND symb_decoder(16#ab#)) OR
 					(reg_q2211 AND symb_decoder(16#7c#)) OR
 					(reg_q2211 AND symb_decoder(16#22#)) OR
 					(reg_q2211 AND symb_decoder(16#10#)) OR
 					(reg_q2211 AND symb_decoder(16#68#)) OR
 					(reg_q2211 AND symb_decoder(16#98#)) OR
 					(reg_q2211 AND symb_decoder(16#c8#)) OR
 					(reg_q2211 AND symb_decoder(16#44#)) OR
 					(reg_q2211 AND symb_decoder(16#37#)) OR
 					(reg_q2211 AND symb_decoder(16#fe#)) OR
 					(reg_q2211 AND symb_decoder(16#69#)) OR
 					(reg_q2211 AND symb_decoder(16#cc#)) OR
 					(reg_q2211 AND symb_decoder(16#86#)) OR
 					(reg_q2211 AND symb_decoder(16#9e#)) OR
 					(reg_q2211 AND symb_decoder(16#b8#)) OR
 					(reg_q2211 AND symb_decoder(16#a5#)) OR
 					(reg_q2211 AND symb_decoder(16#cf#)) OR
 					(reg_q2211 AND symb_decoder(16#47#)) OR
 					(reg_q2211 AND symb_decoder(16#6d#)) OR
 					(reg_q2211 AND symb_decoder(16#3f#)) OR
 					(reg_q2211 AND symb_decoder(16#e8#)) OR
 					(reg_q2211 AND symb_decoder(16#34#)) OR
 					(reg_q2211 AND symb_decoder(16#e6#)) OR
 					(reg_q2211 AND symb_decoder(16#38#)) OR
 					(reg_q2211 AND symb_decoder(16#77#)) OR
 					(reg_q2211 AND symb_decoder(16#fd#)) OR
 					(reg_q2211 AND symb_decoder(16#ca#)) OR
 					(reg_q2211 AND symb_decoder(16#1d#)) OR
 					(reg_q2211 AND symb_decoder(16#c7#)) OR
 					(reg_q2211 AND symb_decoder(16#c6#)) OR
 					(reg_q2211 AND symb_decoder(16#16#)) OR
 					(reg_q2211 AND symb_decoder(16#e4#)) OR
 					(reg_q2211 AND symb_decoder(16#da#)) OR
 					(reg_q2211 AND symb_decoder(16#1e#)) OR
 					(reg_q2211 AND symb_decoder(16#2c#)) OR
 					(reg_q2211 AND symb_decoder(16#cb#)) OR
 					(reg_q2211 AND symb_decoder(16#52#)) OR
 					(reg_q2211 AND symb_decoder(16#17#)) OR
 					(reg_q2211 AND symb_decoder(16#b4#)) OR
 					(reg_q2211 AND symb_decoder(16#28#)) OR
 					(reg_q2211 AND symb_decoder(16#74#)) OR
 					(reg_q2211 AND symb_decoder(16#6a#)) OR
 					(reg_q2211 AND symb_decoder(16#4a#)) OR
 					(reg_q2211 AND symb_decoder(16#c2#)) OR
 					(reg_q2211 AND symb_decoder(16#13#)) OR
 					(reg_q2211 AND symb_decoder(16#96#)) OR
 					(reg_q2211 AND symb_decoder(16#e1#)) OR
 					(reg_q2211 AND symb_decoder(16#1a#)) OR
 					(reg_q2211 AND symb_decoder(16#dd#)) OR
 					(reg_q2211 AND symb_decoder(16#ac#)) OR
 					(reg_q2211 AND symb_decoder(16#8b#)) OR
 					(reg_q2211 AND symb_decoder(16#f2#)) OR
 					(reg_q2211 AND symb_decoder(16#73#)) OR
 					(reg_q2211 AND symb_decoder(16#cd#)) OR
 					(reg_q2211 AND symb_decoder(16#94#)) OR
 					(reg_q2211 AND symb_decoder(16#19#)) OR
 					(reg_q2211 AND symb_decoder(16#bb#)) OR
 					(reg_q2211 AND symb_decoder(16#04#)) OR
 					(reg_q2211 AND symb_decoder(16#63#)) OR
 					(reg_q2211 AND symb_decoder(16#54#)) OR
 					(reg_q2211 AND symb_decoder(16#e3#)) OR
 					(reg_q2211 AND symb_decoder(16#76#)) OR
 					(reg_q2211 AND symb_decoder(16#3a#)) OR
 					(reg_q2211 AND symb_decoder(16#f6#)) OR
 					(reg_q2211 AND symb_decoder(16#87#)) OR
 					(reg_q2211 AND symb_decoder(16#79#)) OR
 					(reg_q2211 AND symb_decoder(16#c0#)) OR
 					(reg_q2211 AND symb_decoder(16#aa#)) OR
 					(reg_q2211 AND symb_decoder(16#0f#)) OR
 					(reg_q2211 AND symb_decoder(16#0c#)) OR
 					(reg_q2211 AND symb_decoder(16#d8#)) OR
 					(reg_q2211 AND symb_decoder(16#14#)) OR
 					(reg_q2211 AND symb_decoder(16#7d#)) OR
 					(reg_q2211 AND symb_decoder(16#a4#)) OR
 					(reg_q2211 AND symb_decoder(16#33#)) OR
 					(reg_q2211 AND symb_decoder(16#0d#)) OR
 					(reg_q2211 AND symb_decoder(16#97#)) OR
 					(reg_q2211 AND symb_decoder(16#8a#)) OR
 					(reg_q2211 AND symb_decoder(16#bc#)) OR
 					(reg_q2211 AND symb_decoder(16#7b#)) OR
 					(reg_q2211 AND symb_decoder(16#ba#)) OR
 					(reg_q2211 AND symb_decoder(16#70#)) OR
 					(reg_q2211 AND symb_decoder(16#fa#));
reg_q2211_init <= '0' ;
	p_reg_q2211: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2211 <= reg_q2211_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2211 <= reg_q2211_init;
        else
          reg_q2211 <= reg_q2211_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q0_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q0 AND symb_decoder(16#b3#)) OR
 					(reg_q0 AND symb_decoder(16#2b#)) OR
 					(reg_q0 AND symb_decoder(16#34#)) OR
 					(reg_q0 AND symb_decoder(16#3a#)) OR
 					(reg_q0 AND symb_decoder(16#90#)) OR
 					(reg_q0 AND symb_decoder(16#e9#)) OR
 					(reg_q0 AND symb_decoder(16#d3#)) OR
 					(reg_q0 AND symb_decoder(16#d4#)) OR
 					(reg_q0 AND symb_decoder(16#32#)) OR
 					(reg_q0 AND symb_decoder(16#e7#)) OR
 					(reg_q0 AND symb_decoder(16#51#)) OR
 					(reg_q0 AND symb_decoder(16#67#)) OR
 					(reg_q0 AND symb_decoder(16#91#)) OR
 					(reg_q0 AND symb_decoder(16#7e#)) OR
 					(reg_q0 AND symb_decoder(16#53#)) OR
 					(reg_q0 AND symb_decoder(16#6a#)) OR
 					(reg_q0 AND symb_decoder(16#a4#)) OR
 					(reg_q0 AND symb_decoder(16#f9#)) OR
 					(reg_q0 AND symb_decoder(16#bc#)) OR
 					(reg_q0 AND symb_decoder(16#11#)) OR
 					(reg_q0 AND symb_decoder(16#10#)) OR
 					(reg_q0 AND symb_decoder(16#01#)) OR
 					(reg_q0 AND symb_decoder(16#ba#)) OR
 					(reg_q0 AND symb_decoder(16#50#)) OR
 					(reg_q0 AND symb_decoder(16#e4#)) OR
 					(reg_q0 AND symb_decoder(16#65#)) OR
 					(reg_q0 AND symb_decoder(16#e5#)) OR
 					(reg_q0 AND symb_decoder(16#87#)) OR
 					(reg_q0 AND symb_decoder(16#2e#)) OR
 					(reg_q0 AND symb_decoder(16#9b#)) OR
 					(reg_q0 AND symb_decoder(16#c3#)) OR
 					(reg_q0 AND symb_decoder(16#40#)) OR
 					(reg_q0 AND symb_decoder(16#0e#)) OR
 					(reg_q0 AND symb_decoder(16#98#)) OR
 					(reg_q0 AND symb_decoder(16#b8#)) OR
 					(reg_q0 AND symb_decoder(16#60#)) OR
 					(reg_q0 AND symb_decoder(16#52#)) OR
 					(reg_q0 AND symb_decoder(16#22#)) OR
 					(reg_q0 AND symb_decoder(16#5a#)) OR
 					(reg_q0 AND symb_decoder(16#31#)) OR
 					(reg_q0 AND symb_decoder(16#a8#)) OR
 					(reg_q0 AND symb_decoder(16#f8#)) OR
 					(reg_q0 AND symb_decoder(16#80#)) OR
 					(reg_q0 AND symb_decoder(16#77#)) OR
 					(reg_q0 AND symb_decoder(16#ca#)) OR
 					(reg_q0 AND symb_decoder(16#fa#)) OR
 					(reg_q0 AND symb_decoder(16#c2#)) OR
 					(reg_q0 AND symb_decoder(16#ea#)) OR
 					(reg_q0 AND symb_decoder(16#5b#)) OR
 					(reg_q0 AND symb_decoder(16#16#)) OR
 					(reg_q0 AND symb_decoder(16#c1#)) OR
 					(reg_q0 AND symb_decoder(16#9c#)) OR
 					(reg_q0 AND symb_decoder(16#9d#)) OR
 					(reg_q0 AND symb_decoder(16#62#)) OR
 					(reg_q0 AND symb_decoder(16#a7#)) OR
 					(reg_q0 AND symb_decoder(16#b0#)) OR
 					(reg_q0 AND symb_decoder(16#5e#)) OR
 					(reg_q0 AND symb_decoder(16#a1#)) OR
 					(reg_q0 AND symb_decoder(16#fb#)) OR
 					(reg_q0 AND symb_decoder(16#9f#)) OR
 					(reg_q0 AND symb_decoder(16#4e#)) OR
 					(reg_q0 AND symb_decoder(16#2f#)) OR
 					(reg_q0 AND symb_decoder(16#74#)) OR
 					(reg_q0 AND symb_decoder(16#8b#)) OR
 					(reg_q0 AND symb_decoder(16#bf#)) OR
 					(reg_q0 AND symb_decoder(16#8f#)) OR
 					(reg_q0 AND symb_decoder(16#20#)) OR
 					(reg_q0 AND symb_decoder(16#3e#)) OR
 					(reg_q0 AND symb_decoder(16#39#)) OR
 					(reg_q0 AND symb_decoder(16#89#)) OR
 					(reg_q0 AND symb_decoder(16#e8#)) OR
 					(reg_q0 AND symb_decoder(16#5d#)) OR
 					(reg_q0 AND symb_decoder(16#a0#)) OR
 					(reg_q0 AND symb_decoder(16#fd#)) OR
 					(reg_q0 AND symb_decoder(16#ec#)) OR
 					(reg_q0 AND symb_decoder(16#cd#)) OR
 					(reg_q0 AND symb_decoder(16#4a#)) OR
 					(reg_q0 AND symb_decoder(16#a3#)) OR
 					(reg_q0 AND symb_decoder(16#6f#)) OR
 					(reg_q0 AND symb_decoder(16#08#)) OR
 					(reg_q0 AND symb_decoder(16#ff#)) OR
 					(reg_q0 AND symb_decoder(16#c7#)) OR
 					(reg_q0 AND symb_decoder(16#cb#)) OR
 					(reg_q0 AND symb_decoder(16#48#)) OR
 					(reg_q0 AND symb_decoder(16#1d#)) OR
 					(reg_q0 AND symb_decoder(16#a5#)) OR
 					(reg_q0 AND symb_decoder(16#1f#)) OR
 					(reg_q0 AND symb_decoder(16#1e#)) OR
 					(reg_q0 AND symb_decoder(16#47#)) OR
 					(reg_q0 AND symb_decoder(16#64#)) OR
 					(reg_q0 AND symb_decoder(16#f6#)) OR
 					(reg_q0 AND symb_decoder(16#6d#)) OR
 					(reg_q0 AND symb_decoder(16#84#)) OR
 					(reg_q0 AND symb_decoder(16#f1#)) OR
 					(reg_q0 AND symb_decoder(16#03#)) OR
 					(reg_q0 AND symb_decoder(16#46#)) OR
 					(reg_q0 AND symb_decoder(16#6b#)) OR
 					(reg_q0 AND symb_decoder(16#02#)) OR
 					(reg_q0 AND symb_decoder(16#88#)) OR
 					(reg_q0 AND symb_decoder(16#bd#)) OR
 					(reg_q0 AND symb_decoder(16#49#)) OR
 					(reg_q0 AND symb_decoder(16#21#)) OR
 					(reg_q0 AND symb_decoder(16#f5#)) OR
 					(reg_q0 AND symb_decoder(16#25#)) OR
 					(reg_q0 AND symb_decoder(16#c6#)) OR
 					(reg_q0 AND symb_decoder(16#97#)) OR
 					(reg_q0 AND symb_decoder(16#d5#)) OR
 					(reg_q0 AND symb_decoder(16#71#)) OR
 					(reg_q0 AND symb_decoder(16#66#)) OR
 					(reg_q0 AND symb_decoder(16#12#)) OR
 					(reg_q0 AND symb_decoder(16#ee#)) OR
 					(reg_q0 AND symb_decoder(16#35#)) OR
 					(reg_q0 AND symb_decoder(16#59#)) OR
 					(reg_q0 AND symb_decoder(16#81#)) OR
 					(reg_q0 AND symb_decoder(16#99#)) OR
 					(reg_q0 AND symb_decoder(16#2d#)) OR
 					(reg_q0 AND symb_decoder(16#ad#)) OR
 					(reg_q0 AND symb_decoder(16#c4#)) OR
 					(reg_q0 AND symb_decoder(16#83#)) OR
 					(reg_q0 AND symb_decoder(16#61#)) OR
 					(reg_q0 AND symb_decoder(16#e1#)) OR
 					(reg_q0 AND symb_decoder(16#4d#)) OR
 					(reg_q0 AND symb_decoder(16#30#)) OR
 					(reg_q0 AND symb_decoder(16#a9#)) OR
 					(reg_q0 AND symb_decoder(16#4b#)) OR
 					(reg_q0 AND symb_decoder(16#da#)) OR
 					(reg_q0 AND symb_decoder(16#9e#)) OR
 					(reg_q0 AND symb_decoder(16#7b#)) OR
 					(reg_q0 AND symb_decoder(16#f2#)) OR
 					(reg_q0 AND symb_decoder(16#9a#)) OR
 					(reg_q0 AND symb_decoder(16#33#)) OR
 					(reg_q0 AND symb_decoder(16#4c#)) OR
 					(reg_q0 AND symb_decoder(16#78#)) OR
 					(reg_q0 AND symb_decoder(16#18#)) OR
 					(reg_q0 AND symb_decoder(16#ef#)) OR
 					(reg_q0 AND symb_decoder(16#3d#)) OR
 					(reg_q0 AND symb_decoder(16#dc#)) OR
 					(reg_q0 AND symb_decoder(16#cc#)) OR
 					(reg_q0 AND symb_decoder(16#a2#)) OR
 					(reg_q0 AND symb_decoder(16#41#)) OR
 					(reg_q0 AND symb_decoder(16#23#)) OR
 					(reg_q0 AND symb_decoder(16#b4#)) OR
 					(reg_q0 AND symb_decoder(16#38#)) OR
 					(reg_q0 AND symb_decoder(16#75#)) OR
 					(reg_q0 AND symb_decoder(16#56#)) OR
 					(reg_q0 AND symb_decoder(16#af#)) OR
 					(reg_q0 AND symb_decoder(16#8e#)) OR
 					(reg_q0 AND symb_decoder(16#55#)) OR
 					(reg_q0 AND symb_decoder(16#cf#)) OR
 					(reg_q0 AND symb_decoder(16#f7#)) OR
 					(reg_q0 AND symb_decoder(16#a6#)) OR
 					(reg_q0 AND symb_decoder(16#76#)) OR
 					(reg_q0 AND symb_decoder(16#1b#)) OR
 					(reg_q0 AND symb_decoder(16#00#)) OR
 					(reg_q0 AND symb_decoder(16#09#)) OR
 					(reg_q0 AND symb_decoder(16#7f#)) OR
 					(reg_q0 AND symb_decoder(16#d1#)) OR
 					(reg_q0 AND symb_decoder(16#17#)) OR
 					(reg_q0 AND symb_decoder(16#c8#)) OR
 					(reg_q0 AND symb_decoder(16#d2#)) OR
 					(reg_q0 AND symb_decoder(16#29#)) OR
 					(reg_q0 AND symb_decoder(16#ac#)) OR
 					(reg_q0 AND symb_decoder(16#94#)) OR
 					(reg_q0 AND symb_decoder(16#86#)) OR
 					(reg_q0 AND symb_decoder(16#ae#)) OR
 					(reg_q0 AND symb_decoder(16#14#)) OR
 					(reg_q0 AND symb_decoder(16#b2#)) OR
 					(reg_q0 AND symb_decoder(16#b1#)) OR
 					(reg_q0 AND symb_decoder(16#ed#)) OR
 					(reg_q0 AND symb_decoder(16#d7#)) OR
 					(reg_q0 AND symb_decoder(16#44#)) OR
 					(reg_q0 AND symb_decoder(16#5c#)) OR
 					(reg_q0 AND symb_decoder(16#06#)) OR
 					(reg_q0 AND symb_decoder(16#19#)) OR
 					(reg_q0 AND symb_decoder(16#c0#)) OR
 					(reg_q0 AND symb_decoder(16#fe#)) OR
 					(reg_q0 AND symb_decoder(16#fc#)) OR
 					(reg_q0 AND symb_decoder(16#05#)) OR
 					(reg_q0 AND symb_decoder(16#3f#)) OR
 					(reg_q0 AND symb_decoder(16#1c#)) OR
 					(reg_q0 AND symb_decoder(16#7c#)) OR
 					(reg_q0 AND symb_decoder(16#e2#)) OR
 					(reg_q0 AND symb_decoder(16#6c#)) OR
 					(reg_q0 AND symb_decoder(16#e0#)) OR
 					(reg_q0 AND symb_decoder(16#36#)) OR
 					(reg_q0 AND symb_decoder(16#aa#)) OR
 					(reg_q0 AND symb_decoder(16#27#)) OR
 					(reg_q0 AND symb_decoder(16#d8#)) OR
 					(reg_q0 AND symb_decoder(16#73#)) OR
 					(reg_q0 AND symb_decoder(16#eb#)) OR
 					(reg_q0 AND symb_decoder(16#85#)) OR
 					(reg_q0 AND symb_decoder(16#54#)) OR
 					(reg_q0 AND symb_decoder(16#69#)) OR
 					(reg_q0 AND symb_decoder(16#13#)) OR
 					(reg_q0 AND symb_decoder(16#f0#)) OR
 					(reg_q0 AND symb_decoder(16#57#)) OR
 					(reg_q0 AND symb_decoder(16#e3#)) OR
 					(reg_q0 AND symb_decoder(16#0a#)) OR
 					(reg_q0 AND symb_decoder(16#42#)) OR
 					(reg_q0 AND symb_decoder(16#95#)) OR
 					(reg_q0 AND symb_decoder(16#b5#)) OR
 					(reg_q0 AND symb_decoder(16#ce#)) OR
 					(reg_q0 AND symb_decoder(16#c5#)) OR
 					(reg_q0 AND symb_decoder(16#26#)) OR
 					(reg_q0 AND symb_decoder(16#96#)) OR
 					(reg_q0 AND symb_decoder(16#63#)) OR
 					(reg_q0 AND symb_decoder(16#ab#)) OR
 					(reg_q0 AND symb_decoder(16#04#)) OR
 					(reg_q0 AND symb_decoder(16#b6#)) OR
 					(reg_q0 AND symb_decoder(16#7a#)) OR
 					(reg_q0 AND symb_decoder(16#0d#)) OR
 					(reg_q0 AND symb_decoder(16#93#)) OR
 					(reg_q0 AND symb_decoder(16#68#)) OR
 					(reg_q0 AND symb_decoder(16#0b#)) OR
 					(reg_q0 AND symb_decoder(16#d6#)) OR
 					(reg_q0 AND symb_decoder(16#b7#)) OR
 					(reg_q0 AND symb_decoder(16#2a#)) OR
 					(reg_q0 AND symb_decoder(16#24#)) OR
 					(reg_q0 AND symb_decoder(16#3c#)) OR
 					(reg_q0 AND symb_decoder(16#3b#)) OR
 					(reg_q0 AND symb_decoder(16#2c#)) OR
 					(reg_q0 AND symb_decoder(16#43#)) OR
 					(reg_q0 AND symb_decoder(16#37#)) OR
 					(reg_q0 AND symb_decoder(16#de#)) OR
 					(reg_q0 AND symb_decoder(16#f3#)) OR
 					(reg_q0 AND symb_decoder(16#c9#)) OR
 					(reg_q0 AND symb_decoder(16#db#)) OR
 					(reg_q0 AND symb_decoder(16#45#)) OR
 					(reg_q0 AND symb_decoder(16#be#)) OR
 					(reg_q0 AND symb_decoder(16#d0#)) OR
 					(reg_q0 AND symb_decoder(16#79#)) OR
 					(reg_q0 AND symb_decoder(16#58#)) OR
 					(reg_q0 AND symb_decoder(16#0f#)) OR
 					(reg_q0 AND symb_decoder(16#8a#)) OR
 					(reg_q0 AND symb_decoder(16#dd#)) OR
 					(reg_q0 AND symb_decoder(16#d9#)) OR
 					(reg_q0 AND symb_decoder(16#07#)) OR
 					(reg_q0 AND symb_decoder(16#28#)) OR
 					(reg_q0 AND symb_decoder(16#1a#)) OR
 					(reg_q0 AND symb_decoder(16#8d#)) OR
 					(reg_q0 AND symb_decoder(16#6e#)) OR
 					(reg_q0 AND symb_decoder(16#8c#)) OR
 					(reg_q0 AND symb_decoder(16#e6#)) OR
 					(reg_q0 AND symb_decoder(16#0c#)) OR
 					(reg_q0 AND symb_decoder(16#70#)) OR
 					(reg_q0 AND symb_decoder(16#15#)) OR
 					(reg_q0 AND symb_decoder(16#92#)) OR
 					(reg_q0 AND symb_decoder(16#bb#)) OR
 					(reg_q0 AND symb_decoder(16#df#)) OR
 					(reg_q0 AND symb_decoder(16#b9#)) OR
 					(reg_q0 AND symb_decoder(16#72#)) OR
 					(reg_q0 AND symb_decoder(16#7d#)) OR
 					(reg_q0 AND symb_decoder(16#5f#)) OR
 					(reg_q0 AND symb_decoder(16#f4#)) OR
 					(reg_q0 AND symb_decoder(16#4f#)) OR
 					(reg_q0 AND symb_decoder(16#82#));
reg_q0_init <= '0' ;
	p_reg_q0: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q0 <= reg_q0_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q0 <= reg_q0_init;
        else
          reg_q0 <= reg_q0_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q303_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q303 AND symb_decoder(16#1c#)) OR
 					(reg_q303 AND symb_decoder(16#26#)) OR
 					(reg_q303 AND symb_decoder(16#77#)) OR
 					(reg_q303 AND symb_decoder(16#95#)) OR
 					(reg_q303 AND symb_decoder(16#86#)) OR
 					(reg_q303 AND symb_decoder(16#53#)) OR
 					(reg_q303 AND symb_decoder(16#5d#)) OR
 					(reg_q303 AND symb_decoder(16#ac#)) OR
 					(reg_q303 AND symb_decoder(16#07#)) OR
 					(reg_q303 AND symb_decoder(16#af#)) OR
 					(reg_q303 AND symb_decoder(16#4b#)) OR
 					(reg_q303 AND symb_decoder(16#de#)) OR
 					(reg_q303 AND symb_decoder(16#9b#)) OR
 					(reg_q303 AND symb_decoder(16#41#)) OR
 					(reg_q303 AND symb_decoder(16#02#)) OR
 					(reg_q303 AND symb_decoder(16#58#)) OR
 					(reg_q303 AND symb_decoder(16#12#)) OR
 					(reg_q303 AND symb_decoder(16#01#)) OR
 					(reg_q303 AND symb_decoder(16#ce#)) OR
 					(reg_q303 AND symb_decoder(16#dd#)) OR
 					(reg_q303 AND symb_decoder(16#70#)) OR
 					(reg_q303 AND symb_decoder(16#e8#)) OR
 					(reg_q303 AND symb_decoder(16#27#)) OR
 					(reg_q303 AND symb_decoder(16#cf#)) OR
 					(reg_q303 AND symb_decoder(16#ec#)) OR
 					(reg_q303 AND symb_decoder(16#f2#)) OR
 					(reg_q303 AND symb_decoder(16#7d#)) OR
 					(reg_q303 AND symb_decoder(16#46#)) OR
 					(reg_q303 AND symb_decoder(16#a3#)) OR
 					(reg_q303 AND symb_decoder(16#3b#)) OR
 					(reg_q303 AND symb_decoder(16#35#)) OR
 					(reg_q303 AND symb_decoder(16#d7#)) OR
 					(reg_q303 AND symb_decoder(16#2a#)) OR
 					(reg_q303 AND symb_decoder(16#df#)) OR
 					(reg_q303 AND symb_decoder(16#f5#)) OR
 					(reg_q303 AND symb_decoder(16#55#)) OR
 					(reg_q303 AND symb_decoder(16#36#)) OR
 					(reg_q303 AND symb_decoder(16#72#)) OR
 					(reg_q303 AND symb_decoder(16#3c#)) OR
 					(reg_q303 AND symb_decoder(16#43#)) OR
 					(reg_q303 AND symb_decoder(16#bc#)) OR
 					(reg_q303 AND symb_decoder(16#11#)) OR
 					(reg_q303 AND symb_decoder(16#fe#)) OR
 					(reg_q303 AND symb_decoder(16#6e#)) OR
 					(reg_q303 AND symb_decoder(16#33#)) OR
 					(reg_q303 AND symb_decoder(16#23#)) OR
 					(reg_q303 AND symb_decoder(16#c9#)) OR
 					(reg_q303 AND symb_decoder(16#24#)) OR
 					(reg_q303 AND symb_decoder(16#e6#)) OR
 					(reg_q303 AND symb_decoder(16#a7#)) OR
 					(reg_q303 AND symb_decoder(16#b9#)) OR
 					(reg_q303 AND symb_decoder(16#f8#)) OR
 					(reg_q303 AND symb_decoder(16#34#)) OR
 					(reg_q303 AND symb_decoder(16#88#)) OR
 					(reg_q303 AND symb_decoder(16#81#)) OR
 					(reg_q303 AND symb_decoder(16#c1#)) OR
 					(reg_q303 AND symb_decoder(16#d5#)) OR
 					(reg_q303 AND symb_decoder(16#3d#)) OR
 					(reg_q303 AND symb_decoder(16#32#)) OR
 					(reg_q303 AND symb_decoder(16#4a#)) OR
 					(reg_q303 AND symb_decoder(16#ff#)) OR
 					(reg_q303 AND symb_decoder(16#5c#)) OR
 					(reg_q303 AND symb_decoder(16#60#)) OR
 					(reg_q303 AND symb_decoder(16#b7#)) OR
 					(reg_q303 AND symb_decoder(16#fd#)) OR
 					(reg_q303 AND symb_decoder(16#eb#)) OR
 					(reg_q303 AND symb_decoder(16#21#)) OR
 					(reg_q303 AND symb_decoder(16#5a#)) OR
 					(reg_q303 AND symb_decoder(16#f7#)) OR
 					(reg_q303 AND symb_decoder(16#59#)) OR
 					(reg_q303 AND symb_decoder(16#18#)) OR
 					(reg_q303 AND symb_decoder(16#13#)) OR
 					(reg_q303 AND symb_decoder(16#56#)) OR
 					(reg_q303 AND symb_decoder(16#ab#)) OR
 					(reg_q303 AND symb_decoder(16#dc#)) OR
 					(reg_q303 AND symb_decoder(16#8b#)) OR
 					(reg_q303 AND symb_decoder(16#68#)) OR
 					(reg_q303 AND symb_decoder(16#76#)) OR
 					(reg_q303 AND symb_decoder(16#b0#)) OR
 					(reg_q303 AND symb_decoder(16#47#)) OR
 					(reg_q303 AND symb_decoder(16#92#)) OR
 					(reg_q303 AND symb_decoder(16#93#)) OR
 					(reg_q303 AND symb_decoder(16#e4#)) OR
 					(reg_q303 AND symb_decoder(16#2d#)) OR
 					(reg_q303 AND symb_decoder(16#7a#)) OR
 					(reg_q303 AND symb_decoder(16#90#)) OR
 					(reg_q303 AND symb_decoder(16#03#)) OR
 					(reg_q303 AND symb_decoder(16#5e#)) OR
 					(reg_q303 AND symb_decoder(16#d3#)) OR
 					(reg_q303 AND symb_decoder(16#84#)) OR
 					(reg_q303 AND symb_decoder(16#f6#)) OR
 					(reg_q303 AND symb_decoder(16#04#)) OR
 					(reg_q303 AND symb_decoder(16#1b#)) OR
 					(reg_q303 AND symb_decoder(16#d2#)) OR
 					(reg_q303 AND symb_decoder(16#c6#)) OR
 					(reg_q303 AND symb_decoder(16#49#)) OR
 					(reg_q303 AND symb_decoder(16#e2#)) OR
 					(reg_q303 AND symb_decoder(16#b4#)) OR
 					(reg_q303 AND symb_decoder(16#d1#)) OR
 					(reg_q303 AND symb_decoder(16#3f#)) OR
 					(reg_q303 AND symb_decoder(16#1d#)) OR
 					(reg_q303 AND symb_decoder(16#c3#)) OR
 					(reg_q303 AND symb_decoder(16#c4#)) OR
 					(reg_q303 AND symb_decoder(16#50#)) OR
 					(reg_q303 AND symb_decoder(16#5b#)) OR
 					(reg_q303 AND symb_decoder(16#1a#)) OR
 					(reg_q303 AND symb_decoder(16#f4#)) OR
 					(reg_q303 AND symb_decoder(16#15#)) OR
 					(reg_q303 AND symb_decoder(16#d0#)) OR
 					(reg_q303 AND symb_decoder(16#f1#)) OR
 					(reg_q303 AND symb_decoder(16#97#)) OR
 					(reg_q303 AND symb_decoder(16#85#)) OR
 					(reg_q303 AND symb_decoder(16#67#)) OR
 					(reg_q303 AND symb_decoder(16#ee#)) OR
 					(reg_q303 AND symb_decoder(16#0c#)) OR
 					(reg_q303 AND symb_decoder(16#96#)) OR
 					(reg_q303 AND symb_decoder(16#8e#)) OR
 					(reg_q303 AND symb_decoder(16#2e#)) OR
 					(reg_q303 AND symb_decoder(16#4d#)) OR
 					(reg_q303 AND symb_decoder(16#ae#)) OR
 					(reg_q303 AND symb_decoder(16#0a#)) OR
 					(reg_q303 AND symb_decoder(16#16#)) OR
 					(reg_q303 AND symb_decoder(16#8f#)) OR
 					(reg_q303 AND symb_decoder(16#78#)) OR
 					(reg_q303 AND symb_decoder(16#74#)) OR
 					(reg_q303 AND symb_decoder(16#a9#)) OR
 					(reg_q303 AND symb_decoder(16#bd#)) OR
 					(reg_q303 AND symb_decoder(16#c7#)) OR
 					(reg_q303 AND symb_decoder(16#30#)) OR
 					(reg_q303 AND symb_decoder(16#00#)) OR
 					(reg_q303 AND symb_decoder(16#c0#)) OR
 					(reg_q303 AND symb_decoder(16#19#)) OR
 					(reg_q303 AND symb_decoder(16#bb#)) OR
 					(reg_q303 AND symb_decoder(16#7e#)) OR
 					(reg_q303 AND symb_decoder(16#38#)) OR
 					(reg_q303 AND symb_decoder(16#0b#)) OR
 					(reg_q303 AND symb_decoder(16#8d#)) OR
 					(reg_q303 AND symb_decoder(16#7b#)) OR
 					(reg_q303 AND symb_decoder(16#45#)) OR
 					(reg_q303 AND symb_decoder(16#e0#)) OR
 					(reg_q303 AND symb_decoder(16#22#)) OR
 					(reg_q303 AND symb_decoder(16#6b#)) OR
 					(reg_q303 AND symb_decoder(16#87#)) OR
 					(reg_q303 AND symb_decoder(16#d8#)) OR
 					(reg_q303 AND symb_decoder(16#9f#)) OR
 					(reg_q303 AND symb_decoder(16#d9#)) OR
 					(reg_q303 AND symb_decoder(16#fb#)) OR
 					(reg_q303 AND symb_decoder(16#62#)) OR
 					(reg_q303 AND symb_decoder(16#cc#)) OR
 					(reg_q303 AND symb_decoder(16#9d#)) OR
 					(reg_q303 AND symb_decoder(16#a1#)) OR
 					(reg_q303 AND symb_decoder(16#65#)) OR
 					(reg_q303 AND symb_decoder(16#0f#)) OR
 					(reg_q303 AND symb_decoder(16#6a#)) OR
 					(reg_q303 AND symb_decoder(16#6d#)) OR
 					(reg_q303 AND symb_decoder(16#63#)) OR
 					(reg_q303 AND symb_decoder(16#05#)) OR
 					(reg_q303 AND symb_decoder(16#ef#)) OR
 					(reg_q303 AND symb_decoder(16#79#)) OR
 					(reg_q303 AND symb_decoder(16#a5#)) OR
 					(reg_q303 AND symb_decoder(16#17#)) OR
 					(reg_q303 AND symb_decoder(16#da#)) OR
 					(reg_q303 AND symb_decoder(16#6c#)) OR
 					(reg_q303 AND symb_decoder(16#cb#)) OR
 					(reg_q303 AND symb_decoder(16#99#)) OR
 					(reg_q303 AND symb_decoder(16#6f#)) OR
 					(reg_q303 AND symb_decoder(16#ed#)) OR
 					(reg_q303 AND symb_decoder(16#2b#)) OR
 					(reg_q303 AND symb_decoder(16#08#)) OR
 					(reg_q303 AND symb_decoder(16#c2#)) OR
 					(reg_q303 AND symb_decoder(16#82#)) OR
 					(reg_q303 AND symb_decoder(16#ea#)) OR
 					(reg_q303 AND symb_decoder(16#25#)) OR
 					(reg_q303 AND symb_decoder(16#09#)) OR
 					(reg_q303 AND symb_decoder(16#57#)) OR
 					(reg_q303 AND symb_decoder(16#64#)) OR
 					(reg_q303 AND symb_decoder(16#10#)) OR
 					(reg_q303 AND symb_decoder(16#db#)) OR
 					(reg_q303 AND symb_decoder(16#fc#)) OR
 					(reg_q303 AND symb_decoder(16#ad#)) OR
 					(reg_q303 AND symb_decoder(16#83#)) OR
 					(reg_q303 AND symb_decoder(16#4f#)) OR
 					(reg_q303 AND symb_decoder(16#14#)) OR
 					(reg_q303 AND symb_decoder(16#66#)) OR
 					(reg_q303 AND symb_decoder(16#7f#)) OR
 					(reg_q303 AND symb_decoder(16#7c#)) OR
 					(reg_q303 AND symb_decoder(16#b3#)) OR
 					(reg_q303 AND symb_decoder(16#94#)) OR
 					(reg_q303 AND symb_decoder(16#8c#)) OR
 					(reg_q303 AND symb_decoder(16#31#)) OR
 					(reg_q303 AND symb_decoder(16#a2#)) OR
 					(reg_q303 AND symb_decoder(16#b8#)) OR
 					(reg_q303 AND symb_decoder(16#52#)) OR
 					(reg_q303 AND symb_decoder(16#e3#)) OR
 					(reg_q303 AND symb_decoder(16#40#)) OR
 					(reg_q303 AND symb_decoder(16#98#)) OR
 					(reg_q303 AND symb_decoder(16#d6#)) OR
 					(reg_q303 AND symb_decoder(16#5f#)) OR
 					(reg_q303 AND symb_decoder(16#f9#)) OR
 					(reg_q303 AND symb_decoder(16#44#)) OR
 					(reg_q303 AND symb_decoder(16#ba#)) OR
 					(reg_q303 AND symb_decoder(16#71#)) OR
 					(reg_q303 AND symb_decoder(16#39#)) OR
 					(reg_q303 AND symb_decoder(16#3e#)) OR
 					(reg_q303 AND symb_decoder(16#28#)) OR
 					(reg_q303 AND symb_decoder(16#b2#)) OR
 					(reg_q303 AND symb_decoder(16#73#)) OR
 					(reg_q303 AND symb_decoder(16#0d#)) OR
 					(reg_q303 AND symb_decoder(16#69#)) OR
 					(reg_q303 AND symb_decoder(16#cd#)) OR
 					(reg_q303 AND symb_decoder(16#a0#)) OR
 					(reg_q303 AND symb_decoder(16#e1#)) OR
 					(reg_q303 AND symb_decoder(16#75#)) OR
 					(reg_q303 AND symb_decoder(16#51#)) OR
 					(reg_q303 AND symb_decoder(16#54#)) OR
 					(reg_q303 AND symb_decoder(16#91#)) OR
 					(reg_q303 AND symb_decoder(16#fa#)) OR
 					(reg_q303 AND symb_decoder(16#e7#)) OR
 					(reg_q303 AND symb_decoder(16#b6#)) OR
 					(reg_q303 AND symb_decoder(16#29#)) OR
 					(reg_q303 AND symb_decoder(16#8a#)) OR
 					(reg_q303 AND symb_decoder(16#b1#)) OR
 					(reg_q303 AND symb_decoder(16#20#)) OR
 					(reg_q303 AND symb_decoder(16#f3#)) OR
 					(reg_q303 AND symb_decoder(16#a8#)) OR
 					(reg_q303 AND symb_decoder(16#1f#)) OR
 					(reg_q303 AND symb_decoder(16#06#)) OR
 					(reg_q303 AND symb_decoder(16#4c#)) OR
 					(reg_q303 AND symb_decoder(16#9e#)) OR
 					(reg_q303 AND symb_decoder(16#42#)) OR
 					(reg_q303 AND symb_decoder(16#48#)) OR
 					(reg_q303 AND symb_decoder(16#80#)) OR
 					(reg_q303 AND symb_decoder(16#a4#)) OR
 					(reg_q303 AND symb_decoder(16#3a#)) OR
 					(reg_q303 AND symb_decoder(16#0e#)) OR
 					(reg_q303 AND symb_decoder(16#a6#)) OR
 					(reg_q303 AND symb_decoder(16#bf#)) OR
 					(reg_q303 AND symb_decoder(16#d4#)) OR
 					(reg_q303 AND symb_decoder(16#4e#)) OR
 					(reg_q303 AND symb_decoder(16#37#)) OR
 					(reg_q303 AND symb_decoder(16#61#)) OR
 					(reg_q303 AND symb_decoder(16#2f#)) OR
 					(reg_q303 AND symb_decoder(16#2c#)) OR
 					(reg_q303 AND symb_decoder(16#ca#)) OR
 					(reg_q303 AND symb_decoder(16#c5#)) OR
 					(reg_q303 AND symb_decoder(16#be#)) OR
 					(reg_q303 AND symb_decoder(16#c8#)) OR
 					(reg_q303 AND symb_decoder(16#b5#)) OR
 					(reg_q303 AND symb_decoder(16#9c#)) OR
 					(reg_q303 AND symb_decoder(16#9a#)) OR
 					(reg_q303 AND symb_decoder(16#aa#)) OR
 					(reg_q303 AND symb_decoder(16#89#)) OR
 					(reg_q303 AND symb_decoder(16#e5#)) OR
 					(reg_q303 AND symb_decoder(16#f0#)) OR
 					(reg_q303 AND symb_decoder(16#e9#)) OR
 					(reg_q303 AND symb_decoder(16#1e#));
reg_q303_init <= '0' ;
	p_reg_q303: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q303 <= reg_q303_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q303 <= reg_q303_init;
        else
          reg_q303 <= reg_q303_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q247_in <= (reg_q245 AND symb_decoder(16#ff#));
reg_q247_init <= '0' ;
	p_reg_q247: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q247 <= reg_q247_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q247 <= reg_q247_init;
        else
          reg_q247 <= reg_q247_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q249_in <= (reg_q247 AND symb_decoder(16#30#)) OR
 					(reg_q247 AND symb_decoder(16#38#)) OR
 					(reg_q247 AND symb_decoder(16#33#)) OR
 					(reg_q247 AND symb_decoder(16#37#)) OR
 					(reg_q247 AND symb_decoder(16#39#)) OR
 					(reg_q247 AND symb_decoder(16#34#)) OR
 					(reg_q247 AND symb_decoder(16#32#)) OR
 					(reg_q247 AND symb_decoder(16#31#)) OR
 					(reg_q247 AND symb_decoder(16#36#)) OR
 					(reg_q247 AND symb_decoder(16#35#)) OR
 					(reg_q249 AND symb_decoder(16#38#)) OR
 					(reg_q249 AND symb_decoder(16#32#)) OR
 					(reg_q249 AND symb_decoder(16#39#)) OR
 					(reg_q249 AND symb_decoder(16#30#)) OR
 					(reg_q249 AND symb_decoder(16#31#)) OR
 					(reg_q249 AND symb_decoder(16#34#)) OR
 					(reg_q249 AND symb_decoder(16#35#)) OR
 					(reg_q249 AND symb_decoder(16#37#)) OR
 					(reg_q249 AND symb_decoder(16#36#)) OR
 					(reg_q249 AND symb_decoder(16#33#));
reg_q249_init <= '0' ;
	p_reg_q249: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q249 <= reg_q249_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q249 <= reg_q249_init;
        else
          reg_q249 <= reg_q249_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2615_in <= (reg_q2615 AND symb_decoder(16#e2#)) OR
 					(reg_q2615 AND symb_decoder(16#1e#)) OR
 					(reg_q2615 AND symb_decoder(16#35#)) OR
 					(reg_q2615 AND symb_decoder(16#cc#)) OR
 					(reg_q2615 AND symb_decoder(16#49#)) OR
 					(reg_q2615 AND symb_decoder(16#2e#)) OR
 					(reg_q2615 AND symb_decoder(16#b4#)) OR
 					(reg_q2615 AND symb_decoder(16#2f#)) OR
 					(reg_q2615 AND symb_decoder(16#41#)) OR
 					(reg_q2615 AND symb_decoder(16#ec#)) OR
 					(reg_q2615 AND symb_decoder(16#16#)) OR
 					(reg_q2615 AND symb_decoder(16#11#)) OR
 					(reg_q2615 AND symb_decoder(16#47#)) OR
 					(reg_q2615 AND symb_decoder(16#9a#)) OR
 					(reg_q2615 AND symb_decoder(16#53#)) OR
 					(reg_q2615 AND symb_decoder(16#ce#)) OR
 					(reg_q2615 AND symb_decoder(16#46#)) OR
 					(reg_q2615 AND symb_decoder(16#de#)) OR
 					(reg_q2615 AND symb_decoder(16#88#)) OR
 					(reg_q2615 AND symb_decoder(16#86#)) OR
 					(reg_q2615 AND symb_decoder(16#f4#)) OR
 					(reg_q2615 AND symb_decoder(16#59#)) OR
 					(reg_q2615 AND symb_decoder(16#d2#)) OR
 					(reg_q2615 AND symb_decoder(16#61#)) OR
 					(reg_q2615 AND symb_decoder(16#cb#)) OR
 					(reg_q2615 AND symb_decoder(16#00#)) OR
 					(reg_q2615 AND symb_decoder(16#3b#)) OR
 					(reg_q2615 AND symb_decoder(16#55#)) OR
 					(reg_q2615 AND symb_decoder(16#b3#)) OR
 					(reg_q2615 AND symb_decoder(16#bb#)) OR
 					(reg_q2615 AND symb_decoder(16#4a#)) OR
 					(reg_q2615 AND symb_decoder(16#0c#)) OR
 					(reg_q2615 AND symb_decoder(16#4e#)) OR
 					(reg_q2615 AND symb_decoder(16#c2#)) OR
 					(reg_q2615 AND symb_decoder(16#3a#)) OR
 					(reg_q2615 AND symb_decoder(16#1c#)) OR
 					(reg_q2615 AND symb_decoder(16#13#)) OR
 					(reg_q2615 AND symb_decoder(16#c6#)) OR
 					(reg_q2615 AND symb_decoder(16#8a#)) OR
 					(reg_q2615 AND symb_decoder(16#91#)) OR
 					(reg_q2615 AND symb_decoder(16#f2#)) OR
 					(reg_q2615 AND symb_decoder(16#12#)) OR
 					(reg_q2615 AND symb_decoder(16#b8#)) OR
 					(reg_q2615 AND symb_decoder(16#a2#)) OR
 					(reg_q2615 AND symb_decoder(16#97#)) OR
 					(reg_q2615 AND symb_decoder(16#1f#)) OR
 					(reg_q2615 AND symb_decoder(16#c9#)) OR
 					(reg_q2615 AND symb_decoder(16#d7#)) OR
 					(reg_q2615 AND symb_decoder(16#d1#)) OR
 					(reg_q2615 AND symb_decoder(16#ff#)) OR
 					(reg_q2615 AND symb_decoder(16#17#)) OR
 					(reg_q2615 AND symb_decoder(16#06#)) OR
 					(reg_q2615 AND symb_decoder(16#51#)) OR
 					(reg_q2615 AND symb_decoder(16#a0#)) OR
 					(reg_q2615 AND symb_decoder(16#e9#)) OR
 					(reg_q2615 AND symb_decoder(16#98#)) OR
 					(reg_q2615 AND symb_decoder(16#33#)) OR
 					(reg_q2615 AND symb_decoder(16#83#)) OR
 					(reg_q2615 AND symb_decoder(16#23#)) OR
 					(reg_q2615 AND symb_decoder(16#94#)) OR
 					(reg_q2615 AND symb_decoder(16#74#)) OR
 					(reg_q2615 AND symb_decoder(16#79#)) OR
 					(reg_q2615 AND symb_decoder(16#8c#)) OR
 					(reg_q2615 AND symb_decoder(16#bf#)) OR
 					(reg_q2615 AND symb_decoder(16#f6#)) OR
 					(reg_q2615 AND symb_decoder(16#7f#)) OR
 					(reg_q2615 AND symb_decoder(16#7a#)) OR
 					(reg_q2615 AND symb_decoder(16#be#)) OR
 					(reg_q2615 AND symb_decoder(16#70#)) OR
 					(reg_q2615 AND symb_decoder(16#6b#)) OR
 					(reg_q2615 AND symb_decoder(16#bd#)) OR
 					(reg_q2615 AND symb_decoder(16#5e#)) OR
 					(reg_q2615 AND symb_decoder(16#73#)) OR
 					(reg_q2615 AND symb_decoder(16#77#)) OR
 					(reg_q2615 AND symb_decoder(16#07#)) OR
 					(reg_q2615 AND symb_decoder(16#6c#)) OR
 					(reg_q2615 AND symb_decoder(16#c3#)) OR
 					(reg_q2615 AND symb_decoder(16#4c#)) OR
 					(reg_q2615 AND symb_decoder(16#1d#)) OR
 					(reg_q2615 AND symb_decoder(16#03#)) OR
 					(reg_q2615 AND symb_decoder(16#ef#)) OR
 					(reg_q2615 AND symb_decoder(16#cd#)) OR
 					(reg_q2615 AND symb_decoder(16#32#)) OR
 					(reg_q2615 AND symb_decoder(16#fd#)) OR
 					(reg_q2615 AND symb_decoder(16#93#)) OR
 					(reg_q2615 AND symb_decoder(16#f9#)) OR
 					(reg_q2615 AND symb_decoder(16#4f#)) OR
 					(reg_q2615 AND symb_decoder(16#f8#)) OR
 					(reg_q2615 AND symb_decoder(16#18#)) OR
 					(reg_q2615 AND symb_decoder(16#df#)) OR
 					(reg_q2615 AND symb_decoder(16#db#)) OR
 					(reg_q2615 AND symb_decoder(16#e4#)) OR
 					(reg_q2615 AND symb_decoder(16#a1#)) OR
 					(reg_q2615 AND symb_decoder(16#37#)) OR
 					(reg_q2615 AND symb_decoder(16#e3#)) OR
 					(reg_q2615 AND symb_decoder(16#9d#)) OR
 					(reg_q2615 AND symb_decoder(16#b5#)) OR
 					(reg_q2615 AND symb_decoder(16#b9#)) OR
 					(reg_q2615 AND symb_decoder(16#5a#)) OR
 					(reg_q2615 AND symb_decoder(16#fb#)) OR
 					(reg_q2615 AND symb_decoder(16#b2#)) OR
 					(reg_q2615 AND symb_decoder(16#99#)) OR
 					(reg_q2615 AND symb_decoder(16#8b#)) OR
 					(reg_q2615 AND symb_decoder(16#39#)) OR
 					(reg_q2615 AND symb_decoder(16#6f#)) OR
 					(reg_q2615 AND symb_decoder(16#b7#)) OR
 					(reg_q2615 AND symb_decoder(16#81#)) OR
 					(reg_q2615 AND symb_decoder(16#80#)) OR
 					(reg_q2615 AND symb_decoder(16#20#)) OR
 					(reg_q2615 AND symb_decoder(16#e7#)) OR
 					(reg_q2615 AND symb_decoder(16#19#)) OR
 					(reg_q2615 AND symb_decoder(16#a4#)) OR
 					(reg_q2615 AND symb_decoder(16#d3#)) OR
 					(reg_q2615 AND symb_decoder(16#a8#)) OR
 					(reg_q2615 AND symb_decoder(16#d0#)) OR
 					(reg_q2615 AND symb_decoder(16#eb#)) OR
 					(reg_q2615 AND symb_decoder(16#72#)) OR
 					(reg_q2615 AND symb_decoder(16#27#)) OR
 					(reg_q2615 AND symb_decoder(16#54#)) OR
 					(reg_q2615 AND symb_decoder(16#2a#)) OR
 					(reg_q2615 AND symb_decoder(16#af#)) OR
 					(reg_q2615 AND symb_decoder(16#42#)) OR
 					(reg_q2615 AND symb_decoder(16#e1#)) OR
 					(reg_q2615 AND symb_decoder(16#6d#)) OR
 					(reg_q2615 AND symb_decoder(16#fc#)) OR
 					(reg_q2615 AND symb_decoder(16#6e#)) OR
 					(reg_q2615 AND symb_decoder(16#57#)) OR
 					(reg_q2615 AND symb_decoder(16#dc#)) OR
 					(reg_q2615 AND symb_decoder(16#a5#)) OR
 					(reg_q2615 AND symb_decoder(16#d9#)) OR
 					(reg_q2615 AND symb_decoder(16#21#)) OR
 					(reg_q2615 AND symb_decoder(16#31#)) OR
 					(reg_q2615 AND symb_decoder(16#22#)) OR
 					(reg_q2615 AND symb_decoder(16#e5#)) OR
 					(reg_q2615 AND symb_decoder(16#9e#)) OR
 					(reg_q2615 AND symb_decoder(16#ed#)) OR
 					(reg_q2615 AND symb_decoder(16#fe#)) OR
 					(reg_q2615 AND symb_decoder(16#85#)) OR
 					(reg_q2615 AND symb_decoder(16#7e#)) OR
 					(reg_q2615 AND symb_decoder(16#08#)) OR
 					(reg_q2615 AND symb_decoder(16#ac#)) OR
 					(reg_q2615 AND symb_decoder(16#5d#)) OR
 					(reg_q2615 AND symb_decoder(16#a6#)) OR
 					(reg_q2615 AND symb_decoder(16#a9#)) OR
 					(reg_q2615 AND symb_decoder(16#d8#)) OR
 					(reg_q2615 AND symb_decoder(16#26#)) OR
 					(reg_q2615 AND symb_decoder(16#e8#)) OR
 					(reg_q2615 AND symb_decoder(16#c8#)) OR
 					(reg_q2615 AND symb_decoder(16#63#)) OR
 					(reg_q2615 AND symb_decoder(16#71#)) OR
 					(reg_q2615 AND symb_decoder(16#9b#)) OR
 					(reg_q2615 AND symb_decoder(16#ae#)) OR
 					(reg_q2615 AND symb_decoder(16#24#)) OR
 					(reg_q2615 AND symb_decoder(16#36#)) OR
 					(reg_q2615 AND symb_decoder(16#05#)) OR
 					(reg_q2615 AND symb_decoder(16#67#)) OR
 					(reg_q2615 AND symb_decoder(16#84#)) OR
 					(reg_q2615 AND symb_decoder(16#1a#)) OR
 					(reg_q2615 AND symb_decoder(16#89#)) OR
 					(reg_q2615 AND symb_decoder(16#92#)) OR
 					(reg_q2615 AND symb_decoder(16#a3#)) OR
 					(reg_q2615 AND symb_decoder(16#45#)) OR
 					(reg_q2615 AND symb_decoder(16#f5#)) OR
 					(reg_q2615 AND symb_decoder(16#29#)) OR
 					(reg_q2615 AND symb_decoder(16#7b#)) OR
 					(reg_q2615 AND symb_decoder(16#3c#)) OR
 					(reg_q2615 AND symb_decoder(16#5c#)) OR
 					(reg_q2615 AND symb_decoder(16#62#)) OR
 					(reg_q2615 AND symb_decoder(16#fa#)) OR
 					(reg_q2615 AND symb_decoder(16#3e#)) OR
 					(reg_q2615 AND symb_decoder(16#90#)) OR
 					(reg_q2615 AND symb_decoder(16#bc#)) OR
 					(reg_q2615 AND symb_decoder(16#f0#)) OR
 					(reg_q2615 AND symb_decoder(16#5f#)) OR
 					(reg_q2615 AND symb_decoder(16#65#)) OR
 					(reg_q2615 AND symb_decoder(16#da#)) OR
 					(reg_q2615 AND symb_decoder(16#f3#)) OR
 					(reg_q2615 AND symb_decoder(16#1b#)) OR
 					(reg_q2615 AND symb_decoder(16#ad#)) OR
 					(reg_q2615 AND symb_decoder(16#0f#)) OR
 					(reg_q2615 AND symb_decoder(16#5b#)) OR
 					(reg_q2615 AND symb_decoder(16#66#)) OR
 					(reg_q2615 AND symb_decoder(16#02#)) OR
 					(reg_q2615 AND symb_decoder(16#ea#)) OR
 					(reg_q2615 AND symb_decoder(16#f7#)) OR
 					(reg_q2615 AND symb_decoder(16#34#)) OR
 					(reg_q2615 AND symb_decoder(16#c0#)) OR
 					(reg_q2615 AND symb_decoder(16#7c#)) OR
 					(reg_q2615 AND symb_decoder(16#3f#)) OR
 					(reg_q2615 AND symb_decoder(16#4d#)) OR
 					(reg_q2615 AND symb_decoder(16#f1#)) OR
 					(reg_q2615 AND symb_decoder(16#30#)) OR
 					(reg_q2615 AND symb_decoder(16#c1#)) OR
 					(reg_q2615 AND symb_decoder(16#b1#)) OR
 					(reg_q2615 AND symb_decoder(16#cf#)) OR
 					(reg_q2615 AND symb_decoder(16#68#)) OR
 					(reg_q2615 AND symb_decoder(16#7d#)) OR
 					(reg_q2615 AND symb_decoder(16#4b#)) OR
 					(reg_q2615 AND symb_decoder(16#10#)) OR
 					(reg_q2615 AND symb_decoder(16#64#)) OR
 					(reg_q2615 AND symb_decoder(16#58#)) OR
 					(reg_q2615 AND symb_decoder(16#8d#)) OR
 					(reg_q2615 AND symb_decoder(16#b6#)) OR
 					(reg_q2615 AND symb_decoder(16#01#)) OR
 					(reg_q2615 AND symb_decoder(16#e0#)) OR
 					(reg_q2615 AND symb_decoder(16#b0#)) OR
 					(reg_q2615 AND symb_decoder(16#d5#)) OR
 					(reg_q2615 AND symb_decoder(16#2b#)) OR
 					(reg_q2615 AND symb_decoder(16#43#)) OR
 					(reg_q2615 AND symb_decoder(16#ca#)) OR
 					(reg_q2615 AND symb_decoder(16#52#)) OR
 					(reg_q2615 AND symb_decoder(16#6a#)) OR
 					(reg_q2615 AND symb_decoder(16#d4#)) OR
 					(reg_q2615 AND symb_decoder(16#04#)) OR
 					(reg_q2615 AND symb_decoder(16#ba#)) OR
 					(reg_q2615 AND symb_decoder(16#3d#)) OR
 					(reg_q2615 AND symb_decoder(16#e6#)) OR
 					(reg_q2615 AND symb_decoder(16#25#)) OR
 					(reg_q2615 AND symb_decoder(16#9c#)) OR
 					(reg_q2615 AND symb_decoder(16#50#)) OR
 					(reg_q2615 AND symb_decoder(16#14#)) OR
 					(reg_q2615 AND symb_decoder(16#56#)) OR
 					(reg_q2615 AND symb_decoder(16#60#)) OR
 					(reg_q2615 AND symb_decoder(16#dd#)) OR
 					(reg_q2615 AND symb_decoder(16#09#)) OR
 					(reg_q2615 AND symb_decoder(16#96#)) OR
 					(reg_q2615 AND symb_decoder(16#c5#)) OR
 					(reg_q2615 AND symb_decoder(16#82#)) OR
 					(reg_q2615 AND symb_decoder(16#38#)) OR
 					(reg_q2615 AND symb_decoder(16#75#)) OR
 					(reg_q2615 AND symb_decoder(16#40#)) OR
 					(reg_q2615 AND symb_decoder(16#a7#)) OR
 					(reg_q2615 AND symb_decoder(16#c4#)) OR
 					(reg_q2615 AND symb_decoder(16#0b#)) OR
 					(reg_q2615 AND symb_decoder(16#15#)) OR
 					(reg_q2615 AND symb_decoder(16#28#)) OR
 					(reg_q2615 AND symb_decoder(16#69#)) OR
 					(reg_q2615 AND symb_decoder(16#9f#)) OR
 					(reg_q2615 AND symb_decoder(16#95#)) OR
 					(reg_q2615 AND symb_decoder(16#2c#)) OR
 					(reg_q2615 AND symb_decoder(16#87#)) OR
 					(reg_q2615 AND symb_decoder(16#ab#)) OR
 					(reg_q2615 AND symb_decoder(16#0e#)) OR
 					(reg_q2615 AND symb_decoder(16#8e#)) OR
 					(reg_q2615 AND symb_decoder(16#c7#)) OR
 					(reg_q2615 AND symb_decoder(16#ee#)) OR
 					(reg_q2615 AND symb_decoder(16#8f#)) OR
 					(reg_q2615 AND symb_decoder(16#78#)) OR
 					(reg_q2615 AND symb_decoder(16#aa#)) OR
 					(reg_q2615 AND symb_decoder(16#d6#)) OR
 					(reg_q2615 AND symb_decoder(16#2d#)) OR
 					(reg_q2615 AND symb_decoder(16#76#)) OR
 					(reg_q2615 AND symb_decoder(16#48#)) OR
 					(reg_q2615 AND symb_decoder(16#44#)) OR
 					(reg_q2579 AND symb_decoder(16#a3#)) OR
 					(reg_q2579 AND symb_decoder(16#ac#)) OR
 					(reg_q2579 AND symb_decoder(16#0b#)) OR
 					(reg_q2579 AND symb_decoder(16#57#)) OR
 					(reg_q2579 AND symb_decoder(16#7c#)) OR
 					(reg_q2579 AND symb_decoder(16#e0#)) OR
 					(reg_q2579 AND symb_decoder(16#9a#)) OR
 					(reg_q2579 AND symb_decoder(16#73#)) OR
 					(reg_q2579 AND symb_decoder(16#99#)) OR
 					(reg_q2579 AND symb_decoder(16#f1#)) OR
 					(reg_q2579 AND symb_decoder(16#c5#)) OR
 					(reg_q2579 AND symb_decoder(16#d5#)) OR
 					(reg_q2579 AND symb_decoder(16#6e#)) OR
 					(reg_q2579 AND symb_decoder(16#03#)) OR
 					(reg_q2579 AND symb_decoder(16#58#)) OR
 					(reg_q2579 AND symb_decoder(16#72#)) OR
 					(reg_q2579 AND symb_decoder(16#01#)) OR
 					(reg_q2579 AND symb_decoder(16#17#)) OR
 					(reg_q2579 AND symb_decoder(16#23#)) OR
 					(reg_q2579 AND symb_decoder(16#95#)) OR
 					(reg_q2579 AND symb_decoder(16#fb#)) OR
 					(reg_q2579 AND symb_decoder(16#a9#)) OR
 					(reg_q2579 AND symb_decoder(16#41#)) OR
 					(reg_q2579 AND symb_decoder(16#dd#)) OR
 					(reg_q2579 AND symb_decoder(16#fc#)) OR
 					(reg_q2579 AND symb_decoder(16#88#)) OR
 					(reg_q2579 AND symb_decoder(16#c7#)) OR
 					(reg_q2579 AND symb_decoder(16#bb#)) OR
 					(reg_q2579 AND symb_decoder(16#5b#)) OR
 					(reg_q2579 AND symb_decoder(16#56#)) OR
 					(reg_q2579 AND symb_decoder(16#e4#)) OR
 					(reg_q2579 AND symb_decoder(16#87#)) OR
 					(reg_q2579 AND symb_decoder(16#35#)) OR
 					(reg_q2579 AND symb_decoder(16#e6#)) OR
 					(reg_q2579 AND symb_decoder(16#1e#)) OR
 					(reg_q2579 AND symb_decoder(16#bd#)) OR
 					(reg_q2579 AND symb_decoder(16#b2#)) OR
 					(reg_q2579 AND symb_decoder(16#de#)) OR
 					(reg_q2579 AND symb_decoder(16#6c#)) OR
 					(reg_q2579 AND symb_decoder(16#42#)) OR
 					(reg_q2579 AND symb_decoder(16#e3#)) OR
 					(reg_q2579 AND symb_decoder(16#20#)) OR
 					(reg_q2579 AND symb_decoder(16#b7#)) OR
 					(reg_q2579 AND symb_decoder(16#90#)) OR
 					(reg_q2579 AND symb_decoder(16#c6#)) OR
 					(reg_q2579 AND symb_decoder(16#c3#)) OR
 					(reg_q2579 AND symb_decoder(16#19#)) OR
 					(reg_q2579 AND symb_decoder(16#ee#)) OR
 					(reg_q2579 AND symb_decoder(16#13#)) OR
 					(reg_q2579 AND symb_decoder(16#9f#)) OR
 					(reg_q2579 AND symb_decoder(16#34#)) OR
 					(reg_q2579 AND symb_decoder(16#68#)) OR
 					(reg_q2579 AND symb_decoder(16#84#)) OR
 					(reg_q2579 AND symb_decoder(16#43#)) OR
 					(reg_q2579 AND symb_decoder(16#91#)) OR
 					(reg_q2579 AND symb_decoder(16#50#)) OR
 					(reg_q2579 AND symb_decoder(16#79#)) OR
 					(reg_q2579 AND symb_decoder(16#aa#)) OR
 					(reg_q2579 AND symb_decoder(16#1f#)) OR
 					(reg_q2579 AND symb_decoder(16#d1#)) OR
 					(reg_q2579 AND symb_decoder(16#1a#)) OR
 					(reg_q2579 AND symb_decoder(16#39#)) OR
 					(reg_q2579 AND symb_decoder(16#18#)) OR
 					(reg_q2579 AND symb_decoder(16#b5#)) OR
 					(reg_q2579 AND symb_decoder(16#00#)) OR
 					(reg_q2579 AND symb_decoder(16#64#)) OR
 					(reg_q2579 AND symb_decoder(16#77#)) OR
 					(reg_q2579 AND symb_decoder(16#2c#)) OR
 					(reg_q2579 AND symb_decoder(16#30#)) OR
 					(reg_q2579 AND symb_decoder(16#b0#)) OR
 					(reg_q2579 AND symb_decoder(16#33#)) OR
 					(reg_q2579 AND symb_decoder(16#ec#)) OR
 					(reg_q2579 AND symb_decoder(16#25#)) OR
 					(reg_q2579 AND symb_decoder(16#b9#)) OR
 					(reg_q2579 AND symb_decoder(16#9b#)) OR
 					(reg_q2579 AND symb_decoder(16#ba#)) OR
 					(reg_q2579 AND symb_decoder(16#2e#)) OR
 					(reg_q2579 AND symb_decoder(16#f6#)) OR
 					(reg_q2579 AND symb_decoder(16#d0#)) OR
 					(reg_q2579 AND symb_decoder(16#92#)) OR
 					(reg_q2579 AND symb_decoder(16#e5#)) OR
 					(reg_q2579 AND symb_decoder(16#7a#)) OR
 					(reg_q2579 AND symb_decoder(16#d8#)) OR
 					(reg_q2579 AND symb_decoder(16#05#)) OR
 					(reg_q2579 AND symb_decoder(16#5e#)) OR
 					(reg_q2579 AND symb_decoder(16#5d#)) OR
 					(reg_q2579 AND symb_decoder(16#a1#)) OR
 					(reg_q2579 AND symb_decoder(16#4c#)) OR
 					(reg_q2579 AND symb_decoder(16#6f#)) OR
 					(reg_q2579 AND symb_decoder(16#0e#)) OR
 					(reg_q2579 AND symb_decoder(16#7b#)) OR
 					(reg_q2579 AND symb_decoder(16#97#)) OR
 					(reg_q2579 AND symb_decoder(16#bc#)) OR
 					(reg_q2579 AND symb_decoder(16#cc#)) OR
 					(reg_q2579 AND symb_decoder(16#85#)) OR
 					(reg_q2579 AND symb_decoder(16#3a#)) OR
 					(reg_q2579 AND symb_decoder(16#53#)) OR
 					(reg_q2579 AND symb_decoder(16#0f#)) OR
 					(reg_q2579 AND symb_decoder(16#1b#)) OR
 					(reg_q2579 AND symb_decoder(16#a5#)) OR
 					(reg_q2579 AND symb_decoder(16#4f#)) OR
 					(reg_q2579 AND symb_decoder(16#11#)) OR
 					(reg_q2579 AND symb_decoder(16#74#)) OR
 					(reg_q2579 AND symb_decoder(16#21#)) OR
 					(reg_q2579 AND symb_decoder(16#93#)) OR
 					(reg_q2579 AND symb_decoder(16#83#)) OR
 					(reg_q2579 AND symb_decoder(16#be#)) OR
 					(reg_q2579 AND symb_decoder(16#8d#)) OR
 					(reg_q2579 AND symb_decoder(16#08#)) OR
 					(reg_q2579 AND symb_decoder(16#da#)) OR
 					(reg_q2579 AND symb_decoder(16#3b#)) OR
 					(reg_q2579 AND symb_decoder(16#c8#)) OR
 					(reg_q2579 AND symb_decoder(16#a0#)) OR
 					(reg_q2579 AND symb_decoder(16#1c#)) OR
 					(reg_q2579 AND symb_decoder(16#98#)) OR
 					(reg_q2579 AND symb_decoder(16#4b#)) OR
 					(reg_q2579 AND symb_decoder(16#96#)) OR
 					(reg_q2579 AND symb_decoder(16#45#)) OR
 					(reg_q2579 AND symb_decoder(16#40#)) OR
 					(reg_q2579 AND symb_decoder(16#c0#)) OR
 					(reg_q2579 AND symb_decoder(16#a6#)) OR
 					(reg_q2579 AND symb_decoder(16#6a#)) OR
 					(reg_q2579 AND symb_decoder(16#2f#)) OR
 					(reg_q2579 AND symb_decoder(16#d2#)) OR
 					(reg_q2579 AND symb_decoder(16#89#)) OR
 					(reg_q2579 AND symb_decoder(16#7e#)) OR
 					(reg_q2579 AND symb_decoder(16#44#)) OR
 					(reg_q2579 AND symb_decoder(16#a2#)) OR
 					(reg_q2579 AND symb_decoder(16#e7#)) OR
 					(reg_q2579 AND symb_decoder(16#df#)) OR
 					(reg_q2579 AND symb_decoder(16#80#)) OR
 					(reg_q2579 AND symb_decoder(16#9c#)) OR
 					(reg_q2579 AND symb_decoder(16#69#)) OR
 					(reg_q2579 AND symb_decoder(16#8b#)) OR
 					(reg_q2579 AND symb_decoder(16#82#)) OR
 					(reg_q2579 AND symb_decoder(16#71#)) OR
 					(reg_q2579 AND symb_decoder(16#14#)) OR
 					(reg_q2579 AND symb_decoder(16#f5#)) OR
 					(reg_q2579 AND symb_decoder(16#d6#)) OR
 					(reg_q2579 AND symb_decoder(16#3f#)) OR
 					(reg_q2579 AND symb_decoder(16#54#)) OR
 					(reg_q2579 AND symb_decoder(16#27#)) OR
 					(reg_q2579 AND symb_decoder(16#ea#)) OR
 					(reg_q2579 AND symb_decoder(16#76#)) OR
 					(reg_q2579 AND symb_decoder(16#09#)) OR
 					(reg_q2579 AND symb_decoder(16#37#)) OR
 					(reg_q2579 AND symb_decoder(16#3c#)) OR
 					(reg_q2579 AND symb_decoder(16#70#)) OR
 					(reg_q2579 AND symb_decoder(16#ca#)) OR
 					(reg_q2579 AND symb_decoder(16#38#)) OR
 					(reg_q2579 AND symb_decoder(16#4d#)) OR
 					(reg_q2579 AND symb_decoder(16#5c#)) OR
 					(reg_q2579 AND symb_decoder(16#1d#)) OR
 					(reg_q2579 AND symb_decoder(16#28#)) OR
 					(reg_q2579 AND symb_decoder(16#2b#)) OR
 					(reg_q2579 AND symb_decoder(16#4e#)) OR
 					(reg_q2579 AND symb_decoder(16#b4#)) OR
 					(reg_q2579 AND symb_decoder(16#fa#)) OR
 					(reg_q2579 AND symb_decoder(16#8c#)) OR
 					(reg_q2579 AND symb_decoder(16#32#)) OR
 					(reg_q2579 AND symb_decoder(16#81#)) OR
 					(reg_q2579 AND symb_decoder(16#2a#)) OR
 					(reg_q2579 AND symb_decoder(16#59#)) OR
 					(reg_q2579 AND symb_decoder(16#8a#)) OR
 					(reg_q2579 AND symb_decoder(16#cd#)) OR
 					(reg_q2579 AND symb_decoder(16#12#)) OR
 					(reg_q2579 AND symb_decoder(16#3d#)) OR
 					(reg_q2579 AND symb_decoder(16#f8#)) OR
 					(reg_q2579 AND symb_decoder(16#02#)) OR
 					(reg_q2579 AND symb_decoder(16#eb#)) OR
 					(reg_q2579 AND symb_decoder(16#d3#)) OR
 					(reg_q2579 AND symb_decoder(16#f7#)) OR
 					(reg_q2579 AND symb_decoder(16#b3#)) OR
 					(reg_q2579 AND symb_decoder(16#ab#)) OR
 					(reg_q2579 AND symb_decoder(16#f0#)) OR
 					(reg_q2579 AND symb_decoder(16#bf#)) OR
 					(reg_q2579 AND symb_decoder(16#e9#)) OR
 					(reg_q2579 AND symb_decoder(16#c1#)) OR
 					(reg_q2579 AND symb_decoder(16#10#)) OR
 					(reg_q2579 AND symb_decoder(16#a4#)) OR
 					(reg_q2579 AND symb_decoder(16#7f#)) OR
 					(reg_q2579 AND symb_decoder(16#b6#)) OR
 					(reg_q2579 AND symb_decoder(16#52#)) OR
 					(reg_q2579 AND symb_decoder(16#cb#)) OR
 					(reg_q2579 AND symb_decoder(16#ae#)) OR
 					(reg_q2579 AND symb_decoder(16#94#)) OR
 					(reg_q2579 AND symb_decoder(16#b1#)) OR
 					(reg_q2579 AND symb_decoder(16#e2#)) OR
 					(reg_q2579 AND symb_decoder(16#55#)) OR
 					(reg_q2579 AND symb_decoder(16#06#)) OR
 					(reg_q2579 AND symb_decoder(16#29#)) OR
 					(reg_q2579 AND symb_decoder(16#4a#)) OR
 					(reg_q2579 AND symb_decoder(16#6b#)) OR
 					(reg_q2579 AND symb_decoder(16#9d#)) OR
 					(reg_q2579 AND symb_decoder(16#a8#)) OR
 					(reg_q2579 AND symb_decoder(16#3e#)) OR
 					(reg_q2579 AND symb_decoder(16#ad#)) OR
 					(reg_q2579 AND symb_decoder(16#65#)) OR
 					(reg_q2579 AND symb_decoder(16#0c#)) OR
 					(reg_q2579 AND symb_decoder(16#fd#)) OR
 					(reg_q2579 AND symb_decoder(16#36#)) OR
 					(reg_q2579 AND symb_decoder(16#f3#)) OR
 					(reg_q2579 AND symb_decoder(16#2d#)) OR
 					(reg_q2579 AND symb_decoder(16#f4#)) OR
 					(reg_q2579 AND symb_decoder(16#f9#)) OR
 					(reg_q2579 AND symb_decoder(16#cf#)) OR
 					(reg_q2579 AND symb_decoder(16#07#)) OR
 					(reg_q2579 AND symb_decoder(16#8f#)) OR
 					(reg_q2579 AND symb_decoder(16#22#)) OR
 					(reg_q2579 AND symb_decoder(16#a7#)) OR
 					(reg_q2579 AND symb_decoder(16#26#)) OR
 					(reg_q2579 AND symb_decoder(16#67#)) OR
 					(reg_q2579 AND symb_decoder(16#24#)) OR
 					(reg_q2579 AND symb_decoder(16#15#)) OR
 					(reg_q2579 AND symb_decoder(16#dc#)) OR
 					(reg_q2579 AND symb_decoder(16#47#)) OR
 					(reg_q2579 AND symb_decoder(16#16#)) OR
 					(reg_q2579 AND symb_decoder(16#51#)) OR
 					(reg_q2579 AND symb_decoder(16#af#)) OR
 					(reg_q2579 AND symb_decoder(16#fe#)) OR
 					(reg_q2579 AND symb_decoder(16#31#)) OR
 					(reg_q2579 AND symb_decoder(16#61#)) OR
 					(reg_q2579 AND symb_decoder(16#66#)) OR
 					(reg_q2579 AND symb_decoder(16#5a#)) OR
 					(reg_q2579 AND symb_decoder(16#49#)) OR
 					(reg_q2579 AND symb_decoder(16#8e#)) OR
 					(reg_q2579 AND symb_decoder(16#63#)) OR
 					(reg_q2579 AND symb_decoder(16#ce#)) OR
 					(reg_q2579 AND symb_decoder(16#9e#)) OR
 					(reg_q2579 AND symb_decoder(16#db#)) OR
 					(reg_q2579 AND symb_decoder(16#04#)) OR
 					(reg_q2579 AND symb_decoder(16#d4#)) OR
 					(reg_q2579 AND symb_decoder(16#e1#)) OR
 					(reg_q2579 AND symb_decoder(16#ef#)) OR
 					(reg_q2579 AND symb_decoder(16#86#)) OR
 					(reg_q2579 AND symb_decoder(16#c2#)) OR
 					(reg_q2579 AND symb_decoder(16#f2#)) OR
 					(reg_q2579 AND symb_decoder(16#46#)) OR
 					(reg_q2579 AND symb_decoder(16#d9#)) OR
 					(reg_q2579 AND symb_decoder(16#6d#)) OR
 					(reg_q2579 AND symb_decoder(16#7d#)) OR
 					(reg_q2579 AND symb_decoder(16#78#)) OR
 					(reg_q2579 AND symb_decoder(16#5f#)) OR
 					(reg_q2579 AND symb_decoder(16#48#)) OR
 					(reg_q2579 AND symb_decoder(16#75#)) OR
 					(reg_q2579 AND symb_decoder(16#e8#)) OR
 					(reg_q2579 AND symb_decoder(16#ed#)) OR
 					(reg_q2579 AND symb_decoder(16#ff#)) OR
 					(reg_q2579 AND symb_decoder(16#60#)) OR
 					(reg_q2579 AND symb_decoder(16#62#)) OR
 					(reg_q2579 AND symb_decoder(16#d7#)) OR
 					(reg_q2579 AND symb_decoder(16#c4#)) OR
 					(reg_q2579 AND symb_decoder(16#c9#)) OR
 					(reg_q2579 AND symb_decoder(16#b8#));
reg_q2615_init <= '0' ;
	p_reg_q2615: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2615 <= reg_q2615_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2615 <= reg_q2615_init;
        else
          reg_q2615 <= reg_q2615_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2518_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2518 AND symb_decoder(16#80#)) OR
 					(reg_q2518 AND symb_decoder(16#92#)) OR
 					(reg_q2518 AND symb_decoder(16#52#)) OR
 					(reg_q2518 AND symb_decoder(16#75#)) OR
 					(reg_q2518 AND symb_decoder(16#28#)) OR
 					(reg_q2518 AND symb_decoder(16#e1#)) OR
 					(reg_q2518 AND symb_decoder(16#54#)) OR
 					(reg_q2518 AND symb_decoder(16#77#)) OR
 					(reg_q2518 AND symb_decoder(16#6d#)) OR
 					(reg_q2518 AND symb_decoder(16#42#)) OR
 					(reg_q2518 AND symb_decoder(16#a3#)) OR
 					(reg_q2518 AND symb_decoder(16#fc#)) OR
 					(reg_q2518 AND symb_decoder(16#88#)) OR
 					(reg_q2518 AND symb_decoder(16#2f#)) OR
 					(reg_q2518 AND symb_decoder(16#b7#)) OR
 					(reg_q2518 AND symb_decoder(16#26#)) OR
 					(reg_q2518 AND symb_decoder(16#7d#)) OR
 					(reg_q2518 AND symb_decoder(16#55#)) OR
 					(reg_q2518 AND symb_decoder(16#9f#)) OR
 					(reg_q2518 AND symb_decoder(16#ec#)) OR
 					(reg_q2518 AND symb_decoder(16#cb#)) OR
 					(reg_q2518 AND symb_decoder(16#39#)) OR
 					(reg_q2518 AND symb_decoder(16#c9#)) OR
 					(reg_q2518 AND symb_decoder(16#d6#)) OR
 					(reg_q2518 AND symb_decoder(16#e2#)) OR
 					(reg_q2518 AND symb_decoder(16#9e#)) OR
 					(reg_q2518 AND symb_decoder(16#bf#)) OR
 					(reg_q2518 AND symb_decoder(16#79#)) OR
 					(reg_q2518 AND symb_decoder(16#8e#)) OR
 					(reg_q2518 AND symb_decoder(16#63#)) OR
 					(reg_q2518 AND symb_decoder(16#1f#)) OR
 					(reg_q2518 AND symb_decoder(16#2e#)) OR
 					(reg_q2518 AND symb_decoder(16#cc#)) OR
 					(reg_q2518 AND symb_decoder(16#3b#)) OR
 					(reg_q2518 AND symb_decoder(16#27#)) OR
 					(reg_q2518 AND symb_decoder(16#12#)) OR
 					(reg_q2518 AND symb_decoder(16#e7#)) OR
 					(reg_q2518 AND symb_decoder(16#f3#)) OR
 					(reg_q2518 AND symb_decoder(16#03#)) OR
 					(reg_q2518 AND symb_decoder(16#db#)) OR
 					(reg_q2518 AND symb_decoder(16#1d#)) OR
 					(reg_q2518 AND symb_decoder(16#b8#)) OR
 					(reg_q2518 AND symb_decoder(16#ab#)) OR
 					(reg_q2518 AND symb_decoder(16#45#)) OR
 					(reg_q2518 AND symb_decoder(16#6c#)) OR
 					(reg_q2518 AND symb_decoder(16#e0#)) OR
 					(reg_q2518 AND symb_decoder(16#1c#)) OR
 					(reg_q2518 AND symb_decoder(16#f0#)) OR
 					(reg_q2518 AND symb_decoder(16#38#)) OR
 					(reg_q2518 AND symb_decoder(16#7a#)) OR
 					(reg_q2518 AND symb_decoder(16#30#)) OR
 					(reg_q2518 AND symb_decoder(16#3e#)) OR
 					(reg_q2518 AND symb_decoder(16#c5#)) OR
 					(reg_q2518 AND symb_decoder(16#d7#)) OR
 					(reg_q2518 AND symb_decoder(16#59#)) OR
 					(reg_q2518 AND symb_decoder(16#06#)) OR
 					(reg_q2518 AND symb_decoder(16#fb#)) OR
 					(reg_q2518 AND symb_decoder(16#eb#)) OR
 					(reg_q2518 AND symb_decoder(16#31#)) OR
 					(reg_q2518 AND symb_decoder(16#af#)) OR
 					(reg_q2518 AND symb_decoder(16#46#)) OR
 					(reg_q2518 AND symb_decoder(16#29#)) OR
 					(reg_q2518 AND symb_decoder(16#47#)) OR
 					(reg_q2518 AND symb_decoder(16#96#)) OR
 					(reg_q2518 AND symb_decoder(16#e5#)) OR
 					(reg_q2518 AND symb_decoder(16#b9#)) OR
 					(reg_q2518 AND symb_decoder(16#d1#)) OR
 					(reg_q2518 AND symb_decoder(16#41#)) OR
 					(reg_q2518 AND symb_decoder(16#fa#)) OR
 					(reg_q2518 AND symb_decoder(16#74#)) OR
 					(reg_q2518 AND symb_decoder(16#f9#)) OR
 					(reg_q2518 AND symb_decoder(16#f1#)) OR
 					(reg_q2518 AND symb_decoder(16#7c#)) OR
 					(reg_q2518 AND symb_decoder(16#be#)) OR
 					(reg_q2518 AND symb_decoder(16#b6#)) OR
 					(reg_q2518 AND symb_decoder(16#f2#)) OR
 					(reg_q2518 AND symb_decoder(16#71#)) OR
 					(reg_q2518 AND symb_decoder(16#d2#)) OR
 					(reg_q2518 AND symb_decoder(16#85#)) OR
 					(reg_q2518 AND symb_decoder(16#ad#)) OR
 					(reg_q2518 AND symb_decoder(16#d4#)) OR
 					(reg_q2518 AND symb_decoder(16#0f#)) OR
 					(reg_q2518 AND symb_decoder(16#e8#)) OR
 					(reg_q2518 AND symb_decoder(16#94#)) OR
 					(reg_q2518 AND symb_decoder(16#a8#)) OR
 					(reg_q2518 AND symb_decoder(16#aa#)) OR
 					(reg_q2518 AND symb_decoder(16#ae#)) OR
 					(reg_q2518 AND symb_decoder(16#10#)) OR
 					(reg_q2518 AND symb_decoder(16#14#)) OR
 					(reg_q2518 AND symb_decoder(16#c1#)) OR
 					(reg_q2518 AND symb_decoder(16#90#)) OR
 					(reg_q2518 AND symb_decoder(16#c4#)) OR
 					(reg_q2518 AND symb_decoder(16#d3#)) OR
 					(reg_q2518 AND symb_decoder(16#6a#)) OR
 					(reg_q2518 AND symb_decoder(16#1b#)) OR
 					(reg_q2518 AND symb_decoder(16#49#)) OR
 					(reg_q2518 AND symb_decoder(16#d8#)) OR
 					(reg_q2518 AND symb_decoder(16#e9#)) OR
 					(reg_q2518 AND symb_decoder(16#cf#)) OR
 					(reg_q2518 AND symb_decoder(16#6b#)) OR
 					(reg_q2518 AND symb_decoder(16#7b#)) OR
 					(reg_q2518 AND symb_decoder(16#1e#)) OR
 					(reg_q2518 AND symb_decoder(16#c8#)) OR
 					(reg_q2518 AND symb_decoder(16#04#)) OR
 					(reg_q2518 AND symb_decoder(16#c2#)) OR
 					(reg_q2518 AND symb_decoder(16#4e#)) OR
 					(reg_q2518 AND symb_decoder(16#6e#)) OR
 					(reg_q2518 AND symb_decoder(16#9b#)) OR
 					(reg_q2518 AND symb_decoder(16#35#)) OR
 					(reg_q2518 AND symb_decoder(16#84#)) OR
 					(reg_q2518 AND symb_decoder(16#b4#)) OR
 					(reg_q2518 AND symb_decoder(16#4c#)) OR
 					(reg_q2518 AND symb_decoder(16#2b#)) OR
 					(reg_q2518 AND symb_decoder(16#72#)) OR
 					(reg_q2518 AND symb_decoder(16#9c#)) OR
 					(reg_q2518 AND symb_decoder(16#82#)) OR
 					(reg_q2518 AND symb_decoder(16#dc#)) OR
 					(reg_q2518 AND symb_decoder(16#3d#)) OR
 					(reg_q2518 AND symb_decoder(16#ce#)) OR
 					(reg_q2518 AND symb_decoder(16#5f#)) OR
 					(reg_q2518 AND symb_decoder(16#76#)) OR
 					(reg_q2518 AND symb_decoder(16#fe#)) OR
 					(reg_q2518 AND symb_decoder(16#60#)) OR
 					(reg_q2518 AND symb_decoder(16#de#)) OR
 					(reg_q2518 AND symb_decoder(16#17#)) OR
 					(reg_q2518 AND symb_decoder(16#c0#)) OR
 					(reg_q2518 AND symb_decoder(16#40#)) OR
 					(reg_q2518 AND symb_decoder(16#da#)) OR
 					(reg_q2518 AND symb_decoder(16#05#)) OR
 					(reg_q2518 AND symb_decoder(16#22#)) OR
 					(reg_q2518 AND symb_decoder(16#56#)) OR
 					(reg_q2518 AND symb_decoder(16#00#)) OR
 					(reg_q2518 AND symb_decoder(16#bb#)) OR
 					(reg_q2518 AND symb_decoder(16#d0#)) OR
 					(reg_q2518 AND symb_decoder(16#a9#)) OR
 					(reg_q2518 AND symb_decoder(16#64#)) OR
 					(reg_q2518 AND symb_decoder(16#b2#)) OR
 					(reg_q2518 AND symb_decoder(16#48#)) OR
 					(reg_q2518 AND symb_decoder(16#8f#)) OR
 					(reg_q2518 AND symb_decoder(16#ee#)) OR
 					(reg_q2518 AND symb_decoder(16#9a#)) OR
 					(reg_q2518 AND symb_decoder(16#dd#)) OR
 					(reg_q2518 AND symb_decoder(16#61#)) OR
 					(reg_q2518 AND symb_decoder(16#97#)) OR
 					(reg_q2518 AND symb_decoder(16#fd#)) OR
 					(reg_q2518 AND symb_decoder(16#1a#)) OR
 					(reg_q2518 AND symb_decoder(16#44#)) OR
 					(reg_q2518 AND symb_decoder(16#95#)) OR
 					(reg_q2518 AND symb_decoder(16#ed#)) OR
 					(reg_q2518 AND symb_decoder(16#81#)) OR
 					(reg_q2518 AND symb_decoder(16#5a#)) OR
 					(reg_q2518 AND symb_decoder(16#b1#)) OR
 					(reg_q2518 AND symb_decoder(16#f7#)) OR
 					(reg_q2518 AND symb_decoder(16#78#)) OR
 					(reg_q2518 AND symb_decoder(16#02#)) OR
 					(reg_q2518 AND symb_decoder(16#24#)) OR
 					(reg_q2518 AND symb_decoder(16#0a#)) OR
 					(reg_q2518 AND symb_decoder(16#18#)) OR
 					(reg_q2518 AND symb_decoder(16#09#)) OR
 					(reg_q2518 AND symb_decoder(16#62#)) OR
 					(reg_q2518 AND symb_decoder(16#2c#)) OR
 					(reg_q2518 AND symb_decoder(16#bc#)) OR
 					(reg_q2518 AND symb_decoder(16#13#)) OR
 					(reg_q2518 AND symb_decoder(16#69#)) OR
 					(reg_q2518 AND symb_decoder(16#3c#)) OR
 					(reg_q2518 AND symb_decoder(16#37#)) OR
 					(reg_q2518 AND symb_decoder(16#32#)) OR
 					(reg_q2518 AND symb_decoder(16#08#)) OR
 					(reg_q2518 AND symb_decoder(16#f8#)) OR
 					(reg_q2518 AND symb_decoder(16#3f#)) OR
 					(reg_q2518 AND symb_decoder(16#21#)) OR
 					(reg_q2518 AND symb_decoder(16#0d#)) OR
 					(reg_q2518 AND symb_decoder(16#2d#)) OR
 					(reg_q2518 AND symb_decoder(16#f4#)) OR
 					(reg_q2518 AND symb_decoder(16#e4#)) OR
 					(reg_q2518 AND symb_decoder(16#50#)) OR
 					(reg_q2518 AND symb_decoder(16#70#)) OR
 					(reg_q2518 AND symb_decoder(16#df#)) OR
 					(reg_q2518 AND symb_decoder(16#87#)) OR
 					(reg_q2518 AND symb_decoder(16#5c#)) OR
 					(reg_q2518 AND symb_decoder(16#e6#)) OR
 					(reg_q2518 AND symb_decoder(16#a7#)) OR
 					(reg_q2518 AND symb_decoder(16#ba#)) OR
 					(reg_q2518 AND symb_decoder(16#6f#)) OR
 					(reg_q2518 AND symb_decoder(16#19#)) OR
 					(reg_q2518 AND symb_decoder(16#11#)) OR
 					(reg_q2518 AND symb_decoder(16#c7#)) OR
 					(reg_q2518 AND symb_decoder(16#4d#)) OR
 					(reg_q2518 AND symb_decoder(16#0c#)) OR
 					(reg_q2518 AND symb_decoder(16#89#)) OR
 					(reg_q2518 AND symb_decoder(16#43#)) OR
 					(reg_q2518 AND symb_decoder(16#0e#)) OR
 					(reg_q2518 AND symb_decoder(16#01#)) OR
 					(reg_q2518 AND symb_decoder(16#93#)) OR
 					(reg_q2518 AND symb_decoder(16#07#)) OR
 					(reg_q2518 AND symb_decoder(16#d9#)) OR
 					(reg_q2518 AND symb_decoder(16#ef#)) OR
 					(reg_q2518 AND symb_decoder(16#e3#)) OR
 					(reg_q2518 AND symb_decoder(16#98#)) OR
 					(reg_q2518 AND symb_decoder(16#53#)) OR
 					(reg_q2518 AND symb_decoder(16#5e#)) OR
 					(reg_q2518 AND symb_decoder(16#68#)) OR
 					(reg_q2518 AND symb_decoder(16#a4#)) OR
 					(reg_q2518 AND symb_decoder(16#34#)) OR
 					(reg_q2518 AND symb_decoder(16#8c#)) OR
 					(reg_q2518 AND symb_decoder(16#67#)) OR
 					(reg_q2518 AND symb_decoder(16#23#)) OR
 					(reg_q2518 AND symb_decoder(16#a1#)) OR
 					(reg_q2518 AND symb_decoder(16#51#)) OR
 					(reg_q2518 AND symb_decoder(16#99#)) OR
 					(reg_q2518 AND symb_decoder(16#66#)) OR
 					(reg_q2518 AND symb_decoder(16#b3#)) OR
 					(reg_q2518 AND symb_decoder(16#ca#)) OR
 					(reg_q2518 AND symb_decoder(16#f5#)) OR
 					(reg_q2518 AND symb_decoder(16#4f#)) OR
 					(reg_q2518 AND symb_decoder(16#83#)) OR
 					(reg_q2518 AND symb_decoder(16#9d#)) OR
 					(reg_q2518 AND symb_decoder(16#73#)) OR
 					(reg_q2518 AND symb_decoder(16#8d#)) OR
 					(reg_q2518 AND symb_decoder(16#4a#)) OR
 					(reg_q2518 AND symb_decoder(16#b0#)) OR
 					(reg_q2518 AND symb_decoder(16#15#)) OR
 					(reg_q2518 AND symb_decoder(16#8b#)) OR
 					(reg_q2518 AND symb_decoder(16#a6#)) OR
 					(reg_q2518 AND symb_decoder(16#5d#)) OR
 					(reg_q2518 AND symb_decoder(16#a5#)) OR
 					(reg_q2518 AND symb_decoder(16#d5#)) OR
 					(reg_q2518 AND symb_decoder(16#16#)) OR
 					(reg_q2518 AND symb_decoder(16#25#)) OR
 					(reg_q2518 AND symb_decoder(16#3a#)) OR
 					(reg_q2518 AND symb_decoder(16#58#)) OR
 					(reg_q2518 AND symb_decoder(16#bd#)) OR
 					(reg_q2518 AND symb_decoder(16#4b#)) OR
 					(reg_q2518 AND symb_decoder(16#ea#)) OR
 					(reg_q2518 AND symb_decoder(16#86#)) OR
 					(reg_q2518 AND symb_decoder(16#91#)) OR
 					(reg_q2518 AND symb_decoder(16#cd#)) OR
 					(reg_q2518 AND symb_decoder(16#33#)) OR
 					(reg_q2518 AND symb_decoder(16#a2#)) OR
 					(reg_q2518 AND symb_decoder(16#f6#)) OR
 					(reg_q2518 AND symb_decoder(16#ff#)) OR
 					(reg_q2518 AND symb_decoder(16#20#)) OR
 					(reg_q2518 AND symb_decoder(16#b5#)) OR
 					(reg_q2518 AND symb_decoder(16#65#)) OR
 					(reg_q2518 AND symb_decoder(16#57#)) OR
 					(reg_q2518 AND symb_decoder(16#7f#)) OR
 					(reg_q2518 AND symb_decoder(16#8a#)) OR
 					(reg_q2518 AND symb_decoder(16#a0#)) OR
 					(reg_q2518 AND symb_decoder(16#c6#)) OR
 					(reg_q2518 AND symb_decoder(16#2a#)) OR
 					(reg_q2518 AND symb_decoder(16#7e#)) OR
 					(reg_q2518 AND symb_decoder(16#5b#)) OR
 					(reg_q2518 AND symb_decoder(16#ac#)) OR
 					(reg_q2518 AND symb_decoder(16#0b#)) OR
 					(reg_q2518 AND symb_decoder(16#c3#)) OR
 					(reg_q2518 AND symb_decoder(16#36#));
reg_q2518_init <= '0' ;
	p_reg_q2518: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2518 <= reg_q2518_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2518 <= reg_q2518_init;
        else
          reg_q2518 <= reg_q2518_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q791_in <= (reg_q789 AND symb_decoder(16#5e#));
reg_q791_init <= '0' ;
	p_reg_q791: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q791 <= reg_q791_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q791 <= reg_q791_init;
        else
          reg_q791 <= reg_q791_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q828_in <= (reg_q826 AND symb_decoder(16#5e#));
reg_q828_init <= '0' ;
	p_reg_q828: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q828 <= reg_q828_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q828 <= reg_q828_init;
        else
          reg_q828 <= reg_q828_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q848_in <= (reg_q828 AND symb_decoder(16#3d#)) OR
 					(reg_q828 AND symb_decoder(16#30#)) OR
 					(reg_q828 AND symb_decoder(16#85#)) OR
 					(reg_q828 AND symb_decoder(16#8a#)) OR
 					(reg_q828 AND symb_decoder(16#e5#)) OR
 					(reg_q828 AND symb_decoder(16#bb#)) OR
 					(reg_q828 AND symb_decoder(16#90#)) OR
 					(reg_q828 AND symb_decoder(16#3e#)) OR
 					(reg_q828 AND symb_decoder(16#c7#)) OR
 					(reg_q828 AND symb_decoder(16#ef#)) OR
 					(reg_q828 AND symb_decoder(16#91#)) OR
 					(reg_q828 AND symb_decoder(16#83#)) OR
 					(reg_q828 AND symb_decoder(16#b2#)) OR
 					(reg_q828 AND symb_decoder(16#5f#)) OR
 					(reg_q828 AND symb_decoder(16#34#)) OR
 					(reg_q828 AND symb_decoder(16#b1#)) OR
 					(reg_q828 AND symb_decoder(16#a9#)) OR
 					(reg_q828 AND symb_decoder(16#4a#)) OR
 					(reg_q828 AND symb_decoder(16#74#)) OR
 					(reg_q828 AND symb_decoder(16#45#)) OR
 					(reg_q828 AND symb_decoder(16#8c#)) OR
 					(reg_q828 AND symb_decoder(16#bd#)) OR
 					(reg_q828 AND symb_decoder(16#15#)) OR
 					(reg_q828 AND symb_decoder(16#59#)) OR
 					(reg_q828 AND symb_decoder(16#5c#)) OR
 					(reg_q828 AND symb_decoder(16#0b#)) OR
 					(reg_q828 AND symb_decoder(16#af#)) OR
 					(reg_q828 AND symb_decoder(16#95#)) OR
 					(reg_q828 AND symb_decoder(16#9f#)) OR
 					(reg_q828 AND symb_decoder(16#23#)) OR
 					(reg_q828 AND symb_decoder(16#1b#)) OR
 					(reg_q828 AND symb_decoder(16#e2#)) OR
 					(reg_q828 AND symb_decoder(16#35#)) OR
 					(reg_q828 AND symb_decoder(16#8e#)) OR
 					(reg_q828 AND symb_decoder(16#aa#)) OR
 					(reg_q828 AND symb_decoder(16#d0#)) OR
 					(reg_q828 AND symb_decoder(16#ec#)) OR
 					(reg_q828 AND symb_decoder(16#c0#)) OR
 					(reg_q828 AND symb_decoder(16#c5#)) OR
 					(reg_q828 AND symb_decoder(16#08#)) OR
 					(reg_q828 AND symb_decoder(16#77#)) OR
 					(reg_q828 AND symb_decoder(16#be#)) OR
 					(reg_q828 AND symb_decoder(16#39#)) OR
 					(reg_q828 AND symb_decoder(16#52#)) OR
 					(reg_q828 AND symb_decoder(16#98#)) OR
 					(reg_q828 AND symb_decoder(16#33#)) OR
 					(reg_q828 AND symb_decoder(16#bc#)) OR
 					(reg_q828 AND symb_decoder(16#71#)) OR
 					(reg_q828 AND symb_decoder(16#54#)) OR
 					(reg_q828 AND symb_decoder(16#37#)) OR
 					(reg_q828 AND symb_decoder(16#94#)) OR
 					(reg_q828 AND symb_decoder(16#97#)) OR
 					(reg_q828 AND symb_decoder(16#a8#)) OR
 					(reg_q828 AND symb_decoder(16#0f#)) OR
 					(reg_q828 AND symb_decoder(16#cf#)) OR
 					(reg_q828 AND symb_decoder(16#40#)) OR
 					(reg_q828 AND symb_decoder(16#c6#)) OR
 					(reg_q828 AND symb_decoder(16#9a#)) OR
 					(reg_q828 AND symb_decoder(16#f2#)) OR
 					(reg_q828 AND symb_decoder(16#eb#)) OR
 					(reg_q828 AND symb_decoder(16#de#)) OR
 					(reg_q828 AND symb_decoder(16#c4#)) OR
 					(reg_q828 AND symb_decoder(16#d9#)) OR
 					(reg_q828 AND symb_decoder(16#86#)) OR
 					(reg_q828 AND symb_decoder(16#f6#)) OR
 					(reg_q828 AND symb_decoder(16#bf#)) OR
 					(reg_q828 AND symb_decoder(16#a7#)) OR
 					(reg_q828 AND symb_decoder(16#2d#)) OR
 					(reg_q828 AND symb_decoder(16#70#)) OR
 					(reg_q828 AND symb_decoder(16#d2#)) OR
 					(reg_q828 AND symb_decoder(16#ac#)) OR
 					(reg_q828 AND symb_decoder(16#e1#)) OR
 					(reg_q828 AND symb_decoder(16#56#)) OR
 					(reg_q828 AND symb_decoder(16#1f#)) OR
 					(reg_q828 AND symb_decoder(16#e6#)) OR
 					(reg_q828 AND symb_decoder(16#41#)) OR
 					(reg_q828 AND symb_decoder(16#7f#)) OR
 					(reg_q828 AND symb_decoder(16#21#)) OR
 					(reg_q828 AND symb_decoder(16#51#)) OR
 					(reg_q828 AND symb_decoder(16#93#)) OR
 					(reg_q828 AND symb_decoder(16#4b#)) OR
 					(reg_q828 AND symb_decoder(16#2a#)) OR
 					(reg_q828 AND symb_decoder(16#5a#)) OR
 					(reg_q828 AND symb_decoder(16#c2#)) OR
 					(reg_q828 AND symb_decoder(16#fe#)) OR
 					(reg_q828 AND symb_decoder(16#3b#)) OR
 					(reg_q828 AND symb_decoder(16#27#)) OR
 					(reg_q828 AND symb_decoder(16#4c#)) OR
 					(reg_q828 AND symb_decoder(16#f3#)) OR
 					(reg_q828 AND symb_decoder(16#76#)) OR
 					(reg_q828 AND symb_decoder(16#7c#)) OR
 					(reg_q828 AND symb_decoder(16#31#)) OR
 					(reg_q828 AND symb_decoder(16#3c#)) OR
 					(reg_q828 AND symb_decoder(16#cb#)) OR
 					(reg_q828 AND symb_decoder(16#a1#)) OR
 					(reg_q828 AND symb_decoder(16#e9#)) OR
 					(reg_q828 AND symb_decoder(16#c3#)) OR
 					(reg_q828 AND symb_decoder(16#f7#)) OR
 					(reg_q828 AND symb_decoder(16#2f#)) OR
 					(reg_q828 AND symb_decoder(16#1d#)) OR
 					(reg_q828 AND symb_decoder(16#18#)) OR
 					(reg_q828 AND symb_decoder(16#ce#)) OR
 					(reg_q828 AND symb_decoder(16#36#)) OR
 					(reg_q828 AND symb_decoder(16#5e#)) OR
 					(reg_q828 AND symb_decoder(16#38#)) OR
 					(reg_q828 AND symb_decoder(16#61#)) OR
 					(reg_q828 AND symb_decoder(16#e8#)) OR
 					(reg_q828 AND symb_decoder(16#22#)) OR
 					(reg_q828 AND symb_decoder(16#b9#)) OR
 					(reg_q828 AND symb_decoder(16#89#)) OR
 					(reg_q828 AND symb_decoder(16#88#)) OR
 					(reg_q828 AND symb_decoder(16#c9#)) OR
 					(reg_q828 AND symb_decoder(16#25#)) OR
 					(reg_q828 AND symb_decoder(16#0e#)) OR
 					(reg_q828 AND symb_decoder(16#d6#)) OR
 					(reg_q828 AND symb_decoder(16#1c#)) OR
 					(reg_q828 AND symb_decoder(16#b6#)) OR
 					(reg_q828 AND symb_decoder(16#6f#)) OR
 					(reg_q828 AND symb_decoder(16#db#)) OR
 					(reg_q828 AND symb_decoder(16#96#)) OR
 					(reg_q828 AND symb_decoder(16#20#)) OR
 					(reg_q828 AND symb_decoder(16#6d#)) OR
 					(reg_q828 AND symb_decoder(16#fb#)) OR
 					(reg_q828 AND symb_decoder(16#49#)) OR
 					(reg_q828 AND symb_decoder(16#02#)) OR
 					(reg_q828 AND symb_decoder(16#a6#)) OR
 					(reg_q828 AND symb_decoder(16#04#)) OR
 					(reg_q828 AND symb_decoder(16#d1#)) OR
 					(reg_q828 AND symb_decoder(16#32#)) OR
 					(reg_q828 AND symb_decoder(16#9e#)) OR
 					(reg_q828 AND symb_decoder(16#78#)) OR
 					(reg_q828 AND symb_decoder(16#65#)) OR
 					(reg_q828 AND symb_decoder(16#64#)) OR
 					(reg_q828 AND symb_decoder(16#12#)) OR
 					(reg_q828 AND symb_decoder(16#5b#)) OR
 					(reg_q828 AND symb_decoder(16#ee#)) OR
 					(reg_q828 AND symb_decoder(16#df#)) OR
 					(reg_q828 AND symb_decoder(16#05#)) OR
 					(reg_q828 AND symb_decoder(16#58#)) OR
 					(reg_q828 AND symb_decoder(16#69#)) OR
 					(reg_q828 AND symb_decoder(16#ae#)) OR
 					(reg_q828 AND symb_decoder(16#6b#)) OR
 					(reg_q828 AND symb_decoder(16#68#)) OR
 					(reg_q828 AND symb_decoder(16#d4#)) OR
 					(reg_q828 AND symb_decoder(16#13#)) OR
 					(reg_q828 AND symb_decoder(16#28#)) OR
 					(reg_q828 AND symb_decoder(16#dc#)) OR
 					(reg_q828 AND symb_decoder(16#55#)) OR
 					(reg_q828 AND symb_decoder(16#43#)) OR
 					(reg_q828 AND symb_decoder(16#01#)) OR
 					(reg_q828 AND symb_decoder(16#16#)) OR
 					(reg_q828 AND symb_decoder(16#b4#)) OR
 					(reg_q828 AND symb_decoder(16#f5#)) OR
 					(reg_q828 AND symb_decoder(16#b0#)) OR
 					(reg_q828 AND symb_decoder(16#3a#)) OR
 					(reg_q828 AND symb_decoder(16#a4#)) OR
 					(reg_q828 AND symb_decoder(16#4d#)) OR
 					(reg_q828 AND symb_decoder(16#80#)) OR
 					(reg_q828 AND symb_decoder(16#d3#)) OR
 					(reg_q828 AND symb_decoder(16#3f#)) OR
 					(reg_q828 AND symb_decoder(16#2b#)) OR
 					(reg_q828 AND symb_decoder(16#7d#)) OR
 					(reg_q828 AND symb_decoder(16#fd#)) OR
 					(reg_q828 AND symb_decoder(16#75#)) OR
 					(reg_q828 AND symb_decoder(16#42#)) OR
 					(reg_q828 AND symb_decoder(16#8f#)) OR
 					(reg_q828 AND symb_decoder(16#f8#)) OR
 					(reg_q828 AND symb_decoder(16#82#)) OR
 					(reg_q828 AND symb_decoder(16#f9#)) OR
 					(reg_q828 AND symb_decoder(16#cd#)) OR
 					(reg_q828 AND symb_decoder(16#7b#)) OR
 					(reg_q828 AND symb_decoder(16#ba#)) OR
 					(reg_q828 AND symb_decoder(16#d8#)) OR
 					(reg_q828 AND symb_decoder(16#e0#)) OR
 					(reg_q828 AND symb_decoder(16#4e#)) OR
 					(reg_q828 AND symb_decoder(16#a0#)) OR
 					(reg_q828 AND symb_decoder(16#ad#)) OR
 					(reg_q828 AND symb_decoder(16#14#)) OR
 					(reg_q828 AND symb_decoder(16#03#)) OR
 					(reg_q828 AND symb_decoder(16#24#)) OR
 					(reg_q828 AND symb_decoder(16#c8#)) OR
 					(reg_q828 AND symb_decoder(16#2c#)) OR
 					(reg_q828 AND symb_decoder(16#e3#)) OR
 					(reg_q828 AND symb_decoder(16#f4#)) OR
 					(reg_q828 AND symb_decoder(16#72#)) OR
 					(reg_q828 AND symb_decoder(16#b8#)) OR
 					(reg_q828 AND symb_decoder(16#0c#)) OR
 					(reg_q828 AND symb_decoder(16#63#)) OR
 					(reg_q828 AND symb_decoder(16#66#)) OR
 					(reg_q828 AND symb_decoder(16#d7#)) OR
 					(reg_q828 AND symb_decoder(16#e4#)) OR
 					(reg_q828 AND symb_decoder(16#b3#)) OR
 					(reg_q828 AND symb_decoder(16#4f#)) OR
 					(reg_q828 AND symb_decoder(16#19#)) OR
 					(reg_q828 AND symb_decoder(16#6c#)) OR
 					(reg_q828 AND symb_decoder(16#ed#)) OR
 					(reg_q828 AND symb_decoder(16#9d#)) OR
 					(reg_q828 AND symb_decoder(16#b5#)) OR
 					(reg_q828 AND symb_decoder(16#67#)) OR
 					(reg_q828 AND symb_decoder(16#da#)) OR
 					(reg_q828 AND symb_decoder(16#48#)) OR
 					(reg_q828 AND symb_decoder(16#e7#)) OR
 					(reg_q828 AND symb_decoder(16#ca#)) OR
 					(reg_q828 AND symb_decoder(16#ab#)) OR
 					(reg_q828 AND symb_decoder(16#fa#)) OR
 					(reg_q828 AND symb_decoder(16#cc#)) OR
 					(reg_q828 AND symb_decoder(16#62#)) OR
 					(reg_q828 AND symb_decoder(16#99#)) OR
 					(reg_q828 AND symb_decoder(16#9b#)) OR
 					(reg_q828 AND symb_decoder(16#73#)) OR
 					(reg_q828 AND symb_decoder(16#07#)) OR
 					(reg_q828 AND symb_decoder(16#a5#)) OR
 					(reg_q828 AND symb_decoder(16#09#)) OR
 					(reg_q828 AND symb_decoder(16#10#)) OR
 					(reg_q828 AND symb_decoder(16#a2#)) OR
 					(reg_q828 AND symb_decoder(16#ff#)) OR
 					(reg_q828 AND symb_decoder(16#44#)) OR
 					(reg_q828 AND symb_decoder(16#6a#)) OR
 					(reg_q828 AND symb_decoder(16#60#)) OR
 					(reg_q828 AND symb_decoder(16#29#)) OR
 					(reg_q828 AND symb_decoder(16#00#)) OR
 					(reg_q828 AND symb_decoder(16#47#)) OR
 					(reg_q828 AND symb_decoder(16#8b#)) OR
 					(reg_q828 AND symb_decoder(16#7e#)) OR
 					(reg_q828 AND symb_decoder(16#2e#)) OR
 					(reg_q828 AND symb_decoder(16#92#)) OR
 					(reg_q828 AND symb_decoder(16#06#)) OR
 					(reg_q828 AND symb_decoder(16#fc#)) OR
 					(reg_q828 AND symb_decoder(16#6e#)) OR
 					(reg_q828 AND symb_decoder(16#5d#)) OR
 					(reg_q828 AND symb_decoder(16#11#)) OR
 					(reg_q828 AND symb_decoder(16#81#)) OR
 					(reg_q828 AND symb_decoder(16#7a#)) OR
 					(reg_q828 AND symb_decoder(16#f0#)) OR
 					(reg_q828 AND symb_decoder(16#57#)) OR
 					(reg_q828 AND symb_decoder(16#dd#)) OR
 					(reg_q828 AND symb_decoder(16#79#)) OR
 					(reg_q828 AND symb_decoder(16#46#)) OR
 					(reg_q828 AND symb_decoder(16#8d#)) OR
 					(reg_q828 AND symb_decoder(16#a3#)) OR
 					(reg_q828 AND symb_decoder(16#84#)) OR
 					(reg_q828 AND symb_decoder(16#b7#)) OR
 					(reg_q828 AND symb_decoder(16#c1#)) OR
 					(reg_q828 AND symb_decoder(16#d5#)) OR
 					(reg_q828 AND symb_decoder(16#9c#)) OR
 					(reg_q828 AND symb_decoder(16#f1#)) OR
 					(reg_q828 AND symb_decoder(16#53#)) OR
 					(reg_q828 AND symb_decoder(16#26#)) OR
 					(reg_q828 AND symb_decoder(16#ea#)) OR
 					(reg_q828 AND symb_decoder(16#17#)) OR
 					(reg_q828 AND symb_decoder(16#1a#)) OR
 					(reg_q828 AND symb_decoder(16#87#)) OR
 					(reg_q828 AND symb_decoder(16#1e#)) OR
 					(reg_q828 AND symb_decoder(16#50#)) OR
 					(reg_q848 AND symb_decoder(16#ac#)) OR
 					(reg_q848 AND symb_decoder(16#77#)) OR
 					(reg_q848 AND symb_decoder(16#27#)) OR
 					(reg_q848 AND symb_decoder(16#cf#)) OR
 					(reg_q848 AND symb_decoder(16#c3#)) OR
 					(reg_q848 AND symb_decoder(16#43#)) OR
 					(reg_q848 AND symb_decoder(16#49#)) OR
 					(reg_q848 AND symb_decoder(16#42#)) OR
 					(reg_q848 AND symb_decoder(16#b4#)) OR
 					(reg_q848 AND symb_decoder(16#d5#)) OR
 					(reg_q848 AND symb_decoder(16#95#)) OR
 					(reg_q848 AND symb_decoder(16#dd#)) OR
 					(reg_q848 AND symb_decoder(16#61#)) OR
 					(reg_q848 AND symb_decoder(16#a7#)) OR
 					(reg_q848 AND symb_decoder(16#ce#)) OR
 					(reg_q848 AND symb_decoder(16#b5#)) OR
 					(reg_q848 AND symb_decoder(16#2b#)) OR
 					(reg_q848 AND symb_decoder(16#7e#)) OR
 					(reg_q848 AND symb_decoder(16#90#)) OR
 					(reg_q848 AND symb_decoder(16#3e#)) OR
 					(reg_q848 AND symb_decoder(16#a4#)) OR
 					(reg_q848 AND symb_decoder(16#d2#)) OR
 					(reg_q848 AND symb_decoder(16#bd#)) OR
 					(reg_q848 AND symb_decoder(16#28#)) OR
 					(reg_q848 AND symb_decoder(16#aa#)) OR
 					(reg_q848 AND symb_decoder(16#c1#)) OR
 					(reg_q848 AND symb_decoder(16#86#)) OR
 					(reg_q848 AND symb_decoder(16#b1#)) OR
 					(reg_q848 AND symb_decoder(16#fc#)) OR
 					(reg_q848 AND symb_decoder(16#d1#)) OR
 					(reg_q848 AND symb_decoder(16#38#)) OR
 					(reg_q848 AND symb_decoder(16#4c#)) OR
 					(reg_q848 AND symb_decoder(16#5f#)) OR
 					(reg_q848 AND symb_decoder(16#26#)) OR
 					(reg_q848 AND symb_decoder(16#35#)) OR
 					(reg_q848 AND symb_decoder(16#19#)) OR
 					(reg_q848 AND symb_decoder(16#8e#)) OR
 					(reg_q848 AND symb_decoder(16#81#)) OR
 					(reg_q848 AND symb_decoder(16#6e#)) OR
 					(reg_q848 AND symb_decoder(16#2e#)) OR
 					(reg_q848 AND symb_decoder(16#17#)) OR
 					(reg_q848 AND symb_decoder(16#7b#)) OR
 					(reg_q848 AND symb_decoder(16#55#)) OR
 					(reg_q848 AND symb_decoder(16#c4#)) OR
 					(reg_q848 AND symb_decoder(16#70#)) OR
 					(reg_q848 AND symb_decoder(16#f7#)) OR
 					(reg_q848 AND symb_decoder(16#32#)) OR
 					(reg_q848 AND symb_decoder(16#c7#)) OR
 					(reg_q848 AND symb_decoder(16#bc#)) OR
 					(reg_q848 AND symb_decoder(16#df#)) OR
 					(reg_q848 AND symb_decoder(16#5a#)) OR
 					(reg_q848 AND symb_decoder(16#ad#)) OR
 					(reg_q848 AND symb_decoder(16#30#)) OR
 					(reg_q848 AND symb_decoder(16#c0#)) OR
 					(reg_q848 AND symb_decoder(16#d9#)) OR
 					(reg_q848 AND symb_decoder(16#b8#)) OR
 					(reg_q848 AND symb_decoder(16#1d#)) OR
 					(reg_q848 AND symb_decoder(16#2a#)) OR
 					(reg_q848 AND symb_decoder(16#24#)) OR
 					(reg_q848 AND symb_decoder(16#a8#)) OR
 					(reg_q848 AND symb_decoder(16#f6#)) OR
 					(reg_q848 AND symb_decoder(16#58#)) OR
 					(reg_q848 AND symb_decoder(16#3f#)) OR
 					(reg_q848 AND symb_decoder(16#72#)) OR
 					(reg_q848 AND symb_decoder(16#c5#)) OR
 					(reg_q848 AND symb_decoder(16#7c#)) OR
 					(reg_q848 AND symb_decoder(16#bb#)) OR
 					(reg_q848 AND symb_decoder(16#34#)) OR
 					(reg_q848 AND symb_decoder(16#fb#)) OR
 					(reg_q848 AND symb_decoder(16#5e#)) OR
 					(reg_q848 AND symb_decoder(16#b7#)) OR
 					(reg_q848 AND symb_decoder(16#53#)) OR
 					(reg_q848 AND symb_decoder(16#0c#)) OR
 					(reg_q848 AND symb_decoder(16#5b#)) OR
 					(reg_q848 AND symb_decoder(16#2f#)) OR
 					(reg_q848 AND symb_decoder(16#87#)) OR
 					(reg_q848 AND symb_decoder(16#0f#)) OR
 					(reg_q848 AND symb_decoder(16#e5#)) OR
 					(reg_q848 AND symb_decoder(16#4a#)) OR
 					(reg_q848 AND symb_decoder(16#cb#)) OR
 					(reg_q848 AND symb_decoder(16#85#)) OR
 					(reg_q848 AND symb_decoder(16#5c#)) OR
 					(reg_q848 AND symb_decoder(16#1f#)) OR
 					(reg_q848 AND symb_decoder(16#a9#)) OR
 					(reg_q848 AND symb_decoder(16#51#)) OR
 					(reg_q848 AND symb_decoder(16#23#)) OR
 					(reg_q848 AND symb_decoder(16#06#)) OR
 					(reg_q848 AND symb_decoder(16#fe#)) OR
 					(reg_q848 AND symb_decoder(16#8f#)) OR
 					(reg_q848 AND symb_decoder(16#08#)) OR
 					(reg_q848 AND symb_decoder(16#02#)) OR
 					(reg_q848 AND symb_decoder(16#62#)) OR
 					(reg_q848 AND symb_decoder(16#33#)) OR
 					(reg_q848 AND symb_decoder(16#66#)) OR
 					(reg_q848 AND symb_decoder(16#59#)) OR
 					(reg_q848 AND symb_decoder(16#1c#)) OR
 					(reg_q848 AND symb_decoder(16#76#)) OR
 					(reg_q848 AND symb_decoder(16#c6#)) OR
 					(reg_q848 AND symb_decoder(16#71#)) OR
 					(reg_q848 AND symb_decoder(16#56#)) OR
 					(reg_q848 AND symb_decoder(16#04#)) OR
 					(reg_q848 AND symb_decoder(16#e6#)) OR
 					(reg_q848 AND symb_decoder(16#ff#)) OR
 					(reg_q848 AND symb_decoder(16#11#)) OR
 					(reg_q848 AND symb_decoder(16#c8#)) OR
 					(reg_q848 AND symb_decoder(16#ca#)) OR
 					(reg_q848 AND symb_decoder(16#6a#)) OR
 					(reg_q848 AND symb_decoder(16#68#)) OR
 					(reg_q848 AND symb_decoder(16#de#)) OR
 					(reg_q848 AND symb_decoder(16#82#)) OR
 					(reg_q848 AND symb_decoder(16#f3#)) OR
 					(reg_q848 AND symb_decoder(16#13#)) OR
 					(reg_q848 AND symb_decoder(16#a0#)) OR
 					(reg_q848 AND symb_decoder(16#97#)) OR
 					(reg_q848 AND symb_decoder(16#a3#)) OR
 					(reg_q848 AND symb_decoder(16#a6#)) OR
 					(reg_q848 AND symb_decoder(16#73#)) OR
 					(reg_q848 AND symb_decoder(16#40#)) OR
 					(reg_q848 AND symb_decoder(16#b3#)) OR
 					(reg_q848 AND symb_decoder(16#1e#)) OR
 					(reg_q848 AND symb_decoder(16#cd#)) OR
 					(reg_q848 AND symb_decoder(16#e1#)) OR
 					(reg_q848 AND symb_decoder(16#ab#)) OR
 					(reg_q848 AND symb_decoder(16#25#)) OR
 					(reg_q848 AND symb_decoder(16#b0#)) OR
 					(reg_q848 AND symb_decoder(16#89#)) OR
 					(reg_q848 AND symb_decoder(16#9a#)) OR
 					(reg_q848 AND symb_decoder(16#99#)) OR
 					(reg_q848 AND symb_decoder(16#7d#)) OR
 					(reg_q848 AND symb_decoder(16#6b#)) OR
 					(reg_q848 AND symb_decoder(16#9b#)) OR
 					(reg_q848 AND symb_decoder(16#47#)) OR
 					(reg_q848 AND symb_decoder(16#3a#)) OR
 					(reg_q848 AND symb_decoder(16#0e#)) OR
 					(reg_q848 AND symb_decoder(16#48#)) OR
 					(reg_q848 AND symb_decoder(16#41#)) OR
 					(reg_q848 AND symb_decoder(16#af#)) OR
 					(reg_q848 AND symb_decoder(16#84#)) OR
 					(reg_q848 AND symb_decoder(16#1a#)) OR
 					(reg_q848 AND symb_decoder(16#dc#)) OR
 					(reg_q848 AND symb_decoder(16#f0#)) OR
 					(reg_q848 AND symb_decoder(16#8d#)) OR
 					(reg_q848 AND symb_decoder(16#10#)) OR
 					(reg_q848 AND symb_decoder(16#93#)) OR
 					(reg_q848 AND symb_decoder(16#31#)) OR
 					(reg_q848 AND symb_decoder(16#ed#)) OR
 					(reg_q848 AND symb_decoder(16#83#)) OR
 					(reg_q848 AND symb_decoder(16#21#)) OR
 					(reg_q848 AND symb_decoder(16#94#)) OR
 					(reg_q848 AND symb_decoder(16#ae#)) OR
 					(reg_q848 AND symb_decoder(16#f4#)) OR
 					(reg_q848 AND symb_decoder(16#e4#)) OR
 					(reg_q848 AND symb_decoder(16#36#)) OR
 					(reg_q848 AND symb_decoder(16#4e#)) OR
 					(reg_q848 AND symb_decoder(16#52#)) OR
 					(reg_q848 AND symb_decoder(16#f2#)) OR
 					(reg_q848 AND symb_decoder(16#4d#)) OR
 					(reg_q848 AND symb_decoder(16#7a#)) OR
 					(reg_q848 AND symb_decoder(16#6d#)) OR
 					(reg_q848 AND symb_decoder(16#20#)) OR
 					(reg_q848 AND symb_decoder(16#60#)) OR
 					(reg_q848 AND symb_decoder(16#b9#)) OR
 					(reg_q848 AND symb_decoder(16#d0#)) OR
 					(reg_q848 AND symb_decoder(16#fd#)) OR
 					(reg_q848 AND symb_decoder(16#e0#)) OR
 					(reg_q848 AND symb_decoder(16#6c#)) OR
 					(reg_q848 AND symb_decoder(16#3d#)) OR
 					(reg_q848 AND symb_decoder(16#eb#)) OR
 					(reg_q848 AND symb_decoder(16#f5#)) OR
 					(reg_q848 AND symb_decoder(16#a2#)) OR
 					(reg_q848 AND symb_decoder(16#c9#)) OR
 					(reg_q848 AND symb_decoder(16#f8#)) OR
 					(reg_q848 AND symb_decoder(16#ec#)) OR
 					(reg_q848 AND symb_decoder(16#f9#)) OR
 					(reg_q848 AND symb_decoder(16#e2#)) OR
 					(reg_q848 AND symb_decoder(16#8b#)) OR
 					(reg_q848 AND symb_decoder(16#80#)) OR
 					(reg_q848 AND symb_decoder(16#5d#)) OR
 					(reg_q848 AND symb_decoder(16#75#)) OR
 					(reg_q848 AND symb_decoder(16#45#)) OR
 					(reg_q848 AND symb_decoder(16#9d#)) OR
 					(reg_q848 AND symb_decoder(16#39#)) OR
 					(reg_q848 AND symb_decoder(16#8a#)) OR
 					(reg_q848 AND symb_decoder(16#e9#)) OR
 					(reg_q848 AND symb_decoder(16#22#)) OR
 					(reg_q848 AND symb_decoder(16#54#)) OR
 					(reg_q848 AND symb_decoder(16#8c#)) OR
 					(reg_q848 AND symb_decoder(16#78#)) OR
 					(reg_q848 AND symb_decoder(16#79#)) OR
 					(reg_q848 AND symb_decoder(16#15#)) OR
 					(reg_q848 AND symb_decoder(16#09#)) OR
 					(reg_q848 AND symb_decoder(16#6f#)) OR
 					(reg_q848 AND symb_decoder(16#fa#)) OR
 					(reg_q848 AND symb_decoder(16#ef#)) OR
 					(reg_q848 AND symb_decoder(16#cc#)) OR
 					(reg_q848 AND symb_decoder(16#67#)) OR
 					(reg_q848 AND symb_decoder(16#c2#)) OR
 					(reg_q848 AND symb_decoder(16#16#)) OR
 					(reg_q848 AND symb_decoder(16#4b#)) OR
 					(reg_q848 AND symb_decoder(16#05#)) OR
 					(reg_q848 AND symb_decoder(16#e8#)) OR
 					(reg_q848 AND symb_decoder(16#1b#)) OR
 					(reg_q848 AND symb_decoder(16#96#)) OR
 					(reg_q848 AND symb_decoder(16#46#)) OR
 					(reg_q848 AND symb_decoder(16#44#)) OR
 					(reg_q848 AND symb_decoder(16#18#)) OR
 					(reg_q848 AND symb_decoder(16#9c#)) OR
 					(reg_q848 AND symb_decoder(16#69#)) OR
 					(reg_q848 AND symb_decoder(16#07#)) OR
 					(reg_q848 AND symb_decoder(16#7f#)) OR
 					(reg_q848 AND symb_decoder(16#01#)) OR
 					(reg_q848 AND symb_decoder(16#03#)) OR
 					(reg_q848 AND symb_decoder(16#a1#)) OR
 					(reg_q848 AND symb_decoder(16#88#)) OR
 					(reg_q848 AND symb_decoder(16#ee#)) OR
 					(reg_q848 AND symb_decoder(16#74#)) OR
 					(reg_q848 AND symb_decoder(16#9f#)) OR
 					(reg_q848 AND symb_decoder(16#12#)) OR
 					(reg_q848 AND symb_decoder(16#57#)) OR
 					(reg_q848 AND symb_decoder(16#37#)) OR
 					(reg_q848 AND symb_decoder(16#63#)) OR
 					(reg_q848 AND symb_decoder(16#92#)) OR
 					(reg_q848 AND symb_decoder(16#d6#)) OR
 					(reg_q848 AND symb_decoder(16#0b#)) OR
 					(reg_q848 AND symb_decoder(16#29#)) OR
 					(reg_q848 AND symb_decoder(16#50#)) OR
 					(reg_q848 AND symb_decoder(16#64#)) OR
 					(reg_q848 AND symb_decoder(16#2c#)) OR
 					(reg_q848 AND symb_decoder(16#4f#)) OR
 					(reg_q848 AND symb_decoder(16#f1#)) OR
 					(reg_q848 AND symb_decoder(16#9e#)) OR
 					(reg_q848 AND symb_decoder(16#b2#)) OR
 					(reg_q848 AND symb_decoder(16#65#)) OR
 					(reg_q848 AND symb_decoder(16#3c#)) OR
 					(reg_q848 AND symb_decoder(16#2d#)) OR
 					(reg_q848 AND symb_decoder(16#d7#)) OR
 					(reg_q848 AND symb_decoder(16#bf#)) OR
 					(reg_q848 AND symb_decoder(16#e3#)) OR
 					(reg_q848 AND symb_decoder(16#91#)) OR
 					(reg_q848 AND symb_decoder(16#98#)) OR
 					(reg_q848 AND symb_decoder(16#e7#)) OR
 					(reg_q848 AND symb_decoder(16#b6#)) OR
 					(reg_q848 AND symb_decoder(16#d4#)) OR
 					(reg_q848 AND symb_decoder(16#d8#)) OR
 					(reg_q848 AND symb_decoder(16#ba#)) OR
 					(reg_q848 AND symb_decoder(16#14#)) OR
 					(reg_q848 AND symb_decoder(16#a5#)) OR
 					(reg_q848 AND symb_decoder(16#be#)) OR
 					(reg_q848 AND symb_decoder(16#00#)) OR
 					(reg_q848 AND symb_decoder(16#d3#)) OR
 					(reg_q848 AND symb_decoder(16#3b#)) OR
 					(reg_q848 AND symb_decoder(16#ea#)) OR
 					(reg_q848 AND symb_decoder(16#da#)) OR
 					(reg_q848 AND symb_decoder(16#db#));
reg_q848_init <= '0' ;
	p_reg_q848: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q848 <= reg_q848_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q848 <= reg_q848_init;
        else
          reg_q848 <= reg_q848_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q119_in <= (reg_q119 AND symb_decoder(16#09#)) OR
 					(reg_q119 AND symb_decoder(16#20#)) OR
 					(reg_q119 AND symb_decoder(16#0a#)) OR
 					(reg_q119 AND symb_decoder(16#0d#)) OR
 					(reg_q119 AND symb_decoder(16#0c#)) OR
 					(reg_q117 AND symb_decoder(16#0a#)) OR
 					(reg_q117 AND symb_decoder(16#0c#)) OR
 					(reg_q117 AND symb_decoder(16#0d#)) OR
 					(reg_q117 AND symb_decoder(16#20#)) OR
 					(reg_q117 AND symb_decoder(16#09#));
reg_q119_init <= '0' ;
	p_reg_q119: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q119 <= reg_q119_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q119 <= reg_q119_init;
        else
          reg_q119 <= reg_q119_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q121_in <= (reg_q119 AND symb_decoder(16#76#)) OR
 					(reg_q119 AND symb_decoder(16#56#));
reg_q121_init <= '0' ;
	p_reg_q121: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q121 <= reg_q121_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q121 <= reg_q121_init;
        else
          reg_q121 <= reg_q121_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1207_in <= (reg_q1207 AND symb_decoder(16#30#)) OR
 					(reg_q1207 AND symb_decoder(16#33#)) OR
 					(reg_q1207 AND symb_decoder(16#37#)) OR
 					(reg_q1207 AND symb_decoder(16#32#)) OR
 					(reg_q1207 AND symb_decoder(16#31#)) OR
 					(reg_q1207 AND symb_decoder(16#38#)) OR
 					(reg_q1207 AND symb_decoder(16#36#)) OR
 					(reg_q1207 AND symb_decoder(16#35#)) OR
 					(reg_q1207 AND symb_decoder(16#34#)) OR
 					(reg_q1207 AND symb_decoder(16#39#)) OR
 					(reg_q1205 AND symb_decoder(16#38#)) OR
 					(reg_q1205 AND symb_decoder(16#34#)) OR
 					(reg_q1205 AND symb_decoder(16#35#)) OR
 					(reg_q1205 AND symb_decoder(16#33#)) OR
 					(reg_q1205 AND symb_decoder(16#32#)) OR
 					(reg_q1205 AND symb_decoder(16#37#)) OR
 					(reg_q1205 AND symb_decoder(16#31#)) OR
 					(reg_q1205 AND symb_decoder(16#39#)) OR
 					(reg_q1205 AND symb_decoder(16#30#)) OR
 					(reg_q1205 AND symb_decoder(16#36#));
reg_q1207_init <= '0' ;
	p_reg_q1207: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1207 <= reg_q1207_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1207 <= reg_q1207_init;
        else
          reg_q1207 <= reg_q1207_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1209_in <= (reg_q1207 AND symb_decoder(16#0c#)) OR
 					(reg_q1207 AND symb_decoder(16#0a#)) OR
 					(reg_q1207 AND symb_decoder(16#0d#)) OR
 					(reg_q1207 AND symb_decoder(16#20#)) OR
 					(reg_q1207 AND symb_decoder(16#09#)) OR
 					(reg_q1209 AND symb_decoder(16#09#)) OR
 					(reg_q1209 AND symb_decoder(16#0d#)) OR
 					(reg_q1209 AND symb_decoder(16#0c#)) OR
 					(reg_q1209 AND symb_decoder(16#20#)) OR
 					(reg_q1209 AND symb_decoder(16#0a#));
reg_q1209_init <= '0' ;
	p_reg_q1209: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1209 <= reg_q1209_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1209 <= reg_q1209_init;
        else
          reg_q1209 <= reg_q1209_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q74_in <= (reg_q72 AND symb_decoder(16#73#)) OR
 					(reg_q72 AND symb_decoder(16#53#));
reg_q74_init <= '0' ;
	p_reg_q74: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q74 <= reg_q74_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q74 <= reg_q74_init;
        else
          reg_q74 <= reg_q74_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q76_in <= (reg_q74 AND symb_decoder(16#45#)) OR
 					(reg_q74 AND symb_decoder(16#65#));
reg_q76_init <= '0' ;
	p_reg_q76: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q76 <= reg_q76_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q76 <= reg_q76_init;
        else
          reg_q76 <= reg_q76_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1189_in <= (reg_q1187 AND symb_decoder(16#42#)) OR
 					(reg_q1187 AND symb_decoder(16#62#));
reg_q1189_init <= '0' ;
	p_reg_q1189: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1189 <= reg_q1189_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1189 <= reg_q1189_init;
        else
          reg_q1189 <= reg_q1189_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1191_in <= (reg_q1189 AND symb_decoder(16#6c#)) OR
 					(reg_q1189 AND symb_decoder(16#4c#));
reg_q1191_init <= '0' ;
	p_reg_q1191: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1191 <= reg_q1191_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1191 <= reg_q1191_init;
        else
          reg_q1191 <= reg_q1191_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q262_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q262 AND symb_decoder(16#12#)) OR
 					(reg_q262 AND symb_decoder(16#61#)) OR
 					(reg_q262 AND symb_decoder(16#e5#)) OR
 					(reg_q262 AND symb_decoder(16#e7#)) OR
 					(reg_q262 AND symb_decoder(16#5f#)) OR
 					(reg_q262 AND symb_decoder(16#02#)) OR
 					(reg_q262 AND symb_decoder(16#89#)) OR
 					(reg_q262 AND symb_decoder(16#b3#)) OR
 					(reg_q262 AND symb_decoder(16#88#)) OR
 					(reg_q262 AND symb_decoder(16#8a#)) OR
 					(reg_q262 AND symb_decoder(16#8b#)) OR
 					(reg_q262 AND symb_decoder(16#34#)) OR
 					(reg_q262 AND symb_decoder(16#d0#)) OR
 					(reg_q262 AND symb_decoder(16#25#)) OR
 					(reg_q262 AND symb_decoder(16#b8#)) OR
 					(reg_q262 AND symb_decoder(16#14#)) OR
 					(reg_q262 AND symb_decoder(16#c4#)) OR
 					(reg_q262 AND symb_decoder(16#d6#)) OR
 					(reg_q262 AND symb_decoder(16#56#)) OR
 					(reg_q262 AND symb_decoder(16#3e#)) OR
 					(reg_q262 AND symb_decoder(16#66#)) OR
 					(reg_q262 AND symb_decoder(16#07#)) OR
 					(reg_q262 AND symb_decoder(16#40#)) OR
 					(reg_q262 AND symb_decoder(16#87#)) OR
 					(reg_q262 AND symb_decoder(16#d1#)) OR
 					(reg_q262 AND symb_decoder(16#de#)) OR
 					(reg_q262 AND symb_decoder(16#df#)) OR
 					(reg_q262 AND symb_decoder(16#9f#)) OR
 					(reg_q262 AND symb_decoder(16#1d#)) OR
 					(reg_q262 AND symb_decoder(16#80#)) OR
 					(reg_q262 AND symb_decoder(16#c7#)) OR
 					(reg_q262 AND symb_decoder(16#6d#)) OR
 					(reg_q262 AND symb_decoder(16#10#)) OR
 					(reg_q262 AND symb_decoder(16#0d#)) OR
 					(reg_q262 AND symb_decoder(16#f6#)) OR
 					(reg_q262 AND symb_decoder(16#1e#)) OR
 					(reg_q262 AND symb_decoder(16#6b#)) OR
 					(reg_q262 AND symb_decoder(16#21#)) OR
 					(reg_q262 AND symb_decoder(16#82#)) OR
 					(reg_q262 AND symb_decoder(16#2c#)) OR
 					(reg_q262 AND symb_decoder(16#9e#)) OR
 					(reg_q262 AND symb_decoder(16#74#)) OR
 					(reg_q262 AND symb_decoder(16#4d#)) OR
 					(reg_q262 AND symb_decoder(16#1b#)) OR
 					(reg_q262 AND symb_decoder(16#36#)) OR
 					(reg_q262 AND symb_decoder(16#f7#)) OR
 					(reg_q262 AND symb_decoder(16#91#)) OR
 					(reg_q262 AND symb_decoder(16#73#)) OR
 					(reg_q262 AND symb_decoder(16#ad#)) OR
 					(reg_q262 AND symb_decoder(16#b7#)) OR
 					(reg_q262 AND symb_decoder(16#2a#)) OR
 					(reg_q262 AND symb_decoder(16#2d#)) OR
 					(reg_q262 AND symb_decoder(16#75#)) OR
 					(reg_q262 AND symb_decoder(16#4f#)) OR
 					(reg_q262 AND symb_decoder(16#a0#)) OR
 					(reg_q262 AND symb_decoder(16#3c#)) OR
 					(reg_q262 AND symb_decoder(16#aa#)) OR
 					(reg_q262 AND symb_decoder(16#a8#)) OR
 					(reg_q262 AND symb_decoder(16#1a#)) OR
 					(reg_q262 AND symb_decoder(16#13#)) OR
 					(reg_q262 AND symb_decoder(16#3b#)) OR
 					(reg_q262 AND symb_decoder(16#8d#)) OR
 					(reg_q262 AND symb_decoder(16#7b#)) OR
 					(reg_q262 AND symb_decoder(16#42#)) OR
 					(reg_q262 AND symb_decoder(16#06#)) OR
 					(reg_q262 AND symb_decoder(16#b5#)) OR
 					(reg_q262 AND symb_decoder(16#ca#)) OR
 					(reg_q262 AND symb_decoder(16#5b#)) OR
 					(reg_q262 AND symb_decoder(16#64#)) OR
 					(reg_q262 AND symb_decoder(16#31#)) OR
 					(reg_q262 AND symb_decoder(16#35#)) OR
 					(reg_q262 AND symb_decoder(16#92#)) OR
 					(reg_q262 AND symb_decoder(16#4a#)) OR
 					(reg_q262 AND symb_decoder(16#2b#)) OR
 					(reg_q262 AND symb_decoder(16#96#)) OR
 					(reg_q262 AND symb_decoder(16#52#)) OR
 					(reg_q262 AND symb_decoder(16#48#)) OR
 					(reg_q262 AND symb_decoder(16#09#)) OR
 					(reg_q262 AND symb_decoder(16#e3#)) OR
 					(reg_q262 AND symb_decoder(16#cf#)) OR
 					(reg_q262 AND symb_decoder(16#ba#)) OR
 					(reg_q262 AND symb_decoder(16#0a#)) OR
 					(reg_q262 AND symb_decoder(16#a3#)) OR
 					(reg_q262 AND symb_decoder(16#6a#)) OR
 					(reg_q262 AND symb_decoder(16#f0#)) OR
 					(reg_q262 AND symb_decoder(16#00#)) OR
 					(reg_q262 AND symb_decoder(16#65#)) OR
 					(reg_q262 AND symb_decoder(16#1f#)) OR
 					(reg_q262 AND symb_decoder(16#24#)) OR
 					(reg_q262 AND symb_decoder(16#fb#)) OR
 					(reg_q262 AND symb_decoder(16#cc#)) OR
 					(reg_q262 AND symb_decoder(16#23#)) OR
 					(reg_q262 AND symb_decoder(16#01#)) OR
 					(reg_q262 AND symb_decoder(16#29#)) OR
 					(reg_q262 AND symb_decoder(16#57#)) OR
 					(reg_q262 AND symb_decoder(16#d7#)) OR
 					(reg_q262 AND symb_decoder(16#b6#)) OR
 					(reg_q262 AND symb_decoder(16#dd#)) OR
 					(reg_q262 AND symb_decoder(16#c5#)) OR
 					(reg_q262 AND symb_decoder(16#44#)) OR
 					(reg_q262 AND symb_decoder(16#f3#)) OR
 					(reg_q262 AND symb_decoder(16#fc#)) OR
 					(reg_q262 AND symb_decoder(16#9a#)) OR
 					(reg_q262 AND symb_decoder(16#8c#)) OR
 					(reg_q262 AND symb_decoder(16#77#)) OR
 					(reg_q262 AND symb_decoder(16#ec#)) OR
 					(reg_q262 AND symb_decoder(16#c2#)) OR
 					(reg_q262 AND symb_decoder(16#e9#)) OR
 					(reg_q262 AND symb_decoder(16#05#)) OR
 					(reg_q262 AND symb_decoder(16#03#)) OR
 					(reg_q262 AND symb_decoder(16#26#)) OR
 					(reg_q262 AND symb_decoder(16#16#)) OR
 					(reg_q262 AND symb_decoder(16#a5#)) OR
 					(reg_q262 AND symb_decoder(16#a7#)) OR
 					(reg_q262 AND symb_decoder(16#0b#)) OR
 					(reg_q262 AND symb_decoder(16#59#)) OR
 					(reg_q262 AND symb_decoder(16#c8#)) OR
 					(reg_q262 AND symb_decoder(16#53#)) OR
 					(reg_q262 AND symb_decoder(16#3d#)) OR
 					(reg_q262 AND symb_decoder(16#20#)) OR
 					(reg_q262 AND symb_decoder(16#99#)) OR
 					(reg_q262 AND symb_decoder(16#b2#)) OR
 					(reg_q262 AND symb_decoder(16#f1#)) OR
 					(reg_q262 AND symb_decoder(16#ac#)) OR
 					(reg_q262 AND symb_decoder(16#6f#)) OR
 					(reg_q262 AND symb_decoder(16#5e#)) OR
 					(reg_q262 AND symb_decoder(16#a4#)) OR
 					(reg_q262 AND symb_decoder(16#98#)) OR
 					(reg_q262 AND symb_decoder(16#27#)) OR
 					(reg_q262 AND symb_decoder(16#d9#)) OR
 					(reg_q262 AND symb_decoder(16#70#)) OR
 					(reg_q262 AND symb_decoder(16#15#)) OR
 					(reg_q262 AND symb_decoder(16#a9#)) OR
 					(reg_q262 AND symb_decoder(16#4b#)) OR
 					(reg_q262 AND symb_decoder(16#e4#)) OR
 					(reg_q262 AND symb_decoder(16#9b#)) OR
 					(reg_q262 AND symb_decoder(16#19#)) OR
 					(reg_q262 AND symb_decoder(16#90#)) OR
 					(reg_q262 AND symb_decoder(16#a6#)) OR
 					(reg_q262 AND symb_decoder(16#f8#)) OR
 					(reg_q262 AND symb_decoder(16#d3#)) OR
 					(reg_q262 AND symb_decoder(16#5c#)) OR
 					(reg_q262 AND symb_decoder(16#45#)) OR
 					(reg_q262 AND symb_decoder(16#b0#)) OR
 					(reg_q262 AND symb_decoder(16#fa#)) OR
 					(reg_q262 AND symb_decoder(16#54#)) OR
 					(reg_q262 AND symb_decoder(16#d8#)) OR
 					(reg_q262 AND symb_decoder(16#78#)) OR
 					(reg_q262 AND symb_decoder(16#3f#)) OR
 					(reg_q262 AND symb_decoder(16#f2#)) OR
 					(reg_q262 AND symb_decoder(16#4c#)) OR
 					(reg_q262 AND symb_decoder(16#6e#)) OR
 					(reg_q262 AND symb_decoder(16#be#)) OR
 					(reg_q262 AND symb_decoder(16#ce#)) OR
 					(reg_q262 AND symb_decoder(16#e8#)) OR
 					(reg_q262 AND symb_decoder(16#11#)) OR
 					(reg_q262 AND symb_decoder(16#dc#)) OR
 					(reg_q262 AND symb_decoder(16#0f#)) OR
 					(reg_q262 AND symb_decoder(16#b4#)) OR
 					(reg_q262 AND symb_decoder(16#08#)) OR
 					(reg_q262 AND symb_decoder(16#62#)) OR
 					(reg_q262 AND symb_decoder(16#f5#)) OR
 					(reg_q262 AND symb_decoder(16#c3#)) OR
 					(reg_q262 AND symb_decoder(16#60#)) OR
 					(reg_q262 AND symb_decoder(16#cd#)) OR
 					(reg_q262 AND symb_decoder(16#8e#)) OR
 					(reg_q262 AND symb_decoder(16#04#)) OR
 					(reg_q262 AND symb_decoder(16#fe#)) OR
 					(reg_q262 AND symb_decoder(16#7f#)) OR
 					(reg_q262 AND symb_decoder(16#ea#)) OR
 					(reg_q262 AND symb_decoder(16#ef#)) OR
 					(reg_q262 AND symb_decoder(16#71#)) OR
 					(reg_q262 AND symb_decoder(16#7c#)) OR
 					(reg_q262 AND symb_decoder(16#5d#)) OR
 					(reg_q262 AND symb_decoder(16#46#)) OR
 					(reg_q262 AND symb_decoder(16#d4#)) OR
 					(reg_q262 AND symb_decoder(16#d2#)) OR
 					(reg_q262 AND symb_decoder(16#3a#)) OR
 					(reg_q262 AND symb_decoder(16#72#)) OR
 					(reg_q262 AND symb_decoder(16#ee#)) OR
 					(reg_q262 AND symb_decoder(16#58#)) OR
 					(reg_q262 AND symb_decoder(16#79#)) OR
 					(reg_q262 AND symb_decoder(16#76#)) OR
 					(reg_q262 AND symb_decoder(16#2e#)) OR
 					(reg_q262 AND symb_decoder(16#e2#)) OR
 					(reg_q262 AND symb_decoder(16#28#)) OR
 					(reg_q262 AND symb_decoder(16#37#)) OR
 					(reg_q262 AND symb_decoder(16#9d#)) OR
 					(reg_q262 AND symb_decoder(16#1c#)) OR
 					(reg_q262 AND symb_decoder(16#ab#)) OR
 					(reg_q262 AND symb_decoder(16#ff#)) OR
 					(reg_q262 AND symb_decoder(16#33#)) OR
 					(reg_q262 AND symb_decoder(16#bb#)) OR
 					(reg_q262 AND symb_decoder(16#f4#)) OR
 					(reg_q262 AND symb_decoder(16#c1#)) OR
 					(reg_q262 AND symb_decoder(16#6c#)) OR
 					(reg_q262 AND symb_decoder(16#17#)) OR
 					(reg_q262 AND symb_decoder(16#bf#)) OR
 					(reg_q262 AND symb_decoder(16#94#)) OR
 					(reg_q262 AND symb_decoder(16#69#)) OR
 					(reg_q262 AND symb_decoder(16#ae#)) OR
 					(reg_q262 AND symb_decoder(16#4e#)) OR
 					(reg_q262 AND symb_decoder(16#c9#)) OR
 					(reg_q262 AND symb_decoder(16#bc#)) OR
 					(reg_q262 AND symb_decoder(16#30#)) OR
 					(reg_q262 AND symb_decoder(16#39#)) OR
 					(reg_q262 AND symb_decoder(16#e0#)) OR
 					(reg_q262 AND symb_decoder(16#9c#)) OR
 					(reg_q262 AND symb_decoder(16#8f#)) OR
 					(reg_q262 AND symb_decoder(16#b1#)) OR
 					(reg_q262 AND symb_decoder(16#e1#)) OR
 					(reg_q262 AND symb_decoder(16#e6#)) OR
 					(reg_q262 AND symb_decoder(16#93#)) OR
 					(reg_q262 AND symb_decoder(16#51#)) OR
 					(reg_q262 AND symb_decoder(16#da#)) OR
 					(reg_q262 AND symb_decoder(16#67#)) OR
 					(reg_q262 AND symb_decoder(16#7a#)) OR
 					(reg_q262 AND symb_decoder(16#68#)) OR
 					(reg_q262 AND symb_decoder(16#af#)) OR
 					(reg_q262 AND symb_decoder(16#a1#)) OR
 					(reg_q262 AND symb_decoder(16#83#)) OR
 					(reg_q262 AND symb_decoder(16#32#)) OR
 					(reg_q262 AND symb_decoder(16#b9#)) OR
 					(reg_q262 AND symb_decoder(16#d5#)) OR
 					(reg_q262 AND symb_decoder(16#bd#)) OR
 					(reg_q262 AND symb_decoder(16#97#)) OR
 					(reg_q262 AND symb_decoder(16#84#)) OR
 					(reg_q262 AND symb_decoder(16#7e#)) OR
 					(reg_q262 AND symb_decoder(16#db#)) OR
 					(reg_q262 AND symb_decoder(16#fd#)) OR
 					(reg_q262 AND symb_decoder(16#0c#)) OR
 					(reg_q262 AND symb_decoder(16#2f#)) OR
 					(reg_q262 AND symb_decoder(16#0e#)) OR
 					(reg_q262 AND symb_decoder(16#22#)) OR
 					(reg_q262 AND symb_decoder(16#7d#)) OR
 					(reg_q262 AND symb_decoder(16#43#)) OR
 					(reg_q262 AND symb_decoder(16#55#)) OR
 					(reg_q262 AND symb_decoder(16#95#)) OR
 					(reg_q262 AND symb_decoder(16#18#)) OR
 					(reg_q262 AND symb_decoder(16#50#)) OR
 					(reg_q262 AND symb_decoder(16#47#)) OR
 					(reg_q262 AND symb_decoder(16#41#)) OR
 					(reg_q262 AND symb_decoder(16#c6#)) OR
 					(reg_q262 AND symb_decoder(16#ed#)) OR
 					(reg_q262 AND symb_decoder(16#86#)) OR
 					(reg_q262 AND symb_decoder(16#38#)) OR
 					(reg_q262 AND symb_decoder(16#63#)) OR
 					(reg_q262 AND symb_decoder(16#c0#)) OR
 					(reg_q262 AND symb_decoder(16#49#)) OR
 					(reg_q262 AND symb_decoder(16#f9#)) OR
 					(reg_q262 AND symb_decoder(16#5a#)) OR
 					(reg_q262 AND symb_decoder(16#cb#)) OR
 					(reg_q262 AND symb_decoder(16#81#)) OR
 					(reg_q262 AND symb_decoder(16#eb#)) OR
 					(reg_q262 AND symb_decoder(16#85#)) OR
 					(reg_q262 AND symb_decoder(16#a2#));
reg_q262_init <= '0' ;
	p_reg_q262: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q262 <= reg_q262_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q262 <= reg_q262_init;
        else
          reg_q262 <= reg_q262_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1884_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1884 AND symb_decoder(16#d1#)) OR
 					(reg_q1884 AND symb_decoder(16#4f#)) OR
 					(reg_q1884 AND symb_decoder(16#17#)) OR
 					(reg_q1884 AND symb_decoder(16#38#)) OR
 					(reg_q1884 AND symb_decoder(16#23#)) OR
 					(reg_q1884 AND symb_decoder(16#ad#)) OR
 					(reg_q1884 AND symb_decoder(16#12#)) OR
 					(reg_q1884 AND symb_decoder(16#1f#)) OR
 					(reg_q1884 AND symb_decoder(16#c7#)) OR
 					(reg_q1884 AND symb_decoder(16#ec#)) OR
 					(reg_q1884 AND symb_decoder(16#e8#)) OR
 					(reg_q1884 AND symb_decoder(16#27#)) OR
 					(reg_q1884 AND symb_decoder(16#bf#)) OR
 					(reg_q1884 AND symb_decoder(16#33#)) OR
 					(reg_q1884 AND symb_decoder(16#a6#)) OR
 					(reg_q1884 AND symb_decoder(16#78#)) OR
 					(reg_q1884 AND symb_decoder(16#f2#)) OR
 					(reg_q1884 AND symb_decoder(16#00#)) OR
 					(reg_q1884 AND symb_decoder(16#4d#)) OR
 					(reg_q1884 AND symb_decoder(16#34#)) OR
 					(reg_q1884 AND symb_decoder(16#c0#)) OR
 					(reg_q1884 AND symb_decoder(16#a7#)) OR
 					(reg_q1884 AND symb_decoder(16#bd#)) OR
 					(reg_q1884 AND symb_decoder(16#fc#)) OR
 					(reg_q1884 AND symb_decoder(16#92#)) OR
 					(reg_q1884 AND symb_decoder(16#c9#)) OR
 					(reg_q1884 AND symb_decoder(16#ae#)) OR
 					(reg_q1884 AND symb_decoder(16#46#)) OR
 					(reg_q1884 AND symb_decoder(16#ff#)) OR
 					(reg_q1884 AND symb_decoder(16#8a#)) OR
 					(reg_q1884 AND symb_decoder(16#09#)) OR
 					(reg_q1884 AND symb_decoder(16#63#)) OR
 					(reg_q1884 AND symb_decoder(16#3e#)) OR
 					(reg_q1884 AND symb_decoder(16#14#)) OR
 					(reg_q1884 AND symb_decoder(16#1a#)) OR
 					(reg_q1884 AND symb_decoder(16#ab#)) OR
 					(reg_q1884 AND symb_decoder(16#dc#)) OR
 					(reg_q1884 AND symb_decoder(16#e5#)) OR
 					(reg_q1884 AND symb_decoder(16#20#)) OR
 					(reg_q1884 AND symb_decoder(16#60#)) OR
 					(reg_q1884 AND symb_decoder(16#1d#)) OR
 					(reg_q1884 AND symb_decoder(16#d8#)) OR
 					(reg_q1884 AND symb_decoder(16#76#)) OR
 					(reg_q1884 AND symb_decoder(16#55#)) OR
 					(reg_q1884 AND symb_decoder(16#aa#)) OR
 					(reg_q1884 AND symb_decoder(16#d0#)) OR
 					(reg_q1884 AND symb_decoder(16#45#)) OR
 					(reg_q1884 AND symb_decoder(16#56#)) OR
 					(reg_q1884 AND symb_decoder(16#9b#)) OR
 					(reg_q1884 AND symb_decoder(16#3d#)) OR
 					(reg_q1884 AND symb_decoder(16#04#)) OR
 					(reg_q1884 AND symb_decoder(16#85#)) OR
 					(reg_q1884 AND symb_decoder(16#89#)) OR
 					(reg_q1884 AND symb_decoder(16#a3#)) OR
 					(reg_q1884 AND symb_decoder(16#72#)) OR
 					(reg_q1884 AND symb_decoder(16#3b#)) OR
 					(reg_q1884 AND symb_decoder(16#c1#)) OR
 					(reg_q1884 AND symb_decoder(16#36#)) OR
 					(reg_q1884 AND symb_decoder(16#10#)) OR
 					(reg_q1884 AND symb_decoder(16#bb#)) OR
 					(reg_q1884 AND symb_decoder(16#7b#)) OR
 					(reg_q1884 AND symb_decoder(16#98#)) OR
 					(reg_q1884 AND symb_decoder(16#e6#)) OR
 					(reg_q1884 AND symb_decoder(16#db#)) OR
 					(reg_q1884 AND symb_decoder(16#2f#)) OR
 					(reg_q1884 AND symb_decoder(16#6b#)) OR
 					(reg_q1884 AND symb_decoder(16#06#)) OR
 					(reg_q1884 AND symb_decoder(16#95#)) OR
 					(reg_q1884 AND symb_decoder(16#87#)) OR
 					(reg_q1884 AND symb_decoder(16#e9#)) OR
 					(reg_q1884 AND symb_decoder(16#b6#)) OR
 					(reg_q1884 AND symb_decoder(16#de#)) OR
 					(reg_q1884 AND symb_decoder(16#9a#)) OR
 					(reg_q1884 AND symb_decoder(16#a5#)) OR
 					(reg_q1884 AND symb_decoder(16#16#)) OR
 					(reg_q1884 AND symb_decoder(16#3a#)) OR
 					(reg_q1884 AND symb_decoder(16#7e#)) OR
 					(reg_q1884 AND symb_decoder(16#6d#)) OR
 					(reg_q1884 AND symb_decoder(16#11#)) OR
 					(reg_q1884 AND symb_decoder(16#d7#)) OR
 					(reg_q1884 AND symb_decoder(16#f9#)) OR
 					(reg_q1884 AND symb_decoder(16#a0#)) OR
 					(reg_q1884 AND symb_decoder(16#bc#)) OR
 					(reg_q1884 AND symb_decoder(16#79#)) OR
 					(reg_q1884 AND symb_decoder(16#c5#)) OR
 					(reg_q1884 AND symb_decoder(16#7f#)) OR
 					(reg_q1884 AND symb_decoder(16#1e#)) OR
 					(reg_q1884 AND symb_decoder(16#d3#)) OR
 					(reg_q1884 AND symb_decoder(16#94#)) OR
 					(reg_q1884 AND symb_decoder(16#b5#)) OR
 					(reg_q1884 AND symb_decoder(16#0f#)) OR
 					(reg_q1884 AND symb_decoder(16#cf#)) OR
 					(reg_q1884 AND symb_decoder(16#13#)) OR
 					(reg_q1884 AND symb_decoder(16#f8#)) OR
 					(reg_q1884 AND symb_decoder(16#4a#)) OR
 					(reg_q1884 AND symb_decoder(16#62#)) OR
 					(reg_q1884 AND symb_decoder(16#c6#)) OR
 					(reg_q1884 AND symb_decoder(16#ed#)) OR
 					(reg_q1884 AND symb_decoder(16#b9#)) OR
 					(reg_q1884 AND symb_decoder(16#30#)) OR
 					(reg_q1884 AND symb_decoder(16#6f#)) OR
 					(reg_q1884 AND symb_decoder(16#35#)) OR
 					(reg_q1884 AND symb_decoder(16#65#)) OR
 					(reg_q1884 AND symb_decoder(16#82#)) OR
 					(reg_q1884 AND symb_decoder(16#be#)) OR
 					(reg_q1884 AND symb_decoder(16#8e#)) OR
 					(reg_q1884 AND symb_decoder(16#6a#)) OR
 					(reg_q1884 AND symb_decoder(16#40#)) OR
 					(reg_q1884 AND symb_decoder(16#81#)) OR
 					(reg_q1884 AND symb_decoder(16#ce#)) OR
 					(reg_q1884 AND symb_decoder(16#e1#)) OR
 					(reg_q1884 AND symb_decoder(16#7a#)) OR
 					(reg_q1884 AND symb_decoder(16#48#)) OR
 					(reg_q1884 AND symb_decoder(16#42#)) OR
 					(reg_q1884 AND symb_decoder(16#02#)) OR
 					(reg_q1884 AND symb_decoder(16#88#)) OR
 					(reg_q1884 AND symb_decoder(16#2d#)) OR
 					(reg_q1884 AND symb_decoder(16#64#)) OR
 					(reg_q1884 AND symb_decoder(16#5f#)) OR
 					(reg_q1884 AND symb_decoder(16#7d#)) OR
 					(reg_q1884 AND symb_decoder(16#69#)) OR
 					(reg_q1884 AND symb_decoder(16#c8#)) OR
 					(reg_q1884 AND symb_decoder(16#5a#)) OR
 					(reg_q1884 AND symb_decoder(16#df#)) OR
 					(reg_q1884 AND symb_decoder(16#2a#)) OR
 					(reg_q1884 AND symb_decoder(16#84#)) OR
 					(reg_q1884 AND symb_decoder(16#74#)) OR
 					(reg_q1884 AND symb_decoder(16#9c#)) OR
 					(reg_q1884 AND symb_decoder(16#03#)) OR
 					(reg_q1884 AND symb_decoder(16#7c#)) OR
 					(reg_q1884 AND symb_decoder(16#91#)) OR
 					(reg_q1884 AND symb_decoder(16#0b#)) OR
 					(reg_q1884 AND symb_decoder(16#2c#)) OR
 					(reg_q1884 AND symb_decoder(16#e7#)) OR
 					(reg_q1884 AND symb_decoder(16#b3#)) OR
 					(reg_q1884 AND symb_decoder(16#32#)) OR
 					(reg_q1884 AND symb_decoder(16#31#)) OR
 					(reg_q1884 AND symb_decoder(16#f7#)) OR
 					(reg_q1884 AND symb_decoder(16#80#)) OR
 					(reg_q1884 AND symb_decoder(16#41#)) OR
 					(reg_q1884 AND symb_decoder(16#b8#)) OR
 					(reg_q1884 AND symb_decoder(16#d4#)) OR
 					(reg_q1884 AND symb_decoder(16#dd#)) OR
 					(reg_q1884 AND symb_decoder(16#90#)) OR
 					(reg_q1884 AND symb_decoder(16#ba#)) OR
 					(reg_q1884 AND symb_decoder(16#e2#)) OR
 					(reg_q1884 AND symb_decoder(16#70#)) OR
 					(reg_q1884 AND symb_decoder(16#5c#)) OR
 					(reg_q1884 AND symb_decoder(16#f4#)) OR
 					(reg_q1884 AND symb_decoder(16#c4#)) OR
 					(reg_q1884 AND symb_decoder(16#ac#)) OR
 					(reg_q1884 AND symb_decoder(16#05#)) OR
 					(reg_q1884 AND symb_decoder(16#37#)) OR
 					(reg_q1884 AND symb_decoder(16#2b#)) OR
 					(reg_q1884 AND symb_decoder(16#d2#)) OR
 					(reg_q1884 AND symb_decoder(16#8b#)) OR
 					(reg_q1884 AND symb_decoder(16#5d#)) OR
 					(reg_q1884 AND symb_decoder(16#9f#)) OR
 					(reg_q1884 AND symb_decoder(16#22#)) OR
 					(reg_q1884 AND symb_decoder(16#97#)) OR
 					(reg_q1884 AND symb_decoder(16#fb#)) OR
 					(reg_q1884 AND symb_decoder(16#f3#)) OR
 					(reg_q1884 AND symb_decoder(16#fd#)) OR
 					(reg_q1884 AND symb_decoder(16#61#)) OR
 					(reg_q1884 AND symb_decoder(16#4c#)) OR
 					(reg_q1884 AND symb_decoder(16#19#)) OR
 					(reg_q1884 AND symb_decoder(16#6e#)) OR
 					(reg_q1884 AND symb_decoder(16#58#)) OR
 					(reg_q1884 AND symb_decoder(16#6c#)) OR
 					(reg_q1884 AND symb_decoder(16#53#)) OR
 					(reg_q1884 AND symb_decoder(16#93#)) OR
 					(reg_q1884 AND symb_decoder(16#1c#)) OR
 					(reg_q1884 AND symb_decoder(16#f5#)) OR
 					(reg_q1884 AND symb_decoder(16#ee#)) OR
 					(reg_q1884 AND symb_decoder(16#b7#)) OR
 					(reg_q1884 AND symb_decoder(16#50#)) OR
 					(reg_q1884 AND symb_decoder(16#3f#)) OR
 					(reg_q1884 AND symb_decoder(16#cc#)) OR
 					(reg_q1884 AND symb_decoder(16#eb#)) OR
 					(reg_q1884 AND symb_decoder(16#b4#)) OR
 					(reg_q1884 AND symb_decoder(16#f0#)) OR
 					(reg_q1884 AND symb_decoder(16#0c#)) OR
 					(reg_q1884 AND symb_decoder(16#67#)) OR
 					(reg_q1884 AND symb_decoder(16#e4#)) OR
 					(reg_q1884 AND symb_decoder(16#71#)) OR
 					(reg_q1884 AND symb_decoder(16#43#)) OR
 					(reg_q1884 AND symb_decoder(16#fa#)) OR
 					(reg_q1884 AND symb_decoder(16#e0#)) OR
 					(reg_q1884 AND symb_decoder(16#57#)) OR
 					(reg_q1884 AND symb_decoder(16#59#)) OR
 					(reg_q1884 AND symb_decoder(16#83#)) OR
 					(reg_q1884 AND symb_decoder(16#01#)) OR
 					(reg_q1884 AND symb_decoder(16#8f#)) OR
 					(reg_q1884 AND symb_decoder(16#47#)) OR
 					(reg_q1884 AND symb_decoder(16#b1#)) OR
 					(reg_q1884 AND symb_decoder(16#0a#)) OR
 					(reg_q1884 AND symb_decoder(16#28#)) OR
 					(reg_q1884 AND symb_decoder(16#9d#)) OR
 					(reg_q1884 AND symb_decoder(16#96#)) OR
 					(reg_q1884 AND symb_decoder(16#d6#)) OR
 					(reg_q1884 AND symb_decoder(16#25#)) OR
 					(reg_q1884 AND symb_decoder(16#a4#)) OR
 					(reg_q1884 AND symb_decoder(16#99#)) OR
 					(reg_q1884 AND symb_decoder(16#c2#)) OR
 					(reg_q1884 AND symb_decoder(16#54#)) OR
 					(reg_q1884 AND symb_decoder(16#18#)) OR
 					(reg_q1884 AND symb_decoder(16#da#)) OR
 					(reg_q1884 AND symb_decoder(16#73#)) OR
 					(reg_q1884 AND symb_decoder(16#5b#)) OR
 					(reg_q1884 AND symb_decoder(16#08#)) OR
 					(reg_q1884 AND symb_decoder(16#26#)) OR
 					(reg_q1884 AND symb_decoder(16#f6#)) OR
 					(reg_q1884 AND symb_decoder(16#a1#)) OR
 					(reg_q1884 AND symb_decoder(16#3c#)) OR
 					(reg_q1884 AND symb_decoder(16#b0#)) OR
 					(reg_q1884 AND symb_decoder(16#cb#)) OR
 					(reg_q1884 AND symb_decoder(16#1b#)) OR
 					(reg_q1884 AND symb_decoder(16#52#)) OR
 					(reg_q1884 AND symb_decoder(16#68#)) OR
 					(reg_q1884 AND symb_decoder(16#9e#)) OR
 					(reg_q1884 AND symb_decoder(16#a9#)) OR
 					(reg_q1884 AND symb_decoder(16#d9#)) OR
 					(reg_q1884 AND symb_decoder(16#ef#)) OR
 					(reg_q1884 AND symb_decoder(16#d5#)) OR
 					(reg_q1884 AND symb_decoder(16#07#)) OR
 					(reg_q1884 AND symb_decoder(16#66#)) OR
 					(reg_q1884 AND symb_decoder(16#21#)) OR
 					(reg_q1884 AND symb_decoder(16#29#)) OR
 					(reg_q1884 AND symb_decoder(16#0e#)) OR
 					(reg_q1884 AND symb_decoder(16#4b#)) OR
 					(reg_q1884 AND symb_decoder(16#fe#)) OR
 					(reg_q1884 AND symb_decoder(16#44#)) OR
 					(reg_q1884 AND symb_decoder(16#f1#)) OR
 					(reg_q1884 AND symb_decoder(16#a2#)) OR
 					(reg_q1884 AND symb_decoder(16#51#)) OR
 					(reg_q1884 AND symb_decoder(16#4e#)) OR
 					(reg_q1884 AND symb_decoder(16#af#)) OR
 					(reg_q1884 AND symb_decoder(16#b2#)) OR
 					(reg_q1884 AND symb_decoder(16#39#)) OR
 					(reg_q1884 AND symb_decoder(16#8d#)) OR
 					(reg_q1884 AND symb_decoder(16#2e#)) OR
 					(reg_q1884 AND symb_decoder(16#15#)) OR
 					(reg_q1884 AND symb_decoder(16#ea#)) OR
 					(reg_q1884 AND symb_decoder(16#77#)) OR
 					(reg_q1884 AND symb_decoder(16#86#)) OR
 					(reg_q1884 AND symb_decoder(16#a8#)) OR
 					(reg_q1884 AND symb_decoder(16#ca#)) OR
 					(reg_q1884 AND symb_decoder(16#c3#)) OR
 					(reg_q1884 AND symb_decoder(16#0d#)) OR
 					(reg_q1884 AND symb_decoder(16#24#)) OR
 					(reg_q1884 AND symb_decoder(16#e3#)) OR
 					(reg_q1884 AND symb_decoder(16#cd#)) OR
 					(reg_q1884 AND symb_decoder(16#75#)) OR
 					(reg_q1884 AND symb_decoder(16#49#)) OR
 					(reg_q1884 AND symb_decoder(16#5e#)) OR
 					(reg_q1884 AND symb_decoder(16#8c#));
reg_q1884_init <= '0' ;
	p_reg_q1884: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1884 <= reg_q1884_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1884 <= reg_q1884_init;
        else
          reg_q1884 <= reg_q1884_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2383_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2383 AND symb_decoder(16#c4#)) OR
 					(reg_q2383 AND symb_decoder(16#5e#)) OR
 					(reg_q2383 AND symb_decoder(16#96#)) OR
 					(reg_q2383 AND symb_decoder(16#62#)) OR
 					(reg_q2383 AND symb_decoder(16#02#)) OR
 					(reg_q2383 AND symb_decoder(16#45#)) OR
 					(reg_q2383 AND symb_decoder(16#09#)) OR
 					(reg_q2383 AND symb_decoder(16#16#)) OR
 					(reg_q2383 AND symb_decoder(16#b9#)) OR
 					(reg_q2383 AND symb_decoder(16#d4#)) OR
 					(reg_q2383 AND symb_decoder(16#8a#)) OR
 					(reg_q2383 AND symb_decoder(16#0c#)) OR
 					(reg_q2383 AND symb_decoder(16#d5#)) OR
 					(reg_q2383 AND symb_decoder(16#5c#)) OR
 					(reg_q2383 AND symb_decoder(16#55#)) OR
 					(reg_q2383 AND symb_decoder(16#f7#)) OR
 					(reg_q2383 AND symb_decoder(16#83#)) OR
 					(reg_q2383 AND symb_decoder(16#5a#)) OR
 					(reg_q2383 AND symb_decoder(16#ef#)) OR
 					(reg_q2383 AND symb_decoder(16#c9#)) OR
 					(reg_q2383 AND symb_decoder(16#9e#)) OR
 					(reg_q2383 AND symb_decoder(16#08#)) OR
 					(reg_q2383 AND symb_decoder(16#1b#)) OR
 					(reg_q2383 AND symb_decoder(16#3e#)) OR
 					(reg_q2383 AND symb_decoder(16#1a#)) OR
 					(reg_q2383 AND symb_decoder(16#48#)) OR
 					(reg_q2383 AND symb_decoder(16#de#)) OR
 					(reg_q2383 AND symb_decoder(16#63#)) OR
 					(reg_q2383 AND symb_decoder(16#dc#)) OR
 					(reg_q2383 AND symb_decoder(16#05#)) OR
 					(reg_q2383 AND symb_decoder(16#a6#)) OR
 					(reg_q2383 AND symb_decoder(16#46#)) OR
 					(reg_q2383 AND symb_decoder(16#56#)) OR
 					(reg_q2383 AND symb_decoder(16#66#)) OR
 					(reg_q2383 AND symb_decoder(16#e2#)) OR
 					(reg_q2383 AND symb_decoder(16#23#)) OR
 					(reg_q2383 AND symb_decoder(16#f1#)) OR
 					(reg_q2383 AND symb_decoder(16#9c#)) OR
 					(reg_q2383 AND symb_decoder(16#b0#)) OR
 					(reg_q2383 AND symb_decoder(16#f8#)) OR
 					(reg_q2383 AND symb_decoder(16#e0#)) OR
 					(reg_q2383 AND symb_decoder(16#20#)) OR
 					(reg_q2383 AND symb_decoder(16#84#)) OR
 					(reg_q2383 AND symb_decoder(16#29#)) OR
 					(reg_q2383 AND symb_decoder(16#e7#)) OR
 					(reg_q2383 AND symb_decoder(16#99#)) OR
 					(reg_q2383 AND symb_decoder(16#ba#)) OR
 					(reg_q2383 AND symb_decoder(16#34#)) OR
 					(reg_q2383 AND symb_decoder(16#53#)) OR
 					(reg_q2383 AND symb_decoder(16#93#)) OR
 					(reg_q2383 AND symb_decoder(16#fa#)) OR
 					(reg_q2383 AND symb_decoder(16#0a#)) OR
 					(reg_q2383 AND symb_decoder(16#d8#)) OR
 					(reg_q2383 AND symb_decoder(16#d3#)) OR
 					(reg_q2383 AND symb_decoder(16#35#)) OR
 					(reg_q2383 AND symb_decoder(16#b6#)) OR
 					(reg_q2383 AND symb_decoder(16#6a#)) OR
 					(reg_q2383 AND symb_decoder(16#90#)) OR
 					(reg_q2383 AND symb_decoder(16#a3#)) OR
 					(reg_q2383 AND symb_decoder(16#0d#)) OR
 					(reg_q2383 AND symb_decoder(16#1d#)) OR
 					(reg_q2383 AND symb_decoder(16#be#)) OR
 					(reg_q2383 AND symb_decoder(16#15#)) OR
 					(reg_q2383 AND symb_decoder(16#39#)) OR
 					(reg_q2383 AND symb_decoder(16#cf#)) OR
 					(reg_q2383 AND symb_decoder(16#1f#)) OR
 					(reg_q2383 AND symb_decoder(16#76#)) OR
 					(reg_q2383 AND symb_decoder(16#2b#)) OR
 					(reg_q2383 AND symb_decoder(16#c6#)) OR
 					(reg_q2383 AND symb_decoder(16#95#)) OR
 					(reg_q2383 AND symb_decoder(16#b1#)) OR
 					(reg_q2383 AND symb_decoder(16#8f#)) OR
 					(reg_q2383 AND symb_decoder(16#f2#)) OR
 					(reg_q2383 AND symb_decoder(16#c1#)) OR
 					(reg_q2383 AND symb_decoder(16#6e#)) OR
 					(reg_q2383 AND symb_decoder(16#40#)) OR
 					(reg_q2383 AND symb_decoder(16#42#)) OR
 					(reg_q2383 AND symb_decoder(16#a0#)) OR
 					(reg_q2383 AND symb_decoder(16#79#)) OR
 					(reg_q2383 AND symb_decoder(16#64#)) OR
 					(reg_q2383 AND symb_decoder(16#72#)) OR
 					(reg_q2383 AND symb_decoder(16#cd#)) OR
 					(reg_q2383 AND symb_decoder(16#c0#)) OR
 					(reg_q2383 AND symb_decoder(16#d9#)) OR
 					(reg_q2383 AND symb_decoder(16#49#)) OR
 					(reg_q2383 AND symb_decoder(16#a1#)) OR
 					(reg_q2383 AND symb_decoder(16#7c#)) OR
 					(reg_q2383 AND symb_decoder(16#ad#)) OR
 					(reg_q2383 AND symb_decoder(16#a5#)) OR
 					(reg_q2383 AND symb_decoder(16#57#)) OR
 					(reg_q2383 AND symb_decoder(16#df#)) OR
 					(reg_q2383 AND symb_decoder(16#ae#)) OR
 					(reg_q2383 AND symb_decoder(16#f0#)) OR
 					(reg_q2383 AND symb_decoder(16#c3#)) OR
 					(reg_q2383 AND symb_decoder(16#33#)) OR
 					(reg_q2383 AND symb_decoder(16#2a#)) OR
 					(reg_q2383 AND symb_decoder(16#82#)) OR
 					(reg_q2383 AND symb_decoder(16#f9#)) OR
 					(reg_q2383 AND symb_decoder(16#cb#)) OR
 					(reg_q2383 AND symb_decoder(16#9d#)) OR
 					(reg_q2383 AND symb_decoder(16#b5#)) OR
 					(reg_q2383 AND symb_decoder(16#18#)) OR
 					(reg_q2383 AND symb_decoder(16#f5#)) OR
 					(reg_q2383 AND symb_decoder(16#da#)) OR
 					(reg_q2383 AND symb_decoder(16#41#)) OR
 					(reg_q2383 AND symb_decoder(16#71#)) OR
 					(reg_q2383 AND symb_decoder(16#78#)) OR
 					(reg_q2383 AND symb_decoder(16#3f#)) OR
 					(reg_q2383 AND symb_decoder(16#6f#)) OR
 					(reg_q2383 AND symb_decoder(16#c2#)) OR
 					(reg_q2383 AND symb_decoder(16#ff#)) OR
 					(reg_q2383 AND symb_decoder(16#4a#)) OR
 					(reg_q2383 AND symb_decoder(16#a2#)) OR
 					(reg_q2383 AND symb_decoder(16#fc#)) OR
 					(reg_q2383 AND symb_decoder(16#59#)) OR
 					(reg_q2383 AND symb_decoder(16#a9#)) OR
 					(reg_q2383 AND symb_decoder(16#3c#)) OR
 					(reg_q2383 AND symb_decoder(16#e3#)) OR
 					(reg_q2383 AND symb_decoder(16#e1#)) OR
 					(reg_q2383 AND symb_decoder(16#fe#)) OR
 					(reg_q2383 AND symb_decoder(16#13#)) OR
 					(reg_q2383 AND symb_decoder(16#ee#)) OR
 					(reg_q2383 AND symb_decoder(16#2c#)) OR
 					(reg_q2383 AND symb_decoder(16#4f#)) OR
 					(reg_q2383 AND symb_decoder(16#54#)) OR
 					(reg_q2383 AND symb_decoder(16#f4#)) OR
 					(reg_q2383 AND symb_decoder(16#bf#)) OR
 					(reg_q2383 AND symb_decoder(16#2d#)) OR
 					(reg_q2383 AND symb_decoder(16#65#)) OR
 					(reg_q2383 AND symb_decoder(16#ca#)) OR
 					(reg_q2383 AND symb_decoder(16#4b#)) OR
 					(reg_q2383 AND symb_decoder(16#7d#)) OR
 					(reg_q2383 AND symb_decoder(16#0f#)) OR
 					(reg_q2383 AND symb_decoder(16#88#)) OR
 					(reg_q2383 AND symb_decoder(16#bc#)) OR
 					(reg_q2383 AND symb_decoder(16#73#)) OR
 					(reg_q2383 AND symb_decoder(16#6c#)) OR
 					(reg_q2383 AND symb_decoder(16#12#)) OR
 					(reg_q2383 AND symb_decoder(16#4c#)) OR
 					(reg_q2383 AND symb_decoder(16#25#)) OR
 					(reg_q2383 AND symb_decoder(16#ed#)) OR
 					(reg_q2383 AND symb_decoder(16#75#)) OR
 					(reg_q2383 AND symb_decoder(16#c5#)) OR
 					(reg_q2383 AND symb_decoder(16#ce#)) OR
 					(reg_q2383 AND symb_decoder(16#bd#)) OR
 					(reg_q2383 AND symb_decoder(16#36#)) OR
 					(reg_q2383 AND symb_decoder(16#db#)) OR
 					(reg_q2383 AND symb_decoder(16#cc#)) OR
 					(reg_q2383 AND symb_decoder(16#21#)) OR
 					(reg_q2383 AND symb_decoder(16#5d#)) OR
 					(reg_q2383 AND symb_decoder(16#d2#)) OR
 					(reg_q2383 AND symb_decoder(16#4e#)) OR
 					(reg_q2383 AND symb_decoder(16#a4#)) OR
 					(reg_q2383 AND symb_decoder(16#22#)) OR
 					(reg_q2383 AND symb_decoder(16#d6#)) OR
 					(reg_q2383 AND symb_decoder(16#5b#)) OR
 					(reg_q2383 AND symb_decoder(16#8b#)) OR
 					(reg_q2383 AND symb_decoder(16#0e#)) OR
 					(reg_q2383 AND symb_decoder(16#86#)) OR
 					(reg_q2383 AND symb_decoder(16#e9#)) OR
 					(reg_q2383 AND symb_decoder(16#2f#)) OR
 					(reg_q2383 AND symb_decoder(16#4d#)) OR
 					(reg_q2383 AND symb_decoder(16#03#)) OR
 					(reg_q2383 AND symb_decoder(16#d7#)) OR
 					(reg_q2383 AND symb_decoder(16#32#)) OR
 					(reg_q2383 AND symb_decoder(16#80#)) OR
 					(reg_q2383 AND symb_decoder(16#d0#)) OR
 					(reg_q2383 AND symb_decoder(16#7b#)) OR
 					(reg_q2383 AND symb_decoder(16#43#)) OR
 					(reg_q2383 AND symb_decoder(16#aa#)) OR
 					(reg_q2383 AND symb_decoder(16#e4#)) OR
 					(reg_q2383 AND symb_decoder(16#fd#)) OR
 					(reg_q2383 AND symb_decoder(16#77#)) OR
 					(reg_q2383 AND symb_decoder(16#7e#)) OR
 					(reg_q2383 AND symb_decoder(16#89#)) OR
 					(reg_q2383 AND symb_decoder(16#3d#)) OR
 					(reg_q2383 AND symb_decoder(16#b3#)) OR
 					(reg_q2383 AND symb_decoder(16#d1#)) OR
 					(reg_q2383 AND symb_decoder(16#00#)) OR
 					(reg_q2383 AND symb_decoder(16#47#)) OR
 					(reg_q2383 AND symb_decoder(16#61#)) OR
 					(reg_q2383 AND symb_decoder(16#87#)) OR
 					(reg_q2383 AND symb_decoder(16#5f#)) OR
 					(reg_q2383 AND symb_decoder(16#27#)) OR
 					(reg_q2383 AND symb_decoder(16#26#)) OR
 					(reg_q2383 AND symb_decoder(16#30#)) OR
 					(reg_q2383 AND symb_decoder(16#31#)) OR
 					(reg_q2383 AND symb_decoder(16#14#)) OR
 					(reg_q2383 AND symb_decoder(16#f3#)) OR
 					(reg_q2383 AND symb_decoder(16#97#)) OR
 					(reg_q2383 AND symb_decoder(16#1c#)) OR
 					(reg_q2383 AND symb_decoder(16#8c#)) OR
 					(reg_q2383 AND symb_decoder(16#e8#)) OR
 					(reg_q2383 AND symb_decoder(16#24#)) OR
 					(reg_q2383 AND symb_decoder(16#a8#)) OR
 					(reg_q2383 AND symb_decoder(16#70#)) OR
 					(reg_q2383 AND symb_decoder(16#04#)) OR
 					(reg_q2383 AND symb_decoder(16#0b#)) OR
 					(reg_q2383 AND symb_decoder(16#7f#)) OR
 					(reg_q2383 AND symb_decoder(16#06#)) OR
 					(reg_q2383 AND symb_decoder(16#3a#)) OR
 					(reg_q2383 AND symb_decoder(16#10#)) OR
 					(reg_q2383 AND symb_decoder(16#b8#)) OR
 					(reg_q2383 AND symb_decoder(16#51#)) OR
 					(reg_q2383 AND symb_decoder(16#e6#)) OR
 					(reg_q2383 AND symb_decoder(16#81#)) OR
 					(reg_q2383 AND symb_decoder(16#a7#)) OR
 					(reg_q2383 AND symb_decoder(16#69#)) OR
 					(reg_q2383 AND symb_decoder(16#60#)) OR
 					(reg_q2383 AND symb_decoder(16#8d#)) OR
 					(reg_q2383 AND symb_decoder(16#28#)) OR
 					(reg_q2383 AND symb_decoder(16#6d#)) OR
 					(reg_q2383 AND symb_decoder(16#fb#)) OR
 					(reg_q2383 AND symb_decoder(16#1e#)) OR
 					(reg_q2383 AND symb_decoder(16#2e#)) OR
 					(reg_q2383 AND symb_decoder(16#af#)) OR
 					(reg_q2383 AND symb_decoder(16#bb#)) OR
 					(reg_q2383 AND symb_decoder(16#9a#)) OR
 					(reg_q2383 AND symb_decoder(16#52#)) OR
 					(reg_q2383 AND symb_decoder(16#44#)) OR
 					(reg_q2383 AND symb_decoder(16#dd#)) OR
 					(reg_q2383 AND symb_decoder(16#68#)) OR
 					(reg_q2383 AND symb_decoder(16#19#)) OR
 					(reg_q2383 AND symb_decoder(16#07#)) OR
 					(reg_q2383 AND symb_decoder(16#7a#)) OR
 					(reg_q2383 AND symb_decoder(16#37#)) OR
 					(reg_q2383 AND symb_decoder(16#e5#)) OR
 					(reg_q2383 AND symb_decoder(16#eb#)) OR
 					(reg_q2383 AND symb_decoder(16#17#)) OR
 					(reg_q2383 AND symb_decoder(16#6b#)) OR
 					(reg_q2383 AND symb_decoder(16#c8#)) OR
 					(reg_q2383 AND symb_decoder(16#3b#)) OR
 					(reg_q2383 AND symb_decoder(16#ec#)) OR
 					(reg_q2383 AND symb_decoder(16#01#)) OR
 					(reg_q2383 AND symb_decoder(16#ab#)) OR
 					(reg_q2383 AND symb_decoder(16#b2#)) OR
 					(reg_q2383 AND symb_decoder(16#94#)) OR
 					(reg_q2383 AND symb_decoder(16#98#)) OR
 					(reg_q2383 AND symb_decoder(16#11#)) OR
 					(reg_q2383 AND symb_decoder(16#f6#)) OR
 					(reg_q2383 AND symb_decoder(16#85#)) OR
 					(reg_q2383 AND symb_decoder(16#58#)) OR
 					(reg_q2383 AND symb_decoder(16#ac#)) OR
 					(reg_q2383 AND symb_decoder(16#b4#)) OR
 					(reg_q2383 AND symb_decoder(16#38#)) OR
 					(reg_q2383 AND symb_decoder(16#92#)) OR
 					(reg_q2383 AND symb_decoder(16#b7#)) OR
 					(reg_q2383 AND symb_decoder(16#67#)) OR
 					(reg_q2383 AND symb_decoder(16#91#)) OR
 					(reg_q2383 AND symb_decoder(16#ea#)) OR
 					(reg_q2383 AND symb_decoder(16#c7#)) OR
 					(reg_q2383 AND symb_decoder(16#9b#)) OR
 					(reg_q2383 AND symb_decoder(16#9f#)) OR
 					(reg_q2383 AND symb_decoder(16#50#)) OR
 					(reg_q2383 AND symb_decoder(16#74#)) OR
 					(reg_q2383 AND symb_decoder(16#8e#));
reg_q2383_init <= '0' ;
	p_reg_q2383: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2383 <= reg_q2383_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2383 <= reg_q2383_init;
        else
          reg_q2383 <= reg_q2383_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q414_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q414 AND symb_decoder(16#ec#)) OR
 					(reg_q414 AND symb_decoder(16#15#)) OR
 					(reg_q414 AND symb_decoder(16#7c#)) OR
 					(reg_q414 AND symb_decoder(16#6e#)) OR
 					(reg_q414 AND symb_decoder(16#db#)) OR
 					(reg_q414 AND symb_decoder(16#fb#)) OR
 					(reg_q414 AND symb_decoder(16#ff#)) OR
 					(reg_q414 AND symb_decoder(16#1a#)) OR
 					(reg_q414 AND symb_decoder(16#49#)) OR
 					(reg_q414 AND symb_decoder(16#5e#)) OR
 					(reg_q414 AND symb_decoder(16#5a#)) OR
 					(reg_q414 AND symb_decoder(16#3d#)) OR
 					(reg_q414 AND symb_decoder(16#94#)) OR
 					(reg_q414 AND symb_decoder(16#48#)) OR
 					(reg_q414 AND symb_decoder(16#02#)) OR
 					(reg_q414 AND symb_decoder(16#c8#)) OR
 					(reg_q414 AND symb_decoder(16#36#)) OR
 					(reg_q414 AND symb_decoder(16#41#)) OR
 					(reg_q414 AND symb_decoder(16#04#)) OR
 					(reg_q414 AND symb_decoder(16#33#)) OR
 					(reg_q414 AND symb_decoder(16#da#)) OR
 					(reg_q414 AND symb_decoder(16#3a#)) OR
 					(reg_q414 AND symb_decoder(16#7d#)) OR
 					(reg_q414 AND symb_decoder(16#ca#)) OR
 					(reg_q414 AND symb_decoder(16#df#)) OR
 					(reg_q414 AND symb_decoder(16#0e#)) OR
 					(reg_q414 AND symb_decoder(16#16#)) OR
 					(reg_q414 AND symb_decoder(16#6d#)) OR
 					(reg_q414 AND symb_decoder(16#8c#)) OR
 					(reg_q414 AND symb_decoder(16#8e#)) OR
 					(reg_q414 AND symb_decoder(16#96#)) OR
 					(reg_q414 AND symb_decoder(16#c5#)) OR
 					(reg_q414 AND symb_decoder(16#4d#)) OR
 					(reg_q414 AND symb_decoder(16#5d#)) OR
 					(reg_q414 AND symb_decoder(16#a5#)) OR
 					(reg_q414 AND symb_decoder(16#c2#)) OR
 					(reg_q414 AND symb_decoder(16#c6#)) OR
 					(reg_q414 AND symb_decoder(16#fe#)) OR
 					(reg_q414 AND symb_decoder(16#69#)) OR
 					(reg_q414 AND symb_decoder(16#ab#)) OR
 					(reg_q414 AND symb_decoder(16#e4#)) OR
 					(reg_q414 AND symb_decoder(16#be#)) OR
 					(reg_q414 AND symb_decoder(16#c3#)) OR
 					(reg_q414 AND symb_decoder(16#06#)) OR
 					(reg_q414 AND symb_decoder(16#f4#)) OR
 					(reg_q414 AND symb_decoder(16#a7#)) OR
 					(reg_q414 AND symb_decoder(16#20#)) OR
 					(reg_q414 AND symb_decoder(16#e9#)) OR
 					(reg_q414 AND symb_decoder(16#4c#)) OR
 					(reg_q414 AND symb_decoder(16#85#)) OR
 					(reg_q414 AND symb_decoder(16#0c#)) OR
 					(reg_q414 AND symb_decoder(16#14#)) OR
 					(reg_q414 AND symb_decoder(16#e6#)) OR
 					(reg_q414 AND symb_decoder(16#9b#)) OR
 					(reg_q414 AND symb_decoder(16#30#)) OR
 					(reg_q414 AND symb_decoder(16#11#)) OR
 					(reg_q414 AND symb_decoder(16#0a#)) OR
 					(reg_q414 AND symb_decoder(16#95#)) OR
 					(reg_q414 AND symb_decoder(16#38#)) OR
 					(reg_q414 AND symb_decoder(16#24#)) OR
 					(reg_q414 AND symb_decoder(16#f7#)) OR
 					(reg_q414 AND symb_decoder(16#9d#)) OR
 					(reg_q414 AND symb_decoder(16#9f#)) OR
 					(reg_q414 AND symb_decoder(16#fd#)) OR
 					(reg_q414 AND symb_decoder(16#87#)) OR
 					(reg_q414 AND symb_decoder(16#65#)) OR
 					(reg_q414 AND symb_decoder(16#13#)) OR
 					(reg_q414 AND symb_decoder(16#26#)) OR
 					(reg_q414 AND symb_decoder(16#b0#)) OR
 					(reg_q414 AND symb_decoder(16#ad#)) OR
 					(reg_q414 AND symb_decoder(16#91#)) OR
 					(reg_q414 AND symb_decoder(16#6c#)) OR
 					(reg_q414 AND symb_decoder(16#2b#)) OR
 					(reg_q414 AND symb_decoder(16#0b#)) OR
 					(reg_q414 AND symb_decoder(16#af#)) OR
 					(reg_q414 AND symb_decoder(16#5f#)) OR
 					(reg_q414 AND symb_decoder(16#89#)) OR
 					(reg_q414 AND symb_decoder(16#f8#)) OR
 					(reg_q414 AND symb_decoder(16#d2#)) OR
 					(reg_q414 AND symb_decoder(16#66#)) OR
 					(reg_q414 AND symb_decoder(16#b1#)) OR
 					(reg_q414 AND symb_decoder(16#b4#)) OR
 					(reg_q414 AND symb_decoder(16#fa#)) OR
 					(reg_q414 AND symb_decoder(16#22#)) OR
 					(reg_q414 AND symb_decoder(16#34#)) OR
 					(reg_q414 AND symb_decoder(16#4e#)) OR
 					(reg_q414 AND symb_decoder(16#cf#)) OR
 					(reg_q414 AND symb_decoder(16#70#)) OR
 					(reg_q414 AND symb_decoder(16#e0#)) OR
 					(reg_q414 AND symb_decoder(16#b5#)) OR
 					(reg_q414 AND symb_decoder(16#75#)) OR
 					(reg_q414 AND symb_decoder(16#57#)) OR
 					(reg_q414 AND symb_decoder(16#68#)) OR
 					(reg_q414 AND symb_decoder(16#de#)) OR
 					(reg_q414 AND symb_decoder(16#50#)) OR
 					(reg_q414 AND symb_decoder(16#ba#)) OR
 					(reg_q414 AND symb_decoder(16#4b#)) OR
 					(reg_q414 AND symb_decoder(16#c4#)) OR
 					(reg_q414 AND symb_decoder(16#c9#)) OR
 					(reg_q414 AND symb_decoder(16#f6#)) OR
 					(reg_q414 AND symb_decoder(16#e5#)) OR
 					(reg_q414 AND symb_decoder(16#f5#)) OR
 					(reg_q414 AND symb_decoder(16#e2#)) OR
 					(reg_q414 AND symb_decoder(16#6a#)) OR
 					(reg_q414 AND symb_decoder(16#a4#)) OR
 					(reg_q414 AND symb_decoder(16#25#)) OR
 					(reg_q414 AND symb_decoder(16#3e#)) OR
 					(reg_q414 AND symb_decoder(16#97#)) OR
 					(reg_q414 AND symb_decoder(16#44#)) OR
 					(reg_q414 AND symb_decoder(16#8a#)) OR
 					(reg_q414 AND symb_decoder(16#64#)) OR
 					(reg_q414 AND symb_decoder(16#45#)) OR
 					(reg_q414 AND symb_decoder(16#ef#)) OR
 					(reg_q414 AND symb_decoder(16#a1#)) OR
 					(reg_q414 AND symb_decoder(16#8b#)) OR
 					(reg_q414 AND symb_decoder(16#f1#)) OR
 					(reg_q414 AND symb_decoder(16#b3#)) OR
 					(reg_q414 AND symb_decoder(16#1f#)) OR
 					(reg_q414 AND symb_decoder(16#c7#)) OR
 					(reg_q414 AND symb_decoder(16#47#)) OR
 					(reg_q414 AND symb_decoder(16#46#)) OR
 					(reg_q414 AND symb_decoder(16#b2#)) OR
 					(reg_q414 AND symb_decoder(16#cc#)) OR
 					(reg_q414 AND symb_decoder(16#a0#)) OR
 					(reg_q414 AND symb_decoder(16#77#)) OR
 					(reg_q414 AND symb_decoder(16#37#)) OR
 					(reg_q414 AND symb_decoder(16#32#)) OR
 					(reg_q414 AND symb_decoder(16#7a#)) OR
 					(reg_q414 AND symb_decoder(16#d0#)) OR
 					(reg_q414 AND symb_decoder(16#7e#)) OR
 					(reg_q414 AND symb_decoder(16#2a#)) OR
 					(reg_q414 AND symb_decoder(16#29#)) OR
 					(reg_q414 AND symb_decoder(16#55#)) OR
 					(reg_q414 AND symb_decoder(16#ae#)) OR
 					(reg_q414 AND symb_decoder(16#c1#)) OR
 					(reg_q414 AND symb_decoder(16#aa#)) OR
 					(reg_q414 AND symb_decoder(16#b8#)) OR
 					(reg_q414 AND symb_decoder(16#12#)) OR
 					(reg_q414 AND symb_decoder(16#71#)) OR
 					(reg_q414 AND symb_decoder(16#72#)) OR
 					(reg_q414 AND symb_decoder(16#42#)) OR
 					(reg_q414 AND symb_decoder(16#f2#)) OR
 					(reg_q414 AND symb_decoder(16#8d#)) OR
 					(reg_q414 AND symb_decoder(16#59#)) OR
 					(reg_q414 AND symb_decoder(16#d7#)) OR
 					(reg_q414 AND symb_decoder(16#eb#)) OR
 					(reg_q414 AND symb_decoder(16#cd#)) OR
 					(reg_q414 AND symb_decoder(16#0f#)) OR
 					(reg_q414 AND symb_decoder(16#dd#)) OR
 					(reg_q414 AND symb_decoder(16#5b#)) OR
 					(reg_q414 AND symb_decoder(16#d4#)) OR
 					(reg_q414 AND symb_decoder(16#d8#)) OR
 					(reg_q414 AND symb_decoder(16#73#)) OR
 					(reg_q414 AND symb_decoder(16#82#)) OR
 					(reg_q414 AND symb_decoder(16#4a#)) OR
 					(reg_q414 AND symb_decoder(16#86#)) OR
 					(reg_q414 AND symb_decoder(16#2d#)) OR
 					(reg_q414 AND symb_decoder(16#53#)) OR
 					(reg_q414 AND symb_decoder(16#4f#)) OR
 					(reg_q414 AND symb_decoder(16#1d#)) OR
 					(reg_q414 AND symb_decoder(16#ee#)) OR
 					(reg_q414 AND symb_decoder(16#bc#)) OR
 					(reg_q414 AND symb_decoder(16#09#)) OR
 					(reg_q414 AND symb_decoder(16#bb#)) OR
 					(reg_q414 AND symb_decoder(16#61#)) OR
 					(reg_q414 AND symb_decoder(16#fc#)) OR
 					(reg_q414 AND symb_decoder(16#74#)) OR
 					(reg_q414 AND symb_decoder(16#a6#)) OR
 					(reg_q414 AND symb_decoder(16#07#)) OR
 					(reg_q414 AND symb_decoder(16#83#)) OR
 					(reg_q414 AND symb_decoder(16#0d#)) OR
 					(reg_q414 AND symb_decoder(16#93#)) OR
 					(reg_q414 AND symb_decoder(16#81#)) OR
 					(reg_q414 AND symb_decoder(16#17#)) OR
 					(reg_q414 AND symb_decoder(16#43#)) OR
 					(reg_q414 AND symb_decoder(16#84#)) OR
 					(reg_q414 AND symb_decoder(16#d5#)) OR
 					(reg_q414 AND symb_decoder(16#78#)) OR
 					(reg_q414 AND symb_decoder(16#88#)) OR
 					(reg_q414 AND symb_decoder(16#21#)) OR
 					(reg_q414 AND symb_decoder(16#9a#)) OR
 					(reg_q414 AND symb_decoder(16#e7#)) OR
 					(reg_q414 AND symb_decoder(16#a9#)) OR
 					(reg_q414 AND symb_decoder(16#7f#)) OR
 					(reg_q414 AND symb_decoder(16#1c#)) OR
 					(reg_q414 AND symb_decoder(16#79#)) OR
 					(reg_q414 AND symb_decoder(16#2f#)) OR
 					(reg_q414 AND symb_decoder(16#63#)) OR
 					(reg_q414 AND symb_decoder(16#ed#)) OR
 					(reg_q414 AND symb_decoder(16#54#)) OR
 					(reg_q414 AND symb_decoder(16#10#)) OR
 					(reg_q414 AND symb_decoder(16#80#)) OR
 					(reg_q414 AND symb_decoder(16#9e#)) OR
 					(reg_q414 AND symb_decoder(16#ce#)) OR
 					(reg_q414 AND symb_decoder(16#ea#)) OR
 					(reg_q414 AND symb_decoder(16#d9#)) OR
 					(reg_q414 AND symb_decoder(16#39#)) OR
 					(reg_q414 AND symb_decoder(16#6f#)) OR
 					(reg_q414 AND symb_decoder(16#40#)) OR
 					(reg_q414 AND symb_decoder(16#b7#)) OR
 					(reg_q414 AND symb_decoder(16#31#)) OR
 					(reg_q414 AND symb_decoder(16#90#)) OR
 					(reg_q414 AND symb_decoder(16#bd#)) OR
 					(reg_q414 AND symb_decoder(16#b9#)) OR
 					(reg_q414 AND symb_decoder(16#99#)) OR
 					(reg_q414 AND symb_decoder(16#8f#)) OR
 					(reg_q414 AND symb_decoder(16#62#)) OR
 					(reg_q414 AND symb_decoder(16#1b#)) OR
 					(reg_q414 AND symb_decoder(16#35#)) OR
 					(reg_q414 AND symb_decoder(16#e8#)) OR
 					(reg_q414 AND symb_decoder(16#e1#)) OR
 					(reg_q414 AND symb_decoder(16#52#)) OR
 					(reg_q414 AND symb_decoder(16#05#)) OR
 					(reg_q414 AND symb_decoder(16#a3#)) OR
 					(reg_q414 AND symb_decoder(16#7b#)) OR
 					(reg_q414 AND symb_decoder(16#3c#)) OR
 					(reg_q414 AND symb_decoder(16#f9#)) OR
 					(reg_q414 AND symb_decoder(16#bf#)) OR
 					(reg_q414 AND symb_decoder(16#03#)) OR
 					(reg_q414 AND symb_decoder(16#67#)) OR
 					(reg_q414 AND symb_decoder(16#1e#)) OR
 					(reg_q414 AND symb_decoder(16#d1#)) OR
 					(reg_q414 AND symb_decoder(16#58#)) OR
 					(reg_q414 AND symb_decoder(16#98#)) OR
 					(reg_q414 AND symb_decoder(16#cb#)) OR
 					(reg_q414 AND symb_decoder(16#d3#)) OR
 					(reg_q414 AND symb_decoder(16#27#)) OR
 					(reg_q414 AND symb_decoder(16#a8#)) OR
 					(reg_q414 AND symb_decoder(16#56#)) OR
 					(reg_q414 AND symb_decoder(16#f0#)) OR
 					(reg_q414 AND symb_decoder(16#b6#)) OR
 					(reg_q414 AND symb_decoder(16#f3#)) OR
 					(reg_q414 AND symb_decoder(16#08#)) OR
 					(reg_q414 AND symb_decoder(16#60#)) OR
 					(reg_q414 AND symb_decoder(16#18#)) OR
 					(reg_q414 AND symb_decoder(16#dc#)) OR
 					(reg_q414 AND symb_decoder(16#19#)) OR
 					(reg_q414 AND symb_decoder(16#9c#)) OR
 					(reg_q414 AND symb_decoder(16#28#)) OR
 					(reg_q414 AND symb_decoder(16#e3#)) OR
 					(reg_q414 AND symb_decoder(16#01#)) OR
 					(reg_q414 AND symb_decoder(16#3f#)) OR
 					(reg_q414 AND symb_decoder(16#a2#)) OR
 					(reg_q414 AND symb_decoder(16#51#)) OR
 					(reg_q414 AND symb_decoder(16#3b#)) OR
 					(reg_q414 AND symb_decoder(16#2e#)) OR
 					(reg_q414 AND symb_decoder(16#d6#)) OR
 					(reg_q414 AND symb_decoder(16#ac#)) OR
 					(reg_q414 AND symb_decoder(16#c0#)) OR
 					(reg_q414 AND symb_decoder(16#92#)) OR
 					(reg_q414 AND symb_decoder(16#5c#)) OR
 					(reg_q414 AND symb_decoder(16#00#)) OR
 					(reg_q414 AND symb_decoder(16#76#)) OR
 					(reg_q414 AND symb_decoder(16#23#)) OR
 					(reg_q414 AND symb_decoder(16#6b#)) OR
 					(reg_q414 AND symb_decoder(16#2c#));
reg_q414_init <= '0' ;
	p_reg_q414: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q414 <= reg_q414_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q414 <= reg_q414_init;
        else
          reg_q414 <= reg_q414_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2252_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2252 AND symb_decoder(16#63#)) OR
 					(reg_q2252 AND symb_decoder(16#43#)) OR
 					(reg_q2252 AND symb_decoder(16#d2#)) OR
 					(reg_q2252 AND symb_decoder(16#ab#)) OR
 					(reg_q2252 AND symb_decoder(16#a6#)) OR
 					(reg_q2252 AND symb_decoder(16#90#)) OR
 					(reg_q2252 AND symb_decoder(16#0a#)) OR
 					(reg_q2252 AND symb_decoder(16#9e#)) OR
 					(reg_q2252 AND symb_decoder(16#86#)) OR
 					(reg_q2252 AND symb_decoder(16#24#)) OR
 					(reg_q2252 AND symb_decoder(16#ec#)) OR
 					(reg_q2252 AND symb_decoder(16#b0#)) OR
 					(reg_q2252 AND symb_decoder(16#7d#)) OR
 					(reg_q2252 AND symb_decoder(16#1a#)) OR
 					(reg_q2252 AND symb_decoder(16#a3#)) OR
 					(reg_q2252 AND symb_decoder(16#93#)) OR
 					(reg_q2252 AND symb_decoder(16#70#)) OR
 					(reg_q2252 AND symb_decoder(16#d9#)) OR
 					(reg_q2252 AND symb_decoder(16#e5#)) OR
 					(reg_q2252 AND symb_decoder(16#14#)) OR
 					(reg_q2252 AND symb_decoder(16#33#)) OR
 					(reg_q2252 AND symb_decoder(16#9c#)) OR
 					(reg_q2252 AND symb_decoder(16#5e#)) OR
 					(reg_q2252 AND symb_decoder(16#42#)) OR
 					(reg_q2252 AND symb_decoder(16#f5#)) OR
 					(reg_q2252 AND symb_decoder(16#b4#)) OR
 					(reg_q2252 AND symb_decoder(16#64#)) OR
 					(reg_q2252 AND symb_decoder(16#c1#)) OR
 					(reg_q2252 AND symb_decoder(16#f1#)) OR
 					(reg_q2252 AND symb_decoder(16#04#)) OR
 					(reg_q2252 AND symb_decoder(16#29#)) OR
 					(reg_q2252 AND symb_decoder(16#27#)) OR
 					(reg_q2252 AND symb_decoder(16#c4#)) OR
 					(reg_q2252 AND symb_decoder(16#74#)) OR
 					(reg_q2252 AND symb_decoder(16#6c#)) OR
 					(reg_q2252 AND symb_decoder(16#d7#)) OR
 					(reg_q2252 AND symb_decoder(16#ef#)) OR
 					(reg_q2252 AND symb_decoder(16#81#)) OR
 					(reg_q2252 AND symb_decoder(16#77#)) OR
 					(reg_q2252 AND symb_decoder(16#cf#)) OR
 					(reg_q2252 AND symb_decoder(16#ca#)) OR
 					(reg_q2252 AND symb_decoder(16#af#)) OR
 					(reg_q2252 AND symb_decoder(16#51#)) OR
 					(reg_q2252 AND symb_decoder(16#22#)) OR
 					(reg_q2252 AND symb_decoder(16#76#)) OR
 					(reg_q2252 AND symb_decoder(16#79#)) OR
 					(reg_q2252 AND symb_decoder(16#b6#)) OR
 					(reg_q2252 AND symb_decoder(16#7c#)) OR
 					(reg_q2252 AND symb_decoder(16#b5#)) OR
 					(reg_q2252 AND symb_decoder(16#39#)) OR
 					(reg_q2252 AND symb_decoder(16#4a#)) OR
 					(reg_q2252 AND symb_decoder(16#34#)) OR
 					(reg_q2252 AND symb_decoder(16#54#)) OR
 					(reg_q2252 AND symb_decoder(16#80#)) OR
 					(reg_q2252 AND symb_decoder(16#41#)) OR
 					(reg_q2252 AND symb_decoder(16#84#)) OR
 					(reg_q2252 AND symb_decoder(16#d6#)) OR
 					(reg_q2252 AND symb_decoder(16#26#)) OR
 					(reg_q2252 AND symb_decoder(16#be#)) OR
 					(reg_q2252 AND symb_decoder(16#05#)) OR
 					(reg_q2252 AND symb_decoder(16#b1#)) OR
 					(reg_q2252 AND symb_decoder(16#3a#)) OR
 					(reg_q2252 AND symb_decoder(16#0e#)) OR
 					(reg_q2252 AND symb_decoder(16#1c#)) OR
 					(reg_q2252 AND symb_decoder(16#e2#)) OR
 					(reg_q2252 AND symb_decoder(16#1d#)) OR
 					(reg_q2252 AND symb_decoder(16#f3#)) OR
 					(reg_q2252 AND symb_decoder(16#a7#)) OR
 					(reg_q2252 AND symb_decoder(16#da#)) OR
 					(reg_q2252 AND symb_decoder(16#2c#)) OR
 					(reg_q2252 AND symb_decoder(16#5a#)) OR
 					(reg_q2252 AND symb_decoder(16#57#)) OR
 					(reg_q2252 AND symb_decoder(16#cb#)) OR
 					(reg_q2252 AND symb_decoder(16#6f#)) OR
 					(reg_q2252 AND symb_decoder(16#f9#)) OR
 					(reg_q2252 AND symb_decoder(16#8a#)) OR
 					(reg_q2252 AND symb_decoder(16#9a#)) OR
 					(reg_q2252 AND symb_decoder(16#7b#)) OR
 					(reg_q2252 AND symb_decoder(16#58#)) OR
 					(reg_q2252 AND symb_decoder(16#10#)) OR
 					(reg_q2252 AND symb_decoder(16#e9#)) OR
 					(reg_q2252 AND symb_decoder(16#e3#)) OR
 					(reg_q2252 AND symb_decoder(16#2a#)) OR
 					(reg_q2252 AND symb_decoder(16#49#)) OR
 					(reg_q2252 AND symb_decoder(16#eb#)) OR
 					(reg_q2252 AND symb_decoder(16#a4#)) OR
 					(reg_q2252 AND symb_decoder(16#7a#)) OR
 					(reg_q2252 AND symb_decoder(16#c3#)) OR
 					(reg_q2252 AND symb_decoder(16#89#)) OR
 					(reg_q2252 AND symb_decoder(16#aa#)) OR
 					(reg_q2252 AND symb_decoder(16#20#)) OR
 					(reg_q2252 AND symb_decoder(16#d5#)) OR
 					(reg_q2252 AND symb_decoder(16#5c#)) OR
 					(reg_q2252 AND symb_decoder(16#3c#)) OR
 					(reg_q2252 AND symb_decoder(16#0f#)) OR
 					(reg_q2252 AND symb_decoder(16#23#)) OR
 					(reg_q2252 AND symb_decoder(16#c8#)) OR
 					(reg_q2252 AND symb_decoder(16#0d#)) OR
 					(reg_q2252 AND symb_decoder(16#07#)) OR
 					(reg_q2252 AND symb_decoder(16#7f#)) OR
 					(reg_q2252 AND symb_decoder(16#c0#)) OR
 					(reg_q2252 AND symb_decoder(16#b3#)) OR
 					(reg_q2252 AND symb_decoder(16#69#)) OR
 					(reg_q2252 AND symb_decoder(16#08#)) OR
 					(reg_q2252 AND symb_decoder(16#4f#)) OR
 					(reg_q2252 AND symb_decoder(16#a5#)) OR
 					(reg_q2252 AND symb_decoder(16#75#)) OR
 					(reg_q2252 AND symb_decoder(16#56#)) OR
 					(reg_q2252 AND symb_decoder(16#dd#)) OR
 					(reg_q2252 AND symb_decoder(16#8e#)) OR
 					(reg_q2252 AND symb_decoder(16#11#)) OR
 					(reg_q2252 AND symb_decoder(16#28#)) OR
 					(reg_q2252 AND symb_decoder(16#e0#)) OR
 					(reg_q2252 AND symb_decoder(16#12#)) OR
 					(reg_q2252 AND symb_decoder(16#9f#)) OR
 					(reg_q2252 AND symb_decoder(16#ac#)) OR
 					(reg_q2252 AND symb_decoder(16#de#)) OR
 					(reg_q2252 AND symb_decoder(16#3d#)) OR
 					(reg_q2252 AND symb_decoder(16#37#)) OR
 					(reg_q2252 AND symb_decoder(16#62#)) OR
 					(reg_q2252 AND symb_decoder(16#2b#)) OR
 					(reg_q2252 AND symb_decoder(16#f7#)) OR
 					(reg_q2252 AND symb_decoder(16#ff#)) OR
 					(reg_q2252 AND symb_decoder(16#96#)) OR
 					(reg_q2252 AND symb_decoder(16#53#)) OR
 					(reg_q2252 AND symb_decoder(16#bb#)) OR
 					(reg_q2252 AND symb_decoder(16#95#)) OR
 					(reg_q2252 AND symb_decoder(16#e7#)) OR
 					(reg_q2252 AND symb_decoder(16#fd#)) OR
 					(reg_q2252 AND symb_decoder(16#8d#)) OR
 					(reg_q2252 AND symb_decoder(16#87#)) OR
 					(reg_q2252 AND symb_decoder(16#a8#)) OR
 					(reg_q2252 AND symb_decoder(16#85#)) OR
 					(reg_q2252 AND symb_decoder(16#60#)) OR
 					(reg_q2252 AND symb_decoder(16#3f#)) OR
 					(reg_q2252 AND symb_decoder(16#c7#)) OR
 					(reg_q2252 AND symb_decoder(16#f0#)) OR
 					(reg_q2252 AND symb_decoder(16#2e#)) OR
 					(reg_q2252 AND symb_decoder(16#c2#)) OR
 					(reg_q2252 AND symb_decoder(16#cd#)) OR
 					(reg_q2252 AND symb_decoder(16#4c#)) OR
 					(reg_q2252 AND symb_decoder(16#ce#)) OR
 					(reg_q2252 AND symb_decoder(16#94#)) OR
 					(reg_q2252 AND symb_decoder(16#fe#)) OR
 					(reg_q2252 AND symb_decoder(16#52#)) OR
 					(reg_q2252 AND symb_decoder(16#6d#)) OR
 					(reg_q2252 AND symb_decoder(16#19#)) OR
 					(reg_q2252 AND symb_decoder(16#1b#)) OR
 					(reg_q2252 AND symb_decoder(16#15#)) OR
 					(reg_q2252 AND symb_decoder(16#1e#)) OR
 					(reg_q2252 AND symb_decoder(16#4d#)) OR
 					(reg_q2252 AND symb_decoder(16#ba#)) OR
 					(reg_q2252 AND symb_decoder(16#d8#)) OR
 					(reg_q2252 AND symb_decoder(16#a9#)) OR
 					(reg_q2252 AND symb_decoder(16#fc#)) OR
 					(reg_q2252 AND symb_decoder(16#21#)) OR
 					(reg_q2252 AND symb_decoder(16#d4#)) OR
 					(reg_q2252 AND symb_decoder(16#b7#)) OR
 					(reg_q2252 AND symb_decoder(16#09#)) OR
 					(reg_q2252 AND symb_decoder(16#6e#)) OR
 					(reg_q2252 AND symb_decoder(16#dc#)) OR
 					(reg_q2252 AND symb_decoder(16#d0#)) OR
 					(reg_q2252 AND symb_decoder(16#d1#)) OR
 					(reg_q2252 AND symb_decoder(16#bc#)) OR
 					(reg_q2252 AND symb_decoder(16#ea#)) OR
 					(reg_q2252 AND symb_decoder(16#3b#)) OR
 					(reg_q2252 AND symb_decoder(16#d3#)) OR
 					(reg_q2252 AND symb_decoder(16#bf#)) OR
 					(reg_q2252 AND symb_decoder(16#66#)) OR
 					(reg_q2252 AND symb_decoder(16#b2#)) OR
 					(reg_q2252 AND symb_decoder(16#2f#)) OR
 					(reg_q2252 AND symb_decoder(16#6b#)) OR
 					(reg_q2252 AND symb_decoder(16#47#)) OR
 					(reg_q2252 AND symb_decoder(16#8f#)) OR
 					(reg_q2252 AND symb_decoder(16#ad#)) OR
 					(reg_q2252 AND symb_decoder(16#17#)) OR
 					(reg_q2252 AND symb_decoder(16#8b#)) OR
 					(reg_q2252 AND symb_decoder(16#71#)) OR
 					(reg_q2252 AND symb_decoder(16#8c#)) OR
 					(reg_q2252 AND symb_decoder(16#55#)) OR
 					(reg_q2252 AND symb_decoder(16#a2#)) OR
 					(reg_q2252 AND symb_decoder(16#83#)) OR
 					(reg_q2252 AND symb_decoder(16#5b#)) OR
 					(reg_q2252 AND symb_decoder(16#cc#)) OR
 					(reg_q2252 AND symb_decoder(16#b9#)) OR
 					(reg_q2252 AND symb_decoder(16#ed#)) OR
 					(reg_q2252 AND symb_decoder(16#48#)) OR
 					(reg_q2252 AND symb_decoder(16#38#)) OR
 					(reg_q2252 AND symb_decoder(16#7e#)) OR
 					(reg_q2252 AND symb_decoder(16#9b#)) OR
 					(reg_q2252 AND symb_decoder(16#0c#)) OR
 					(reg_q2252 AND symb_decoder(16#2d#)) OR
 					(reg_q2252 AND symb_decoder(16#db#)) OR
 					(reg_q2252 AND symb_decoder(16#78#)) OR
 					(reg_q2252 AND symb_decoder(16#ae#)) OR
 					(reg_q2252 AND symb_decoder(16#44#)) OR
 					(reg_q2252 AND symb_decoder(16#6a#)) OR
 					(reg_q2252 AND symb_decoder(16#68#)) OR
 					(reg_q2252 AND symb_decoder(16#98#)) OR
 					(reg_q2252 AND symb_decoder(16#88#)) OR
 					(reg_q2252 AND symb_decoder(16#97#)) OR
 					(reg_q2252 AND symb_decoder(16#00#)) OR
 					(reg_q2252 AND symb_decoder(16#67#)) OR
 					(reg_q2252 AND symb_decoder(16#31#)) OR
 					(reg_q2252 AND symb_decoder(16#16#)) OR
 					(reg_q2252 AND symb_decoder(16#45#)) OR
 					(reg_q2252 AND symb_decoder(16#5d#)) OR
 					(reg_q2252 AND symb_decoder(16#40#)) OR
 					(reg_q2252 AND symb_decoder(16#a0#)) OR
 					(reg_q2252 AND symb_decoder(16#e1#)) OR
 					(reg_q2252 AND symb_decoder(16#25#)) OR
 					(reg_q2252 AND symb_decoder(16#b8#)) OR
 					(reg_q2252 AND symb_decoder(16#46#)) OR
 					(reg_q2252 AND symb_decoder(16#99#)) OR
 					(reg_q2252 AND symb_decoder(16#9d#)) OR
 					(reg_q2252 AND symb_decoder(16#4e#)) OR
 					(reg_q2252 AND symb_decoder(16#36#)) OR
 					(reg_q2252 AND symb_decoder(16#50#)) OR
 					(reg_q2252 AND symb_decoder(16#01#)) OR
 					(reg_q2252 AND symb_decoder(16#f8#)) OR
 					(reg_q2252 AND symb_decoder(16#df#)) OR
 					(reg_q2252 AND symb_decoder(16#06#)) OR
 					(reg_q2252 AND symb_decoder(16#c5#)) OR
 					(reg_q2252 AND symb_decoder(16#5f#)) OR
 					(reg_q2252 AND symb_decoder(16#f4#)) OR
 					(reg_q2252 AND symb_decoder(16#3e#)) OR
 					(reg_q2252 AND symb_decoder(16#ee#)) OR
 					(reg_q2252 AND symb_decoder(16#f2#)) OR
 					(reg_q2252 AND symb_decoder(16#30#)) OR
 					(reg_q2252 AND symb_decoder(16#73#)) OR
 					(reg_q2252 AND symb_decoder(16#59#)) OR
 					(reg_q2252 AND symb_decoder(16#03#)) OR
 					(reg_q2252 AND symb_decoder(16#fa#)) OR
 					(reg_q2252 AND symb_decoder(16#a1#)) OR
 					(reg_q2252 AND symb_decoder(16#72#)) OR
 					(reg_q2252 AND symb_decoder(16#92#)) OR
 					(reg_q2252 AND symb_decoder(16#82#)) OR
 					(reg_q2252 AND symb_decoder(16#13#)) OR
 					(reg_q2252 AND symb_decoder(16#0b#)) OR
 					(reg_q2252 AND symb_decoder(16#f6#)) OR
 					(reg_q2252 AND symb_decoder(16#1f#)) OR
 					(reg_q2252 AND symb_decoder(16#e4#)) OR
 					(reg_q2252 AND symb_decoder(16#32#)) OR
 					(reg_q2252 AND symb_decoder(16#fb#)) OR
 					(reg_q2252 AND symb_decoder(16#65#)) OR
 					(reg_q2252 AND symb_decoder(16#e8#)) OR
 					(reg_q2252 AND symb_decoder(16#c9#)) OR
 					(reg_q2252 AND symb_decoder(16#bd#)) OR
 					(reg_q2252 AND symb_decoder(16#18#)) OR
 					(reg_q2252 AND symb_decoder(16#c6#)) OR
 					(reg_q2252 AND symb_decoder(16#02#)) OR
 					(reg_q2252 AND symb_decoder(16#e6#)) OR
 					(reg_q2252 AND symb_decoder(16#61#)) OR
 					(reg_q2252 AND symb_decoder(16#35#)) OR
 					(reg_q2252 AND symb_decoder(16#91#)) OR
 					(reg_q2252 AND symb_decoder(16#4b#));
reg_q2252_init <= '0' ;
	p_reg_q2252: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2252 <= reg_q2252_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2252 <= reg_q2252_init;
        else
          reg_q2252 <= reg_q2252_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q913_in <= (reg_q911 AND symb_decoder(16#74#)) OR
 					(reg_q911 AND symb_decoder(16#54#));
reg_q913_init <= '0' ;
	p_reg_q913: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q913 <= reg_q913_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q913 <= reg_q913_init;
        else
          reg_q913 <= reg_q913_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q915_in <= (reg_q913 AND symb_decoder(16#20#)) OR
 					(reg_q913 AND symb_decoder(16#0c#)) OR
 					(reg_q913 AND symb_decoder(16#0d#)) OR
 					(reg_q913 AND symb_decoder(16#0a#)) OR
 					(reg_q913 AND symb_decoder(16#09#)) OR
 					(reg_q915 AND symb_decoder(16#20#)) OR
 					(reg_q915 AND symb_decoder(16#0d#)) OR
 					(reg_q915 AND symb_decoder(16#0a#)) OR
 					(reg_q915 AND symb_decoder(16#09#)) OR
 					(reg_q915 AND symb_decoder(16#0c#));
reg_q915_init <= '0' ;
	p_reg_q915: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q915 <= reg_q915_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q915 <= reg_q915_init;
        else
          reg_q915 <= reg_q915_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2192_in <= (reg_q2190 AND symb_decoder(16#6c#)) OR
 					(reg_q2190 AND symb_decoder(16#4c#));
reg_q2192_init <= '0' ;
	p_reg_q2192: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2192 <= reg_q2192_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2192 <= reg_q2192_init;
        else
          reg_q2192 <= reg_q2192_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2194_in <= (reg_q2192 AND symb_decoder(16#0d#)) OR
 					(reg_q2192 AND symb_decoder(16#0c#)) OR
 					(reg_q2192 AND symb_decoder(16#09#)) OR
 					(reg_q2192 AND symb_decoder(16#20#)) OR
 					(reg_q2192 AND symb_decoder(16#0a#)) OR
 					(reg_q2194 AND symb_decoder(16#0d#)) OR
 					(reg_q2194 AND symb_decoder(16#09#)) OR
 					(reg_q2194 AND symb_decoder(16#0a#)) OR
 					(reg_q2194 AND symb_decoder(16#0c#)) OR
 					(reg_q2194 AND symb_decoder(16#20#));
reg_q2194_init <= '0' ;
	p_reg_q2194: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2194 <= reg_q2194_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2194 <= reg_q2194_init;
        else
          reg_q2194 <= reg_q2194_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q680_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q680 AND symb_decoder(16#d0#)) OR
 					(reg_q680 AND symb_decoder(16#3c#)) OR
 					(reg_q680 AND symb_decoder(16#95#)) OR
 					(reg_q680 AND symb_decoder(16#ee#)) OR
 					(reg_q680 AND symb_decoder(16#9a#)) OR
 					(reg_q680 AND symb_decoder(16#c4#)) OR
 					(reg_q680 AND symb_decoder(16#33#)) OR
 					(reg_q680 AND symb_decoder(16#03#)) OR
 					(reg_q680 AND symb_decoder(16#f8#)) OR
 					(reg_q680 AND symb_decoder(16#11#)) OR
 					(reg_q680 AND symb_decoder(16#26#)) OR
 					(reg_q680 AND symb_decoder(16#f0#)) OR
 					(reg_q680 AND symb_decoder(16#1c#)) OR
 					(reg_q680 AND symb_decoder(16#ae#)) OR
 					(reg_q680 AND symb_decoder(16#7e#)) OR
 					(reg_q680 AND symb_decoder(16#b1#)) OR
 					(reg_q680 AND symb_decoder(16#46#)) OR
 					(reg_q680 AND symb_decoder(16#8c#)) OR
 					(reg_q680 AND symb_decoder(16#ad#)) OR
 					(reg_q680 AND symb_decoder(16#32#)) OR
 					(reg_q680 AND symb_decoder(16#77#)) OR
 					(reg_q680 AND symb_decoder(16#d8#)) OR
 					(reg_q680 AND symb_decoder(16#bb#)) OR
 					(reg_q680 AND symb_decoder(16#e5#)) OR
 					(reg_q680 AND symb_decoder(16#17#)) OR
 					(reg_q680 AND symb_decoder(16#15#)) OR
 					(reg_q680 AND symb_decoder(16#0b#)) OR
 					(reg_q680 AND symb_decoder(16#3e#)) OR
 					(reg_q680 AND symb_decoder(16#ef#)) OR
 					(reg_q680 AND symb_decoder(16#86#)) OR
 					(reg_q680 AND symb_decoder(16#34#)) OR
 					(reg_q680 AND symb_decoder(16#1e#)) OR
 					(reg_q680 AND symb_decoder(16#cd#)) OR
 					(reg_q680 AND symb_decoder(16#0a#)) OR
 					(reg_q680 AND symb_decoder(16#48#)) OR
 					(reg_q680 AND symb_decoder(16#fa#)) OR
 					(reg_q680 AND symb_decoder(16#2c#)) OR
 					(reg_q680 AND symb_decoder(16#81#)) OR
 					(reg_q680 AND symb_decoder(16#55#)) OR
 					(reg_q680 AND symb_decoder(16#66#)) OR
 					(reg_q680 AND symb_decoder(16#35#)) OR
 					(reg_q680 AND symb_decoder(16#e0#)) OR
 					(reg_q680 AND symb_decoder(16#f7#)) OR
 					(reg_q680 AND symb_decoder(16#60#)) OR
 					(reg_q680 AND symb_decoder(16#73#)) OR
 					(reg_q680 AND symb_decoder(16#a2#)) OR
 					(reg_q680 AND symb_decoder(16#c0#)) OR
 					(reg_q680 AND symb_decoder(16#04#)) OR
 					(reg_q680 AND symb_decoder(16#e9#)) OR
 					(reg_q680 AND symb_decoder(16#12#)) OR
 					(reg_q680 AND symb_decoder(16#1d#)) OR
 					(reg_q680 AND symb_decoder(16#19#)) OR
 					(reg_q680 AND symb_decoder(16#75#)) OR
 					(reg_q680 AND symb_decoder(16#2b#)) OR
 					(reg_q680 AND symb_decoder(16#38#)) OR
 					(reg_q680 AND symb_decoder(16#e4#)) OR
 					(reg_q680 AND symb_decoder(16#de#)) OR
 					(reg_q680 AND symb_decoder(16#05#)) OR
 					(reg_q680 AND symb_decoder(16#5e#)) OR
 					(reg_q680 AND symb_decoder(16#f2#)) OR
 					(reg_q680 AND symb_decoder(16#a4#)) OR
 					(reg_q680 AND symb_decoder(16#e1#)) OR
 					(reg_q680 AND symb_decoder(16#4b#)) OR
 					(reg_q680 AND symb_decoder(16#e2#)) OR
 					(reg_q680 AND symb_decoder(16#e8#)) OR
 					(reg_q680 AND symb_decoder(16#3b#)) OR
 					(reg_q680 AND symb_decoder(16#07#)) OR
 					(reg_q680 AND symb_decoder(16#f9#)) OR
 					(reg_q680 AND symb_decoder(16#b2#)) OR
 					(reg_q680 AND symb_decoder(16#80#)) OR
 					(reg_q680 AND symb_decoder(16#5a#)) OR
 					(reg_q680 AND symb_decoder(16#9b#)) OR
 					(reg_q680 AND symb_decoder(16#50#)) OR
 					(reg_q680 AND symb_decoder(16#e7#)) OR
 					(reg_q680 AND symb_decoder(16#02#)) OR
 					(reg_q680 AND symb_decoder(16#7b#)) OR
 					(reg_q680 AND symb_decoder(16#e3#)) OR
 					(reg_q680 AND symb_decoder(16#43#)) OR
 					(reg_q680 AND symb_decoder(16#ca#)) OR
 					(reg_q680 AND symb_decoder(16#21#)) OR
 					(reg_q680 AND symb_decoder(16#8b#)) OR
 					(reg_q680 AND symb_decoder(16#c7#)) OR
 					(reg_q680 AND symb_decoder(16#f3#)) OR
 					(reg_q680 AND symb_decoder(16#0d#)) OR
 					(reg_q680 AND symb_decoder(16#3f#)) OR
 					(reg_q680 AND symb_decoder(16#5c#)) OR
 					(reg_q680 AND symb_decoder(16#20#)) OR
 					(reg_q680 AND symb_decoder(16#1b#)) OR
 					(reg_q680 AND symb_decoder(16#45#)) OR
 					(reg_q680 AND symb_decoder(16#4a#)) OR
 					(reg_q680 AND symb_decoder(16#cb#)) OR
 					(reg_q680 AND symb_decoder(16#31#)) OR
 					(reg_q680 AND symb_decoder(16#f5#)) OR
 					(reg_q680 AND symb_decoder(16#da#)) OR
 					(reg_q680 AND symb_decoder(16#29#)) OR
 					(reg_q680 AND symb_decoder(16#b8#)) OR
 					(reg_q680 AND symb_decoder(16#be#)) OR
 					(reg_q680 AND symb_decoder(16#2f#)) OR
 					(reg_q680 AND symb_decoder(16#d5#)) OR
 					(reg_q680 AND symb_decoder(16#28#)) OR
 					(reg_q680 AND symb_decoder(16#c2#)) OR
 					(reg_q680 AND symb_decoder(16#d6#)) OR
 					(reg_q680 AND symb_decoder(16#e6#)) OR
 					(reg_q680 AND symb_decoder(16#4d#)) OR
 					(reg_q680 AND symb_decoder(16#db#)) OR
 					(reg_q680 AND symb_decoder(16#94#)) OR
 					(reg_q680 AND symb_decoder(16#37#)) OR
 					(reg_q680 AND symb_decoder(16#76#)) OR
 					(reg_q680 AND symb_decoder(16#9e#)) OR
 					(reg_q680 AND symb_decoder(16#99#)) OR
 					(reg_q680 AND symb_decoder(16#8e#)) OR
 					(reg_q680 AND symb_decoder(16#fd#)) OR
 					(reg_q680 AND symb_decoder(16#b3#)) OR
 					(reg_q680 AND symb_decoder(16#ac#)) OR
 					(reg_q680 AND symb_decoder(16#6d#)) OR
 					(reg_q680 AND symb_decoder(16#a8#)) OR
 					(reg_q680 AND symb_decoder(16#3a#)) OR
 					(reg_q680 AND symb_decoder(16#a0#)) OR
 					(reg_q680 AND symb_decoder(16#ed#)) OR
 					(reg_q680 AND symb_decoder(16#92#)) OR
 					(reg_q680 AND symb_decoder(16#eb#)) OR
 					(reg_q680 AND symb_decoder(16#72#)) OR
 					(reg_q680 AND symb_decoder(16#d4#)) OR
 					(reg_q680 AND symb_decoder(16#7d#)) OR
 					(reg_q680 AND symb_decoder(16#c3#)) OR
 					(reg_q680 AND symb_decoder(16#6a#)) OR
 					(reg_q680 AND symb_decoder(16#c8#)) OR
 					(reg_q680 AND symb_decoder(16#4f#)) OR
 					(reg_q680 AND symb_decoder(16#af#)) OR
 					(reg_q680 AND symb_decoder(16#83#)) OR
 					(reg_q680 AND symb_decoder(16#24#)) OR
 					(reg_q680 AND symb_decoder(16#b9#)) OR
 					(reg_q680 AND symb_decoder(16#fe#)) OR
 					(reg_q680 AND symb_decoder(16#cc#)) OR
 					(reg_q680 AND symb_decoder(16#d1#)) OR
 					(reg_q680 AND symb_decoder(16#2a#)) OR
 					(reg_q680 AND symb_decoder(16#2d#)) OR
 					(reg_q680 AND symb_decoder(16#8a#)) OR
 					(reg_q680 AND symb_decoder(16#09#)) OR
 					(reg_q680 AND symb_decoder(16#0f#)) OR
 					(reg_q680 AND symb_decoder(16#c5#)) OR
 					(reg_q680 AND symb_decoder(16#89#)) OR
 					(reg_q680 AND symb_decoder(16#67#)) OR
 					(reg_q680 AND symb_decoder(16#01#)) OR
 					(reg_q680 AND symb_decoder(16#53#)) OR
 					(reg_q680 AND symb_decoder(16#82#)) OR
 					(reg_q680 AND symb_decoder(16#25#)) OR
 					(reg_q680 AND symb_decoder(16#47#)) OR
 					(reg_q680 AND symb_decoder(16#6f#)) OR
 					(reg_q680 AND symb_decoder(16#ce#)) OR
 					(reg_q680 AND symb_decoder(16#a5#)) OR
 					(reg_q680 AND symb_decoder(16#90#)) OR
 					(reg_q680 AND symb_decoder(16#df#)) OR
 					(reg_q680 AND symb_decoder(16#06#)) OR
 					(reg_q680 AND symb_decoder(16#74#)) OR
 					(reg_q680 AND symb_decoder(16#5f#)) OR
 					(reg_q680 AND symb_decoder(16#b7#)) OR
 					(reg_q680 AND symb_decoder(16#52#)) OR
 					(reg_q680 AND symb_decoder(16#a6#)) OR
 					(reg_q680 AND symb_decoder(16#63#)) OR
 					(reg_q680 AND symb_decoder(16#ff#)) OR
 					(reg_q680 AND symb_decoder(16#08#)) OR
 					(reg_q680 AND symb_decoder(16#8f#)) OR
 					(reg_q680 AND symb_decoder(16#51#)) OR
 					(reg_q680 AND symb_decoder(16#b6#)) OR
 					(reg_q680 AND symb_decoder(16#6b#)) OR
 					(reg_q680 AND symb_decoder(16#14#)) OR
 					(reg_q680 AND symb_decoder(16#97#)) OR
 					(reg_q680 AND symb_decoder(16#9f#)) OR
 					(reg_q680 AND symb_decoder(16#7a#)) OR
 					(reg_q680 AND symb_decoder(16#27#)) OR
 					(reg_q680 AND symb_decoder(16#1f#)) OR
 					(reg_q680 AND symb_decoder(16#62#)) OR
 					(reg_q680 AND symb_decoder(16#61#)) OR
 					(reg_q680 AND symb_decoder(16#64#)) OR
 					(reg_q680 AND symb_decoder(16#9d#)) OR
 					(reg_q680 AND symb_decoder(16#58#)) OR
 					(reg_q680 AND symb_decoder(16#fb#)) OR
 					(reg_q680 AND symb_decoder(16#c9#)) OR
 					(reg_q680 AND symb_decoder(16#49#)) OR
 					(reg_q680 AND symb_decoder(16#18#)) OR
 					(reg_q680 AND symb_decoder(16#dd#)) OR
 					(reg_q680 AND symb_decoder(16#c6#)) OR
 					(reg_q680 AND symb_decoder(16#87#)) OR
 					(reg_q680 AND symb_decoder(16#57#)) OR
 					(reg_q680 AND symb_decoder(16#cf#)) OR
 					(reg_q680 AND symb_decoder(16#96#)) OR
 					(reg_q680 AND symb_decoder(16#7f#)) OR
 					(reg_q680 AND symb_decoder(16#0c#)) OR
 					(reg_q680 AND symb_decoder(16#d9#)) OR
 					(reg_q680 AND symb_decoder(16#6e#)) OR
 					(reg_q680 AND symb_decoder(16#93#)) OR
 					(reg_q680 AND symb_decoder(16#69#)) OR
 					(reg_q680 AND symb_decoder(16#4c#)) OR
 					(reg_q680 AND symb_decoder(16#ea#)) OR
 					(reg_q680 AND symb_decoder(16#54#)) OR
 					(reg_q680 AND symb_decoder(16#23#)) OR
 					(reg_q680 AND symb_decoder(16#dc#)) OR
 					(reg_q680 AND symb_decoder(16#16#)) OR
 					(reg_q680 AND symb_decoder(16#ab#)) OR
 					(reg_q680 AND symb_decoder(16#44#)) OR
 					(reg_q680 AND symb_decoder(16#7c#)) OR
 					(reg_q680 AND symb_decoder(16#39#)) OR
 					(reg_q680 AND symb_decoder(16#2e#)) OR
 					(reg_q680 AND symb_decoder(16#71#)) OR
 					(reg_q680 AND symb_decoder(16#bd#)) OR
 					(reg_q680 AND symb_decoder(16#10#)) OR
 					(reg_q680 AND symb_decoder(16#5d#)) OR
 					(reg_q680 AND symb_decoder(16#30#)) OR
 					(reg_q680 AND symb_decoder(16#36#)) OR
 					(reg_q680 AND symb_decoder(16#fc#)) OR
 					(reg_q680 AND symb_decoder(16#b0#)) OR
 					(reg_q680 AND symb_decoder(16#a9#)) OR
 					(reg_q680 AND symb_decoder(16#ba#)) OR
 					(reg_q680 AND symb_decoder(16#b5#)) OR
 					(reg_q680 AND symb_decoder(16#a1#)) OR
 					(reg_q680 AND symb_decoder(16#ec#)) OR
 					(reg_q680 AND symb_decoder(16#d2#)) OR
 					(reg_q680 AND symb_decoder(16#88#)) OR
 					(reg_q680 AND symb_decoder(16#f1#)) OR
 					(reg_q680 AND symb_decoder(16#b4#)) OR
 					(reg_q680 AND symb_decoder(16#aa#)) OR
 					(reg_q680 AND symb_decoder(16#d7#)) OR
 					(reg_q680 AND symb_decoder(16#1a#)) OR
 					(reg_q680 AND symb_decoder(16#78#)) OR
 					(reg_q680 AND symb_decoder(16#00#)) OR
 					(reg_q680 AND symb_decoder(16#79#)) OR
 					(reg_q680 AND symb_decoder(16#13#)) OR
 					(reg_q680 AND symb_decoder(16#91#)) OR
 					(reg_q680 AND symb_decoder(16#56#)) OR
 					(reg_q680 AND symb_decoder(16#22#)) OR
 					(reg_q680 AND symb_decoder(16#4e#)) OR
 					(reg_q680 AND symb_decoder(16#98#)) OR
 					(reg_q680 AND symb_decoder(16#9c#)) OR
 					(reg_q680 AND symb_decoder(16#5b#)) OR
 					(reg_q680 AND symb_decoder(16#85#)) OR
 					(reg_q680 AND symb_decoder(16#bf#)) OR
 					(reg_q680 AND symb_decoder(16#6c#)) OR
 					(reg_q680 AND symb_decoder(16#65#)) OR
 					(reg_q680 AND symb_decoder(16#3d#)) OR
 					(reg_q680 AND symb_decoder(16#70#)) OR
 					(reg_q680 AND symb_decoder(16#40#)) OR
 					(reg_q680 AND symb_decoder(16#f6#)) OR
 					(reg_q680 AND symb_decoder(16#41#)) OR
 					(reg_q680 AND symb_decoder(16#0e#)) OR
 					(reg_q680 AND symb_decoder(16#59#)) OR
 					(reg_q680 AND symb_decoder(16#68#)) OR
 					(reg_q680 AND symb_decoder(16#a3#)) OR
 					(reg_q680 AND symb_decoder(16#f4#)) OR
 					(reg_q680 AND symb_decoder(16#8d#)) OR
 					(reg_q680 AND symb_decoder(16#84#)) OR
 					(reg_q680 AND symb_decoder(16#bc#)) OR
 					(reg_q680 AND symb_decoder(16#d3#)) OR
 					(reg_q680 AND symb_decoder(16#c1#)) OR
 					(reg_q680 AND symb_decoder(16#42#)) OR
 					(reg_q680 AND symb_decoder(16#a7#));
reg_q680_init <= '0' ;
	p_reg_q680: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q680 <= reg_q680_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q680 <= reg_q680_init;
        else
          reg_q680 <= reg_q680_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q452_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q452 AND symb_decoder(16#10#)) OR
 					(reg_q452 AND symb_decoder(16#4c#)) OR
 					(reg_q452 AND symb_decoder(16#fc#)) OR
 					(reg_q452 AND symb_decoder(16#77#)) OR
 					(reg_q452 AND symb_decoder(16#38#)) OR
 					(reg_q452 AND symb_decoder(16#4d#)) OR
 					(reg_q452 AND symb_decoder(16#0a#)) OR
 					(reg_q452 AND symb_decoder(16#e2#)) OR
 					(reg_q452 AND symb_decoder(16#d4#)) OR
 					(reg_q452 AND symb_decoder(16#b8#)) OR
 					(reg_q452 AND symb_decoder(16#23#)) OR
 					(reg_q452 AND symb_decoder(16#48#)) OR
 					(reg_q452 AND symb_decoder(16#24#)) OR
 					(reg_q452 AND symb_decoder(16#39#)) OR
 					(reg_q452 AND symb_decoder(16#4b#)) OR
 					(reg_q452 AND symb_decoder(16#80#)) OR
 					(reg_q452 AND symb_decoder(16#a7#)) OR
 					(reg_q452 AND symb_decoder(16#f8#)) OR
 					(reg_q452 AND symb_decoder(16#e7#)) OR
 					(reg_q452 AND symb_decoder(16#bb#)) OR
 					(reg_q452 AND symb_decoder(16#1e#)) OR
 					(reg_q452 AND symb_decoder(16#46#)) OR
 					(reg_q452 AND symb_decoder(16#e1#)) OR
 					(reg_q452 AND symb_decoder(16#79#)) OR
 					(reg_q452 AND symb_decoder(16#5e#)) OR
 					(reg_q452 AND symb_decoder(16#96#)) OR
 					(reg_q452 AND symb_decoder(16#a4#)) OR
 					(reg_q452 AND symb_decoder(16#8a#)) OR
 					(reg_q452 AND symb_decoder(16#a1#)) OR
 					(reg_q452 AND symb_decoder(16#c1#)) OR
 					(reg_q452 AND symb_decoder(16#36#)) OR
 					(reg_q452 AND symb_decoder(16#3b#)) OR
 					(reg_q452 AND symb_decoder(16#87#)) OR
 					(reg_q452 AND symb_decoder(16#5a#)) OR
 					(reg_q452 AND symb_decoder(16#94#)) OR
 					(reg_q452 AND symb_decoder(16#7b#)) OR
 					(reg_q452 AND symb_decoder(16#28#)) OR
 					(reg_q452 AND symb_decoder(16#1d#)) OR
 					(reg_q452 AND symb_decoder(16#19#)) OR
 					(reg_q452 AND symb_decoder(16#68#)) OR
 					(reg_q452 AND symb_decoder(16#5f#)) OR
 					(reg_q452 AND symb_decoder(16#6e#)) OR
 					(reg_q452 AND symb_decoder(16#ad#)) OR
 					(reg_q452 AND symb_decoder(16#d7#)) OR
 					(reg_q452 AND symb_decoder(16#b7#)) OR
 					(reg_q452 AND symb_decoder(16#e8#)) OR
 					(reg_q452 AND symb_decoder(16#bf#)) OR
 					(reg_q452 AND symb_decoder(16#42#)) OR
 					(reg_q452 AND symb_decoder(16#08#)) OR
 					(reg_q452 AND symb_decoder(16#4f#)) OR
 					(reg_q452 AND symb_decoder(16#44#)) OR
 					(reg_q452 AND symb_decoder(16#a3#)) OR
 					(reg_q452 AND symb_decoder(16#76#)) OR
 					(reg_q452 AND symb_decoder(16#e6#)) OR
 					(reg_q452 AND symb_decoder(16#21#)) OR
 					(reg_q452 AND symb_decoder(16#05#)) OR
 					(reg_q452 AND symb_decoder(16#fe#)) OR
 					(reg_q452 AND symb_decoder(16#9a#)) OR
 					(reg_q452 AND symb_decoder(16#26#)) OR
 					(reg_q452 AND symb_decoder(16#40#)) OR
 					(reg_q452 AND symb_decoder(16#b9#)) OR
 					(reg_q452 AND symb_decoder(16#e3#)) OR
 					(reg_q452 AND symb_decoder(16#1c#)) OR
 					(reg_q452 AND symb_decoder(16#b1#)) OR
 					(reg_q452 AND symb_decoder(16#ca#)) OR
 					(reg_q452 AND symb_decoder(16#b5#)) OR
 					(reg_q452 AND symb_decoder(16#f4#)) OR
 					(reg_q452 AND symb_decoder(16#a8#)) OR
 					(reg_q452 AND symb_decoder(16#2f#)) OR
 					(reg_q452 AND symb_decoder(16#dc#)) OR
 					(reg_q452 AND symb_decoder(16#1f#)) OR
 					(reg_q452 AND symb_decoder(16#5c#)) OR
 					(reg_q452 AND symb_decoder(16#47#)) OR
 					(reg_q452 AND symb_decoder(16#8e#)) OR
 					(reg_q452 AND symb_decoder(16#43#)) OR
 					(reg_q452 AND symb_decoder(16#b2#)) OR
 					(reg_q452 AND symb_decoder(16#4a#)) OR
 					(reg_q452 AND symb_decoder(16#c8#)) OR
 					(reg_q452 AND symb_decoder(16#13#)) OR
 					(reg_q452 AND symb_decoder(16#17#)) OR
 					(reg_q452 AND symb_decoder(16#2c#)) OR
 					(reg_q452 AND symb_decoder(16#70#)) OR
 					(reg_q452 AND symb_decoder(16#45#)) OR
 					(reg_q452 AND symb_decoder(16#c0#)) OR
 					(reg_q452 AND symb_decoder(16#a2#)) OR
 					(reg_q452 AND symb_decoder(16#b0#)) OR
 					(reg_q452 AND symb_decoder(16#6b#)) OR
 					(reg_q452 AND symb_decoder(16#d6#)) OR
 					(reg_q452 AND symb_decoder(16#a9#)) OR
 					(reg_q452 AND symb_decoder(16#9e#)) OR
 					(reg_q452 AND symb_decoder(16#cf#)) OR
 					(reg_q452 AND symb_decoder(16#ae#)) OR
 					(reg_q452 AND symb_decoder(16#89#)) OR
 					(reg_q452 AND symb_decoder(16#fd#)) OR
 					(reg_q452 AND symb_decoder(16#50#)) OR
 					(reg_q452 AND symb_decoder(16#f9#)) OR
 					(reg_q452 AND symb_decoder(16#fa#)) OR
 					(reg_q452 AND symb_decoder(16#9d#)) OR
 					(reg_q452 AND symb_decoder(16#63#)) OR
 					(reg_q452 AND symb_decoder(16#73#)) OR
 					(reg_q452 AND symb_decoder(16#bd#)) OR
 					(reg_q452 AND symb_decoder(16#db#)) OR
 					(reg_q452 AND symb_decoder(16#ea#)) OR
 					(reg_q452 AND symb_decoder(16#09#)) OR
 					(reg_q452 AND symb_decoder(16#7f#)) OR
 					(reg_q452 AND symb_decoder(16#a5#)) OR
 					(reg_q452 AND symb_decoder(16#cb#)) OR
 					(reg_q452 AND symb_decoder(16#83#)) OR
 					(reg_q452 AND symb_decoder(16#97#)) OR
 					(reg_q452 AND symb_decoder(16#71#)) OR
 					(reg_q452 AND symb_decoder(16#90#)) OR
 					(reg_q452 AND symb_decoder(16#a0#)) OR
 					(reg_q452 AND symb_decoder(16#29#)) OR
 					(reg_q452 AND symb_decoder(16#6d#)) OR
 					(reg_q452 AND symb_decoder(16#00#)) OR
 					(reg_q452 AND symb_decoder(16#07#)) OR
 					(reg_q452 AND symb_decoder(16#59#)) OR
 					(reg_q452 AND symb_decoder(16#56#)) OR
 					(reg_q452 AND symb_decoder(16#1a#)) OR
 					(reg_q452 AND symb_decoder(16#3d#)) OR
 					(reg_q452 AND symb_decoder(16#33#)) OR
 					(reg_q452 AND symb_decoder(16#ec#)) OR
 					(reg_q452 AND symb_decoder(16#c7#)) OR
 					(reg_q452 AND symb_decoder(16#72#)) OR
 					(reg_q452 AND symb_decoder(16#01#)) OR
 					(reg_q452 AND symb_decoder(16#81#)) OR
 					(reg_q452 AND symb_decoder(16#cd#)) OR
 					(reg_q452 AND symb_decoder(16#0e#)) OR
 					(reg_q452 AND symb_decoder(16#df#)) OR
 					(reg_q452 AND symb_decoder(16#6f#)) OR
 					(reg_q452 AND symb_decoder(16#a6#)) OR
 					(reg_q452 AND symb_decoder(16#ee#)) OR
 					(reg_q452 AND symb_decoder(16#75#)) OR
 					(reg_q452 AND symb_decoder(16#88#)) OR
 					(reg_q452 AND symb_decoder(16#41#)) OR
 					(reg_q452 AND symb_decoder(16#66#)) OR
 					(reg_q452 AND symb_decoder(16#0f#)) OR
 					(reg_q452 AND symb_decoder(16#93#)) OR
 					(reg_q452 AND symb_decoder(16#aa#)) OR
 					(reg_q452 AND symb_decoder(16#9c#)) OR
 					(reg_q452 AND symb_decoder(16#b6#)) OR
 					(reg_q452 AND symb_decoder(16#de#)) OR
 					(reg_q452 AND symb_decoder(16#f6#)) OR
 					(reg_q452 AND symb_decoder(16#0b#)) OR
 					(reg_q452 AND symb_decoder(16#22#)) OR
 					(reg_q452 AND symb_decoder(16#7d#)) OR
 					(reg_q452 AND symb_decoder(16#15#)) OR
 					(reg_q452 AND symb_decoder(16#20#)) OR
 					(reg_q452 AND symb_decoder(16#f1#)) OR
 					(reg_q452 AND symb_decoder(16#06#)) OR
 					(reg_q452 AND symb_decoder(16#98#)) OR
 					(reg_q452 AND symb_decoder(16#6c#)) OR
 					(reg_q452 AND symb_decoder(16#8f#)) OR
 					(reg_q452 AND symb_decoder(16#d2#)) OR
 					(reg_q452 AND symb_decoder(16#d8#)) OR
 					(reg_q452 AND symb_decoder(16#f5#)) OR
 					(reg_q452 AND symb_decoder(16#c2#)) OR
 					(reg_q452 AND symb_decoder(16#30#)) OR
 					(reg_q452 AND symb_decoder(16#11#)) OR
 					(reg_q452 AND symb_decoder(16#5d#)) OR
 					(reg_q452 AND symb_decoder(16#18#)) OR
 					(reg_q452 AND symb_decoder(16#12#)) OR
 					(reg_q452 AND symb_decoder(16#64#)) OR
 					(reg_q452 AND symb_decoder(16#91#)) OR
 					(reg_q452 AND symb_decoder(16#ed#)) OR
 					(reg_q452 AND symb_decoder(16#2d#)) OR
 					(reg_q452 AND symb_decoder(16#58#)) OR
 					(reg_q452 AND symb_decoder(16#ff#)) OR
 					(reg_q452 AND symb_decoder(16#c5#)) OR
 					(reg_q452 AND symb_decoder(16#03#)) OR
 					(reg_q452 AND symb_decoder(16#86#)) OR
 					(reg_q452 AND symb_decoder(16#14#)) OR
 					(reg_q452 AND symb_decoder(16#8b#)) OR
 					(reg_q452 AND symb_decoder(16#d0#)) OR
 					(reg_q452 AND symb_decoder(16#eb#)) OR
 					(reg_q452 AND symb_decoder(16#7a#)) OR
 					(reg_q452 AND symb_decoder(16#3a#)) OR
 					(reg_q452 AND symb_decoder(16#b4#)) OR
 					(reg_q452 AND symb_decoder(16#2a#)) OR
 					(reg_q452 AND symb_decoder(16#57#)) OR
 					(reg_q452 AND symb_decoder(16#3f#)) OR
 					(reg_q452 AND symb_decoder(16#60#)) OR
 					(reg_q452 AND symb_decoder(16#f2#)) OR
 					(reg_q452 AND symb_decoder(16#74#)) OR
 					(reg_q452 AND symb_decoder(16#e5#)) OR
 					(reg_q452 AND symb_decoder(16#be#)) OR
 					(reg_q452 AND symb_decoder(16#bc#)) OR
 					(reg_q452 AND symb_decoder(16#92#)) OR
 					(reg_q452 AND symb_decoder(16#e4#)) OR
 					(reg_q452 AND symb_decoder(16#5b#)) OR
 					(reg_q452 AND symb_decoder(16#ba#)) OR
 					(reg_q452 AND symb_decoder(16#7e#)) OR
 					(reg_q452 AND symb_decoder(16#ce#)) OR
 					(reg_q452 AND symb_decoder(16#62#)) OR
 					(reg_q452 AND symb_decoder(16#25#)) OR
 					(reg_q452 AND symb_decoder(16#9f#)) OR
 					(reg_q452 AND symb_decoder(16#da#)) OR
 					(reg_q452 AND symb_decoder(16#32#)) OR
 					(reg_q452 AND symb_decoder(16#c6#)) OR
 					(reg_q452 AND symb_decoder(16#9b#)) OR
 					(reg_q452 AND symb_decoder(16#c3#)) OR
 					(reg_q452 AND symb_decoder(16#65#)) OR
 					(reg_q452 AND symb_decoder(16#37#)) OR
 					(reg_q452 AND symb_decoder(16#c9#)) OR
 					(reg_q452 AND symb_decoder(16#d3#)) OR
 					(reg_q452 AND symb_decoder(16#49#)) OR
 					(reg_q452 AND symb_decoder(16#3e#)) OR
 					(reg_q452 AND symb_decoder(16#c4#)) OR
 					(reg_q452 AND symb_decoder(16#ab#)) OR
 					(reg_q452 AND symb_decoder(16#f7#)) OR
 					(reg_q452 AND symb_decoder(16#e0#)) OR
 					(reg_q452 AND symb_decoder(16#99#)) OR
 					(reg_q452 AND symb_decoder(16#ef#)) OR
 					(reg_q452 AND symb_decoder(16#52#)) OR
 					(reg_q452 AND symb_decoder(16#7c#)) OR
 					(reg_q452 AND symb_decoder(16#b3#)) OR
 					(reg_q452 AND symb_decoder(16#67#)) OR
 					(reg_q452 AND symb_decoder(16#78#)) OR
 					(reg_q452 AND symb_decoder(16#27#)) OR
 					(reg_q452 AND symb_decoder(16#f3#)) OR
 					(reg_q452 AND symb_decoder(16#35#)) OR
 					(reg_q452 AND symb_decoder(16#54#)) OR
 					(reg_q452 AND symb_decoder(16#0c#)) OR
 					(reg_q452 AND symb_decoder(16#1b#)) OR
 					(reg_q452 AND symb_decoder(16#04#)) OR
 					(reg_q452 AND symb_decoder(16#d1#)) OR
 					(reg_q452 AND symb_decoder(16#34#)) OR
 					(reg_q452 AND symb_decoder(16#0d#)) OR
 					(reg_q452 AND symb_decoder(16#85#)) OR
 					(reg_q452 AND symb_decoder(16#8d#)) OR
 					(reg_q452 AND symb_decoder(16#69#)) OR
 					(reg_q452 AND symb_decoder(16#95#)) OR
 					(reg_q452 AND symb_decoder(16#4e#)) OR
 					(reg_q452 AND symb_decoder(16#8c#)) OR
 					(reg_q452 AND symb_decoder(16#fb#)) OR
 					(reg_q452 AND symb_decoder(16#af#)) OR
 					(reg_q452 AND symb_decoder(16#cc#)) OR
 					(reg_q452 AND symb_decoder(16#2e#)) OR
 					(reg_q452 AND symb_decoder(16#d9#)) OR
 					(reg_q452 AND symb_decoder(16#61#)) OR
 					(reg_q452 AND symb_decoder(16#6a#)) OR
 					(reg_q452 AND symb_decoder(16#84#)) OR
 					(reg_q452 AND symb_decoder(16#31#)) OR
 					(reg_q452 AND symb_decoder(16#51#)) OR
 					(reg_q452 AND symb_decoder(16#2b#)) OR
 					(reg_q452 AND symb_decoder(16#82#)) OR
 					(reg_q452 AND symb_decoder(16#02#)) OR
 					(reg_q452 AND symb_decoder(16#d5#)) OR
 					(reg_q452 AND symb_decoder(16#e9#)) OR
 					(reg_q452 AND symb_decoder(16#16#)) OR
 					(reg_q452 AND symb_decoder(16#f0#)) OR
 					(reg_q452 AND symb_decoder(16#dd#)) OR
 					(reg_q452 AND symb_decoder(16#55#)) OR
 					(reg_q452 AND symb_decoder(16#ac#)) OR
 					(reg_q452 AND symb_decoder(16#3c#)) OR
 					(reg_q452 AND symb_decoder(16#53#));
reg_q452_init <= '0' ;
	p_reg_q452: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q452 <= reg_q452_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q452 <= reg_q452_init;
        else
          reg_q452 <= reg_q452_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q556_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q556 AND symb_decoder(16#d9#)) OR
 					(reg_q556 AND symb_decoder(16#f4#)) OR
 					(reg_q556 AND symb_decoder(16#cf#)) OR
 					(reg_q556 AND symb_decoder(16#fd#)) OR
 					(reg_q556 AND symb_decoder(16#b2#)) OR
 					(reg_q556 AND symb_decoder(16#74#)) OR
 					(reg_q556 AND symb_decoder(16#63#)) OR
 					(reg_q556 AND symb_decoder(16#c3#)) OR
 					(reg_q556 AND symb_decoder(16#0f#)) OR
 					(reg_q556 AND symb_decoder(16#e6#)) OR
 					(reg_q556 AND symb_decoder(16#b9#)) OR
 					(reg_q556 AND symb_decoder(16#0b#)) OR
 					(reg_q556 AND symb_decoder(16#3d#)) OR
 					(reg_q556 AND symb_decoder(16#e7#)) OR
 					(reg_q556 AND symb_decoder(16#ba#)) OR
 					(reg_q556 AND symb_decoder(16#8c#)) OR
 					(reg_q556 AND symb_decoder(16#92#)) OR
 					(reg_q556 AND symb_decoder(16#a0#)) OR
 					(reg_q556 AND symb_decoder(16#6e#)) OR
 					(reg_q556 AND symb_decoder(16#fc#)) OR
 					(reg_q556 AND symb_decoder(16#15#)) OR
 					(reg_q556 AND symb_decoder(16#85#)) OR
 					(reg_q556 AND symb_decoder(16#68#)) OR
 					(reg_q556 AND symb_decoder(16#48#)) OR
 					(reg_q556 AND symb_decoder(16#a3#)) OR
 					(reg_q556 AND symb_decoder(16#ea#)) OR
 					(reg_q556 AND symb_decoder(16#8d#)) OR
 					(reg_q556 AND symb_decoder(16#f3#)) OR
 					(reg_q556 AND symb_decoder(16#8f#)) OR
 					(reg_q556 AND symb_decoder(16#6a#)) OR
 					(reg_q556 AND symb_decoder(16#96#)) OR
 					(reg_q556 AND symb_decoder(16#30#)) OR
 					(reg_q556 AND symb_decoder(16#47#)) OR
 					(reg_q556 AND symb_decoder(16#f8#)) OR
 					(reg_q556 AND symb_decoder(16#44#)) OR
 					(reg_q556 AND symb_decoder(16#9f#)) OR
 					(reg_q556 AND symb_decoder(16#de#)) OR
 					(reg_q556 AND symb_decoder(16#0a#)) OR
 					(reg_q556 AND symb_decoder(16#13#)) OR
 					(reg_q556 AND symb_decoder(16#3e#)) OR
 					(reg_q556 AND symb_decoder(16#01#)) OR
 					(reg_q556 AND symb_decoder(16#1a#)) OR
 					(reg_q556 AND symb_decoder(16#7a#)) OR
 					(reg_q556 AND symb_decoder(16#10#)) OR
 					(reg_q556 AND symb_decoder(16#1f#)) OR
 					(reg_q556 AND symb_decoder(16#09#)) OR
 					(reg_q556 AND symb_decoder(16#b5#)) OR
 					(reg_q556 AND symb_decoder(16#65#)) OR
 					(reg_q556 AND symb_decoder(16#db#)) OR
 					(reg_q556 AND symb_decoder(16#d1#)) OR
 					(reg_q556 AND symb_decoder(16#a1#)) OR
 					(reg_q556 AND symb_decoder(16#81#)) OR
 					(reg_q556 AND symb_decoder(16#76#)) OR
 					(reg_q556 AND symb_decoder(16#40#)) OR
 					(reg_q556 AND symb_decoder(16#df#)) OR
 					(reg_q556 AND symb_decoder(16#ab#)) OR
 					(reg_q556 AND symb_decoder(16#5e#)) OR
 					(reg_q556 AND symb_decoder(16#0c#)) OR
 					(reg_q556 AND symb_decoder(16#dd#)) OR
 					(reg_q556 AND symb_decoder(16#95#)) OR
 					(reg_q556 AND symb_decoder(16#fa#)) OR
 					(reg_q556 AND symb_decoder(16#14#)) OR
 					(reg_q556 AND symb_decoder(16#b8#)) OR
 					(reg_q556 AND symb_decoder(16#c6#)) OR
 					(reg_q556 AND symb_decoder(16#70#)) OR
 					(reg_q556 AND symb_decoder(16#e8#)) OR
 					(reg_q556 AND symb_decoder(16#43#)) OR
 					(reg_q556 AND symb_decoder(16#60#)) OR
 					(reg_q556 AND symb_decoder(16#50#)) OR
 					(reg_q556 AND symb_decoder(16#d2#)) OR
 					(reg_q556 AND symb_decoder(16#a8#)) OR
 					(reg_q556 AND symb_decoder(16#54#)) OR
 					(reg_q556 AND symb_decoder(16#55#)) OR
 					(reg_q556 AND symb_decoder(16#49#)) OR
 					(reg_q556 AND symb_decoder(16#d8#)) OR
 					(reg_q556 AND symb_decoder(16#d6#)) OR
 					(reg_q556 AND symb_decoder(16#78#)) OR
 					(reg_q556 AND symb_decoder(16#36#)) OR
 					(reg_q556 AND symb_decoder(16#8a#)) OR
 					(reg_q556 AND symb_decoder(16#2b#)) OR
 					(reg_q556 AND symb_decoder(16#c9#)) OR
 					(reg_q556 AND symb_decoder(16#7c#)) OR
 					(reg_q556 AND symb_decoder(16#ee#)) OR
 					(reg_q556 AND symb_decoder(16#21#)) OR
 					(reg_q556 AND symb_decoder(16#4f#)) OR
 					(reg_q556 AND symb_decoder(16#e0#)) OR
 					(reg_q556 AND symb_decoder(16#80#)) OR
 					(reg_q556 AND symb_decoder(16#3a#)) OR
 					(reg_q556 AND symb_decoder(16#39#)) OR
 					(reg_q556 AND symb_decoder(16#f0#)) OR
 					(reg_q556 AND symb_decoder(16#7f#)) OR
 					(reg_q556 AND symb_decoder(16#7b#)) OR
 					(reg_q556 AND symb_decoder(16#12#)) OR
 					(reg_q556 AND symb_decoder(16#93#)) OR
 					(reg_q556 AND symb_decoder(16#46#)) OR
 					(reg_q556 AND symb_decoder(16#1e#)) OR
 					(reg_q556 AND symb_decoder(16#9e#)) OR
 					(reg_q556 AND symb_decoder(16#90#)) OR
 					(reg_q556 AND symb_decoder(16#fe#)) OR
 					(reg_q556 AND symb_decoder(16#6f#)) OR
 					(reg_q556 AND symb_decoder(16#d4#)) OR
 					(reg_q556 AND symb_decoder(16#71#)) OR
 					(reg_q556 AND symb_decoder(16#a5#)) OR
 					(reg_q556 AND symb_decoder(16#b1#)) OR
 					(reg_q556 AND symb_decoder(16#9c#)) OR
 					(reg_q556 AND symb_decoder(16#4a#)) OR
 					(reg_q556 AND symb_decoder(16#2a#)) OR
 					(reg_q556 AND symb_decoder(16#e5#)) OR
 					(reg_q556 AND symb_decoder(16#5c#)) OR
 					(reg_q556 AND symb_decoder(16#d7#)) OR
 					(reg_q556 AND symb_decoder(16#22#)) OR
 					(reg_q556 AND symb_decoder(16#2e#)) OR
 					(reg_q556 AND symb_decoder(16#cb#)) OR
 					(reg_q556 AND symb_decoder(16#79#)) OR
 					(reg_q556 AND symb_decoder(16#a2#)) OR
 					(reg_q556 AND symb_decoder(16#cc#)) OR
 					(reg_q556 AND symb_decoder(16#2f#)) OR
 					(reg_q556 AND symb_decoder(16#c0#)) OR
 					(reg_q556 AND symb_decoder(16#41#)) OR
 					(reg_q556 AND symb_decoder(16#67#)) OR
 					(reg_q556 AND symb_decoder(16#d3#)) OR
 					(reg_q556 AND symb_decoder(16#e3#)) OR
 					(reg_q556 AND symb_decoder(16#82#)) OR
 					(reg_q556 AND symb_decoder(16#19#)) OR
 					(reg_q556 AND symb_decoder(16#06#)) OR
 					(reg_q556 AND symb_decoder(16#9b#)) OR
 					(reg_q556 AND symb_decoder(16#02#)) OR
 					(reg_q556 AND symb_decoder(16#33#)) OR
 					(reg_q556 AND symb_decoder(16#0d#)) OR
 					(reg_q556 AND symb_decoder(16#42#)) OR
 					(reg_q556 AND symb_decoder(16#3c#)) OR
 					(reg_q556 AND symb_decoder(16#bf#)) OR
 					(reg_q556 AND symb_decoder(16#c8#)) OR
 					(reg_q556 AND symb_decoder(16#aa#)) OR
 					(reg_q556 AND symb_decoder(16#7d#)) OR
 					(reg_q556 AND symb_decoder(16#b6#)) OR
 					(reg_q556 AND symb_decoder(16#05#)) OR
 					(reg_q556 AND symb_decoder(16#1d#)) OR
 					(reg_q556 AND symb_decoder(16#17#)) OR
 					(reg_q556 AND symb_decoder(16#f5#)) OR
 					(reg_q556 AND symb_decoder(16#bd#)) OR
 					(reg_q556 AND symb_decoder(16#a6#)) OR
 					(reg_q556 AND symb_decoder(16#af#)) OR
 					(reg_q556 AND symb_decoder(16#56#)) OR
 					(reg_q556 AND symb_decoder(16#11#)) OR
 					(reg_q556 AND symb_decoder(16#f9#)) OR
 					(reg_q556 AND symb_decoder(16#94#)) OR
 					(reg_q556 AND symb_decoder(16#ff#)) OR
 					(reg_q556 AND symb_decoder(16#ed#)) OR
 					(reg_q556 AND symb_decoder(16#e2#)) OR
 					(reg_q556 AND symb_decoder(16#e1#)) OR
 					(reg_q556 AND symb_decoder(16#9d#)) OR
 					(reg_q556 AND symb_decoder(16#5a#)) OR
 					(reg_q556 AND symb_decoder(16#37#)) OR
 					(reg_q556 AND symb_decoder(16#07#)) OR
 					(reg_q556 AND symb_decoder(16#a7#)) OR
 					(reg_q556 AND symb_decoder(16#8b#)) OR
 					(reg_q556 AND symb_decoder(16#98#)) OR
 					(reg_q556 AND symb_decoder(16#84#)) OR
 					(reg_q556 AND symb_decoder(16#c7#)) OR
 					(reg_q556 AND symb_decoder(16#d0#)) OR
 					(reg_q556 AND symb_decoder(16#73#)) OR
 					(reg_q556 AND symb_decoder(16#c1#)) OR
 					(reg_q556 AND symb_decoder(16#2c#)) OR
 					(reg_q556 AND symb_decoder(16#9a#)) OR
 					(reg_q556 AND symb_decoder(16#b4#)) OR
 					(reg_q556 AND symb_decoder(16#e9#)) OR
 					(reg_q556 AND symb_decoder(16#bc#)) OR
 					(reg_q556 AND symb_decoder(16#f7#)) OR
 					(reg_q556 AND symb_decoder(16#f6#)) OR
 					(reg_q556 AND symb_decoder(16#08#)) OR
 					(reg_q556 AND symb_decoder(16#4d#)) OR
 					(reg_q556 AND symb_decoder(16#26#)) OR
 					(reg_q556 AND symb_decoder(16#58#)) OR
 					(reg_q556 AND symb_decoder(16#64#)) OR
 					(reg_q556 AND symb_decoder(16#62#)) OR
 					(reg_q556 AND symb_decoder(16#91#)) OR
 					(reg_q556 AND symb_decoder(16#32#)) OR
 					(reg_q556 AND symb_decoder(16#29#)) OR
 					(reg_q556 AND symb_decoder(16#6c#)) OR
 					(reg_q556 AND symb_decoder(16#99#)) OR
 					(reg_q556 AND symb_decoder(16#ec#)) OR
 					(reg_q556 AND symb_decoder(16#f2#)) OR
 					(reg_q556 AND symb_decoder(16#c5#)) OR
 					(reg_q556 AND symb_decoder(16#72#)) OR
 					(reg_q556 AND symb_decoder(16#52#)) OR
 					(reg_q556 AND symb_decoder(16#00#)) OR
 					(reg_q556 AND symb_decoder(16#53#)) OR
 					(reg_q556 AND symb_decoder(16#89#)) OR
 					(reg_q556 AND symb_decoder(16#ad#)) OR
 					(reg_q556 AND symb_decoder(16#eb#)) OR
 					(reg_q556 AND symb_decoder(16#0e#)) OR
 					(reg_q556 AND symb_decoder(16#be#)) OR
 					(reg_q556 AND symb_decoder(16#ca#)) OR
 					(reg_q556 AND symb_decoder(16#97#)) OR
 					(reg_q556 AND symb_decoder(16#c2#)) OR
 					(reg_q556 AND symb_decoder(16#a4#)) OR
 					(reg_q556 AND symb_decoder(16#6d#)) OR
 					(reg_q556 AND symb_decoder(16#18#)) OR
 					(reg_q556 AND symb_decoder(16#77#)) OR
 					(reg_q556 AND symb_decoder(16#7e#)) OR
 					(reg_q556 AND symb_decoder(16#b0#)) OR
 					(reg_q556 AND symb_decoder(16#57#)) OR
 					(reg_q556 AND symb_decoder(16#da#)) OR
 					(reg_q556 AND symb_decoder(16#16#)) OR
 					(reg_q556 AND symb_decoder(16#8e#)) OR
 					(reg_q556 AND symb_decoder(16#51#)) OR
 					(reg_q556 AND symb_decoder(16#24#)) OR
 					(reg_q556 AND symb_decoder(16#27#)) OR
 					(reg_q556 AND symb_decoder(16#20#)) OR
 					(reg_q556 AND symb_decoder(16#5b#)) OR
 					(reg_q556 AND symb_decoder(16#87#)) OR
 					(reg_q556 AND symb_decoder(16#31#)) OR
 					(reg_q556 AND symb_decoder(16#03#)) OR
 					(reg_q556 AND symb_decoder(16#75#)) OR
 					(reg_q556 AND symb_decoder(16#fb#)) OR
 					(reg_q556 AND symb_decoder(16#4e#)) OR
 					(reg_q556 AND symb_decoder(16#bb#)) OR
 					(reg_q556 AND symb_decoder(16#c4#)) OR
 					(reg_q556 AND symb_decoder(16#d5#)) OR
 					(reg_q556 AND symb_decoder(16#ef#)) OR
 					(reg_q556 AND symb_decoder(16#5d#)) OR
 					(reg_q556 AND symb_decoder(16#ae#)) OR
 					(reg_q556 AND symb_decoder(16#3f#)) OR
 					(reg_q556 AND symb_decoder(16#4b#)) OR
 					(reg_q556 AND symb_decoder(16#3b#)) OR
 					(reg_q556 AND symb_decoder(16#f1#)) OR
 					(reg_q556 AND symb_decoder(16#b3#)) OR
 					(reg_q556 AND symb_decoder(16#28#)) OR
 					(reg_q556 AND symb_decoder(16#86#)) OR
 					(reg_q556 AND symb_decoder(16#38#)) OR
 					(reg_q556 AND symb_decoder(16#59#)) OR
 					(reg_q556 AND symb_decoder(16#25#)) OR
 					(reg_q556 AND symb_decoder(16#6b#)) OR
 					(reg_q556 AND symb_decoder(16#b7#)) OR
 					(reg_q556 AND symb_decoder(16#2d#)) OR
 					(reg_q556 AND symb_decoder(16#66#)) OR
 					(reg_q556 AND symb_decoder(16#35#)) OR
 					(reg_q556 AND symb_decoder(16#34#)) OR
 					(reg_q556 AND symb_decoder(16#e4#)) OR
 					(reg_q556 AND symb_decoder(16#dc#)) OR
 					(reg_q556 AND symb_decoder(16#1c#)) OR
 					(reg_q556 AND symb_decoder(16#45#)) OR
 					(reg_q556 AND symb_decoder(16#88#)) OR
 					(reg_q556 AND symb_decoder(16#04#)) OR
 					(reg_q556 AND symb_decoder(16#23#)) OR
 					(reg_q556 AND symb_decoder(16#ac#)) OR
 					(reg_q556 AND symb_decoder(16#ce#)) OR
 					(reg_q556 AND symb_decoder(16#83#)) OR
 					(reg_q556 AND symb_decoder(16#61#)) OR
 					(reg_q556 AND symb_decoder(16#1b#)) OR
 					(reg_q556 AND symb_decoder(16#4c#)) OR
 					(reg_q556 AND symb_decoder(16#5f#)) OR
 					(reg_q556 AND symb_decoder(16#69#)) OR
 					(reg_q556 AND symb_decoder(16#cd#)) OR
 					(reg_q556 AND symb_decoder(16#a9#));
reg_q556_init <= '0' ;
	p_reg_q556: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q556 <= reg_q556_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q556 <= reg_q556_init;
        else
          reg_q556 <= reg_q556_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1111_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1111 AND symb_decoder(16#ba#)) OR
 					(reg_q1111 AND symb_decoder(16#9b#)) OR
 					(reg_q1111 AND symb_decoder(16#35#)) OR
 					(reg_q1111 AND symb_decoder(16#e3#)) OR
 					(reg_q1111 AND symb_decoder(16#77#)) OR
 					(reg_q1111 AND symb_decoder(16#34#)) OR
 					(reg_q1111 AND symb_decoder(16#d6#)) OR
 					(reg_q1111 AND symb_decoder(16#1f#)) OR
 					(reg_q1111 AND symb_decoder(16#c7#)) OR
 					(reg_q1111 AND symb_decoder(16#b6#)) OR
 					(reg_q1111 AND symb_decoder(16#29#)) OR
 					(reg_q1111 AND symb_decoder(16#f3#)) OR
 					(reg_q1111 AND symb_decoder(16#dc#)) OR
 					(reg_q1111 AND symb_decoder(16#66#)) OR
 					(reg_q1111 AND symb_decoder(16#21#)) OR
 					(reg_q1111 AND symb_decoder(16#00#)) OR
 					(reg_q1111 AND symb_decoder(16#b0#)) OR
 					(reg_q1111 AND symb_decoder(16#f2#)) OR
 					(reg_q1111 AND symb_decoder(16#38#)) OR
 					(reg_q1111 AND symb_decoder(16#78#)) OR
 					(reg_q1111 AND symb_decoder(16#27#)) OR
 					(reg_q1111 AND symb_decoder(16#08#)) OR
 					(reg_q1111 AND symb_decoder(16#bf#)) OR
 					(reg_q1111 AND symb_decoder(16#f4#)) OR
 					(reg_q1111 AND symb_decoder(16#16#)) OR
 					(reg_q1111 AND symb_decoder(16#cc#)) OR
 					(reg_q1111 AND symb_decoder(16#70#)) OR
 					(reg_q1111 AND symb_decoder(16#ff#)) OR
 					(reg_q1111 AND symb_decoder(16#32#)) OR
 					(reg_q1111 AND symb_decoder(16#4c#)) OR
 					(reg_q1111 AND symb_decoder(16#15#)) OR
 					(reg_q1111 AND symb_decoder(16#3b#)) OR
 					(reg_q1111 AND symb_decoder(16#63#)) OR
 					(reg_q1111 AND symb_decoder(16#0a#)) OR
 					(reg_q1111 AND symb_decoder(16#d2#)) OR
 					(reg_q1111 AND symb_decoder(16#8b#)) OR
 					(reg_q1111 AND symb_decoder(16#c6#)) OR
 					(reg_q1111 AND symb_decoder(16#a6#)) OR
 					(reg_q1111 AND symb_decoder(16#86#)) OR
 					(reg_q1111 AND symb_decoder(16#5a#)) OR
 					(reg_q1111 AND symb_decoder(16#72#)) OR
 					(reg_q1111 AND symb_decoder(16#1d#)) OR
 					(reg_q1111 AND symb_decoder(16#57#)) OR
 					(reg_q1111 AND symb_decoder(16#98#)) OR
 					(reg_q1111 AND symb_decoder(16#8d#)) OR
 					(reg_q1111 AND symb_decoder(16#19#)) OR
 					(reg_q1111 AND symb_decoder(16#12#)) OR
 					(reg_q1111 AND symb_decoder(16#53#)) OR
 					(reg_q1111 AND symb_decoder(16#51#)) OR
 					(reg_q1111 AND symb_decoder(16#b8#)) OR
 					(reg_q1111 AND symb_decoder(16#20#)) OR
 					(reg_q1111 AND symb_decoder(16#9e#)) OR
 					(reg_q1111 AND symb_decoder(16#5c#)) OR
 					(reg_q1111 AND symb_decoder(16#ef#)) OR
 					(reg_q1111 AND symb_decoder(16#17#)) OR
 					(reg_q1111 AND symb_decoder(16#9f#)) OR
 					(reg_q1111 AND symb_decoder(16#88#)) OR
 					(reg_q1111 AND symb_decoder(16#92#)) OR
 					(reg_q1111 AND symb_decoder(16#8f#)) OR
 					(reg_q1111 AND symb_decoder(16#62#)) OR
 					(reg_q1111 AND symb_decoder(16#40#)) OR
 					(reg_q1111 AND symb_decoder(16#a3#)) OR
 					(reg_q1111 AND symb_decoder(16#97#)) OR
 					(reg_q1111 AND symb_decoder(16#0d#)) OR
 					(reg_q1111 AND symb_decoder(16#c4#)) OR
 					(reg_q1111 AND symb_decoder(16#06#)) OR
 					(reg_q1111 AND symb_decoder(16#49#)) OR
 					(reg_q1111 AND symb_decoder(16#13#)) OR
 					(reg_q1111 AND symb_decoder(16#6c#)) OR
 					(reg_q1111 AND symb_decoder(16#9c#)) OR
 					(reg_q1111 AND symb_decoder(16#4e#)) OR
 					(reg_q1111 AND symb_decoder(16#67#)) OR
 					(reg_q1111 AND symb_decoder(16#3f#)) OR
 					(reg_q1111 AND symb_decoder(16#25#)) OR
 					(reg_q1111 AND symb_decoder(16#ea#)) OR
 					(reg_q1111 AND symb_decoder(16#3a#)) OR
 					(reg_q1111 AND symb_decoder(16#ad#)) OR
 					(reg_q1111 AND symb_decoder(16#e1#)) OR
 					(reg_q1111 AND symb_decoder(16#a0#)) OR
 					(reg_q1111 AND symb_decoder(16#e4#)) OR
 					(reg_q1111 AND symb_decoder(16#a9#)) OR
 					(reg_q1111 AND symb_decoder(16#d7#)) OR
 					(reg_q1111 AND symb_decoder(16#a7#)) OR
 					(reg_q1111 AND symb_decoder(16#68#)) OR
 					(reg_q1111 AND symb_decoder(16#da#)) OR
 					(reg_q1111 AND symb_decoder(16#6d#)) OR
 					(reg_q1111 AND symb_decoder(16#80#)) OR
 					(reg_q1111 AND symb_decoder(16#d0#)) OR
 					(reg_q1111 AND symb_decoder(16#23#)) OR
 					(reg_q1111 AND symb_decoder(16#75#)) OR
 					(reg_q1111 AND symb_decoder(16#87#)) OR
 					(reg_q1111 AND symb_decoder(16#37#)) OR
 					(reg_q1111 AND symb_decoder(16#dd#)) OR
 					(reg_q1111 AND symb_decoder(16#81#)) OR
 					(reg_q1111 AND symb_decoder(16#d5#)) OR
 					(reg_q1111 AND symb_decoder(16#fc#)) OR
 					(reg_q1111 AND symb_decoder(16#f7#)) OR
 					(reg_q1111 AND symb_decoder(16#1c#)) OR
 					(reg_q1111 AND symb_decoder(16#aa#)) OR
 					(reg_q1111 AND symb_decoder(16#fa#)) OR
 					(reg_q1111 AND symb_decoder(16#c8#)) OR
 					(reg_q1111 AND symb_decoder(16#30#)) OR
 					(reg_q1111 AND symb_decoder(16#48#)) OR
 					(reg_q1111 AND symb_decoder(16#39#)) OR
 					(reg_q1111 AND symb_decoder(16#bc#)) OR
 					(reg_q1111 AND symb_decoder(16#de#)) OR
 					(reg_q1111 AND symb_decoder(16#f5#)) OR
 					(reg_q1111 AND symb_decoder(16#43#)) OR
 					(reg_q1111 AND symb_decoder(16#b4#)) OR
 					(reg_q1111 AND symb_decoder(16#61#)) OR
 					(reg_q1111 AND symb_decoder(16#7e#)) OR
 					(reg_q1111 AND symb_decoder(16#3c#)) OR
 					(reg_q1111 AND symb_decoder(16#a8#)) OR
 					(reg_q1111 AND symb_decoder(16#3d#)) OR
 					(reg_q1111 AND symb_decoder(16#2b#)) OR
 					(reg_q1111 AND symb_decoder(16#01#)) OR
 					(reg_q1111 AND symb_decoder(16#d8#)) OR
 					(reg_q1111 AND symb_decoder(16#a1#)) OR
 					(reg_q1111 AND symb_decoder(16#c3#)) OR
 					(reg_q1111 AND symb_decoder(16#ed#)) OR
 					(reg_q1111 AND symb_decoder(16#99#)) OR
 					(reg_q1111 AND symb_decoder(16#46#)) OR
 					(reg_q1111 AND symb_decoder(16#26#)) OR
 					(reg_q1111 AND symb_decoder(16#83#)) OR
 					(reg_q1111 AND symb_decoder(16#7b#)) OR
 					(reg_q1111 AND symb_decoder(16#6b#)) OR
 					(reg_q1111 AND symb_decoder(16#be#)) OR
 					(reg_q1111 AND symb_decoder(16#96#)) OR
 					(reg_q1111 AND symb_decoder(16#71#)) OR
 					(reg_q1111 AND symb_decoder(16#2e#)) OR
 					(reg_q1111 AND symb_decoder(16#d9#)) OR
 					(reg_q1111 AND symb_decoder(16#6f#)) OR
 					(reg_q1111 AND symb_decoder(16#fb#)) OR
 					(reg_q1111 AND symb_decoder(16#c9#)) OR
 					(reg_q1111 AND symb_decoder(16#22#)) OR
 					(reg_q1111 AND symb_decoder(16#5e#)) OR
 					(reg_q1111 AND symb_decoder(16#2d#)) OR
 					(reg_q1111 AND symb_decoder(16#4b#)) OR
 					(reg_q1111 AND symb_decoder(16#52#)) OR
 					(reg_q1111 AND symb_decoder(16#8e#)) OR
 					(reg_q1111 AND symb_decoder(16#04#)) OR
 					(reg_q1111 AND symb_decoder(16#cb#)) OR
 					(reg_q1111 AND symb_decoder(16#11#)) OR
 					(reg_q1111 AND symb_decoder(16#ec#)) OR
 					(reg_q1111 AND symb_decoder(16#02#)) OR
 					(reg_q1111 AND symb_decoder(16#ae#)) OR
 					(reg_q1111 AND symb_decoder(16#65#)) OR
 					(reg_q1111 AND symb_decoder(16#45#)) OR
 					(reg_q1111 AND symb_decoder(16#db#)) OR
 					(reg_q1111 AND symb_decoder(16#ab#)) OR
 					(reg_q1111 AND symb_decoder(16#fe#)) OR
 					(reg_q1111 AND symb_decoder(16#f9#)) OR
 					(reg_q1111 AND symb_decoder(16#df#)) OR
 					(reg_q1111 AND symb_decoder(16#6e#)) OR
 					(reg_q1111 AND symb_decoder(16#82#)) OR
 					(reg_q1111 AND symb_decoder(16#6a#)) OR
 					(reg_q1111 AND symb_decoder(16#33#)) OR
 					(reg_q1111 AND symb_decoder(16#c1#)) OR
 					(reg_q1111 AND symb_decoder(16#18#)) OR
 					(reg_q1111 AND symb_decoder(16#7c#)) OR
 					(reg_q1111 AND symb_decoder(16#ac#)) OR
 					(reg_q1111 AND symb_decoder(16#0b#)) OR
 					(reg_q1111 AND symb_decoder(16#24#)) OR
 					(reg_q1111 AND symb_decoder(16#1b#)) OR
 					(reg_q1111 AND symb_decoder(16#05#)) OR
 					(reg_q1111 AND symb_decoder(16#e9#)) OR
 					(reg_q1111 AND symb_decoder(16#e5#)) OR
 					(reg_q1111 AND symb_decoder(16#e6#)) OR
 					(reg_q1111 AND symb_decoder(16#10#)) OR
 					(reg_q1111 AND symb_decoder(16#bb#)) OR
 					(reg_q1111 AND symb_decoder(16#c0#)) OR
 					(reg_q1111 AND symb_decoder(16#47#)) OR
 					(reg_q1111 AND symb_decoder(16#1e#)) OR
 					(reg_q1111 AND symb_decoder(16#74#)) OR
 					(reg_q1111 AND symb_decoder(16#5b#)) OR
 					(reg_q1111 AND symb_decoder(16#03#)) OR
 					(reg_q1111 AND symb_decoder(16#59#)) OR
 					(reg_q1111 AND symb_decoder(16#07#)) OR
 					(reg_q1111 AND symb_decoder(16#5d#)) OR
 					(reg_q1111 AND symb_decoder(16#2a#)) OR
 					(reg_q1111 AND symb_decoder(16#cd#)) OR
 					(reg_q1111 AND symb_decoder(16#41#)) OR
 					(reg_q1111 AND symb_decoder(16#a4#)) OR
 					(reg_q1111 AND symb_decoder(16#89#)) OR
 					(reg_q1111 AND symb_decoder(16#d4#)) OR
 					(reg_q1111 AND symb_decoder(16#7a#)) OR
 					(reg_q1111 AND symb_decoder(16#3e#)) OR
 					(reg_q1111 AND symb_decoder(16#fd#)) OR
 					(reg_q1111 AND symb_decoder(16#56#)) OR
 					(reg_q1111 AND symb_decoder(16#31#)) OR
 					(reg_q1111 AND symb_decoder(16#d3#)) OR
 					(reg_q1111 AND symb_decoder(16#b1#)) OR
 					(reg_q1111 AND symb_decoder(16#2c#)) OR
 					(reg_q1111 AND symb_decoder(16#8c#)) OR
 					(reg_q1111 AND symb_decoder(16#76#)) OR
 					(reg_q1111 AND symb_decoder(16#58#)) OR
 					(reg_q1111 AND symb_decoder(16#79#)) OR
 					(reg_q1111 AND symb_decoder(16#5f#)) OR
 					(reg_q1111 AND symb_decoder(16#0f#)) OR
 					(reg_q1111 AND symb_decoder(16#8a#)) OR
 					(reg_q1111 AND symb_decoder(16#4d#)) OR
 					(reg_q1111 AND symb_decoder(16#73#)) OR
 					(reg_q1111 AND symb_decoder(16#54#)) OR
 					(reg_q1111 AND symb_decoder(16#ca#)) OR
 					(reg_q1111 AND symb_decoder(16#b2#)) OR
 					(reg_q1111 AND symb_decoder(16#90#)) OR
 					(reg_q1111 AND symb_decoder(16#cf#)) OR
 					(reg_q1111 AND symb_decoder(16#0c#)) OR
 					(reg_q1111 AND symb_decoder(16#f0#)) OR
 					(reg_q1111 AND symb_decoder(16#69#)) OR
 					(reg_q1111 AND symb_decoder(16#e8#)) OR
 					(reg_q1111 AND symb_decoder(16#c5#)) OR
 					(reg_q1111 AND symb_decoder(16#e7#)) OR
 					(reg_q1111 AND symb_decoder(16#2f#)) OR
 					(reg_q1111 AND symb_decoder(16#e2#)) OR
 					(reg_q1111 AND symb_decoder(16#84#)) OR
 					(reg_q1111 AND symb_decoder(16#af#)) OR
 					(reg_q1111 AND symb_decoder(16#42#)) OR
 					(reg_q1111 AND symb_decoder(16#f1#)) OR
 					(reg_q1111 AND symb_decoder(16#4a#)) OR
 					(reg_q1111 AND symb_decoder(16#1a#)) OR
 					(reg_q1111 AND symb_decoder(16#a2#)) OR
 					(reg_q1111 AND symb_decoder(16#0e#)) OR
 					(reg_q1111 AND symb_decoder(16#9d#)) OR
 					(reg_q1111 AND symb_decoder(16#14#)) OR
 					(reg_q1111 AND symb_decoder(16#b9#)) OR
 					(reg_q1111 AND symb_decoder(16#e0#)) OR
 					(reg_q1111 AND symb_decoder(16#f6#)) OR
 					(reg_q1111 AND symb_decoder(16#ee#)) OR
 					(reg_q1111 AND symb_decoder(16#9a#)) OR
 					(reg_q1111 AND symb_decoder(16#7f#)) OR
 					(reg_q1111 AND symb_decoder(16#28#)) OR
 					(reg_q1111 AND symb_decoder(16#d1#)) OR
 					(reg_q1111 AND symb_decoder(16#95#)) OR
 					(reg_q1111 AND symb_decoder(16#55#)) OR
 					(reg_q1111 AND symb_decoder(16#36#)) OR
 					(reg_q1111 AND symb_decoder(16#b7#)) OR
 					(reg_q1111 AND symb_decoder(16#60#)) OR
 					(reg_q1111 AND symb_decoder(16#c2#)) OR
 					(reg_q1111 AND symb_decoder(16#85#)) OR
 					(reg_q1111 AND symb_decoder(16#b5#)) OR
 					(reg_q1111 AND symb_decoder(16#4f#)) OR
 					(reg_q1111 AND symb_decoder(16#93#)) OR
 					(reg_q1111 AND symb_decoder(16#a5#)) OR
 					(reg_q1111 AND symb_decoder(16#50#)) OR
 					(reg_q1111 AND symb_decoder(16#09#)) OR
 					(reg_q1111 AND symb_decoder(16#f8#)) OR
 					(reg_q1111 AND symb_decoder(16#7d#)) OR
 					(reg_q1111 AND symb_decoder(16#ce#)) OR
 					(reg_q1111 AND symb_decoder(16#64#)) OR
 					(reg_q1111 AND symb_decoder(16#91#)) OR
 					(reg_q1111 AND symb_decoder(16#eb#)) OR
 					(reg_q1111 AND symb_decoder(16#bd#)) OR
 					(reg_q1111 AND symb_decoder(16#94#)) OR
 					(reg_q1111 AND symb_decoder(16#b3#)) OR
 					(reg_q1111 AND symb_decoder(16#44#));
reg_q1111_init <= '0' ;
	p_reg_q1111: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1111 <= reg_q1111_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1111 <= reg_q1111_init;
        else
          reg_q1111 <= reg_q1111_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1644_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1644 AND symb_decoder(16#d0#)) OR
 					(reg_q1644 AND symb_decoder(16#69#)) OR
 					(reg_q1644 AND symb_decoder(16#b4#)) OR
 					(reg_q1644 AND symb_decoder(16#1a#)) OR
 					(reg_q1644 AND symb_decoder(16#76#)) OR
 					(reg_q1644 AND symb_decoder(16#c3#)) OR
 					(reg_q1644 AND symb_decoder(16#b7#)) OR
 					(reg_q1644 AND symb_decoder(16#36#)) OR
 					(reg_q1644 AND symb_decoder(16#03#)) OR
 					(reg_q1644 AND symb_decoder(16#b3#)) OR
 					(reg_q1644 AND symb_decoder(16#15#)) OR
 					(reg_q1644 AND symb_decoder(16#59#)) OR
 					(reg_q1644 AND symb_decoder(16#c7#)) OR
 					(reg_q1644 AND symb_decoder(16#00#)) OR
 					(reg_q1644 AND symb_decoder(16#70#)) OR
 					(reg_q1644 AND symb_decoder(16#ca#)) OR
 					(reg_q1644 AND symb_decoder(16#47#)) OR
 					(reg_q1644 AND symb_decoder(16#1e#)) OR
 					(reg_q1644 AND symb_decoder(16#f6#)) OR
 					(reg_q1644 AND symb_decoder(16#3f#)) OR
 					(reg_q1644 AND symb_decoder(16#4e#)) OR
 					(reg_q1644 AND symb_decoder(16#aa#)) OR
 					(reg_q1644 AND symb_decoder(16#8b#)) OR
 					(reg_q1644 AND symb_decoder(16#37#)) OR
 					(reg_q1644 AND symb_decoder(16#17#)) OR
 					(reg_q1644 AND symb_decoder(16#d9#)) OR
 					(reg_q1644 AND symb_decoder(16#9c#)) OR
 					(reg_q1644 AND symb_decoder(16#a4#)) OR
 					(reg_q1644 AND symb_decoder(16#89#)) OR
 					(reg_q1644 AND symb_decoder(16#61#)) OR
 					(reg_q1644 AND symb_decoder(16#cf#)) OR
 					(reg_q1644 AND symb_decoder(16#19#)) OR
 					(reg_q1644 AND symb_decoder(16#ea#)) OR
 					(reg_q1644 AND symb_decoder(16#07#)) OR
 					(reg_q1644 AND symb_decoder(16#b5#)) OR
 					(reg_q1644 AND symb_decoder(16#02#)) OR
 					(reg_q1644 AND symb_decoder(16#e4#)) OR
 					(reg_q1644 AND symb_decoder(16#66#)) OR
 					(reg_q1644 AND symb_decoder(16#79#)) OR
 					(reg_q1644 AND symb_decoder(16#b2#)) OR
 					(reg_q1644 AND symb_decoder(16#84#)) OR
 					(reg_q1644 AND symb_decoder(16#25#)) OR
 					(reg_q1644 AND symb_decoder(16#0d#)) OR
 					(reg_q1644 AND symb_decoder(16#08#)) OR
 					(reg_q1644 AND symb_decoder(16#35#)) OR
 					(reg_q1644 AND symb_decoder(16#60#)) OR
 					(reg_q1644 AND symb_decoder(16#fd#)) OR
 					(reg_q1644 AND symb_decoder(16#bc#)) OR
 					(reg_q1644 AND symb_decoder(16#98#)) OR
 					(reg_q1644 AND symb_decoder(16#94#)) OR
 					(reg_q1644 AND symb_decoder(16#5f#)) OR
 					(reg_q1644 AND symb_decoder(16#32#)) OR
 					(reg_q1644 AND symb_decoder(16#da#)) OR
 					(reg_q1644 AND symb_decoder(16#2a#)) OR
 					(reg_q1644 AND symb_decoder(16#3a#)) OR
 					(reg_q1644 AND symb_decoder(16#cc#)) OR
 					(reg_q1644 AND symb_decoder(16#88#)) OR
 					(reg_q1644 AND symb_decoder(16#82#)) OR
 					(reg_q1644 AND symb_decoder(16#20#)) OR
 					(reg_q1644 AND symb_decoder(16#c2#)) OR
 					(reg_q1644 AND symb_decoder(16#ee#)) OR
 					(reg_q1644 AND symb_decoder(16#57#)) OR
 					(reg_q1644 AND symb_decoder(16#ad#)) OR
 					(reg_q1644 AND symb_decoder(16#73#)) OR
 					(reg_q1644 AND symb_decoder(16#a0#)) OR
 					(reg_q1644 AND symb_decoder(16#fe#)) OR
 					(reg_q1644 AND symb_decoder(16#95#)) OR
 					(reg_q1644 AND symb_decoder(16#d1#)) OR
 					(reg_q1644 AND symb_decoder(16#7a#)) OR
 					(reg_q1644 AND symb_decoder(16#4a#)) OR
 					(reg_q1644 AND symb_decoder(16#8d#)) OR
 					(reg_q1644 AND symb_decoder(16#64#)) OR
 					(reg_q1644 AND symb_decoder(16#31#)) OR
 					(reg_q1644 AND symb_decoder(16#51#)) OR
 					(reg_q1644 AND symb_decoder(16#ab#)) OR
 					(reg_q1644 AND symb_decoder(16#04#)) OR
 					(reg_q1644 AND symb_decoder(16#81#)) OR
 					(reg_q1644 AND symb_decoder(16#f7#)) OR
 					(reg_q1644 AND symb_decoder(16#46#)) OR
 					(reg_q1644 AND symb_decoder(16#3e#)) OR
 					(reg_q1644 AND symb_decoder(16#0b#)) OR
 					(reg_q1644 AND symb_decoder(16#7e#)) OR
 					(reg_q1644 AND symb_decoder(16#09#)) OR
 					(reg_q1644 AND symb_decoder(16#75#)) OR
 					(reg_q1644 AND symb_decoder(16#41#)) OR
 					(reg_q1644 AND symb_decoder(16#86#)) OR
 					(reg_q1644 AND symb_decoder(16#e1#)) OR
 					(reg_q1644 AND symb_decoder(16#dd#)) OR
 					(reg_q1644 AND symb_decoder(16#c8#)) OR
 					(reg_q1644 AND symb_decoder(16#e2#)) OR
 					(reg_q1644 AND symb_decoder(16#c0#)) OR
 					(reg_q1644 AND symb_decoder(16#65#)) OR
 					(reg_q1644 AND symb_decoder(16#4d#)) OR
 					(reg_q1644 AND symb_decoder(16#fa#)) OR
 					(reg_q1644 AND symb_decoder(16#ec#)) OR
 					(reg_q1644 AND symb_decoder(16#85#)) OR
 					(reg_q1644 AND symb_decoder(16#a8#)) OR
 					(reg_q1644 AND symb_decoder(16#56#)) OR
 					(reg_q1644 AND symb_decoder(16#40#)) OR
 					(reg_q1644 AND symb_decoder(16#de#)) OR
 					(reg_q1644 AND symb_decoder(16#50#)) OR
 					(reg_q1644 AND symb_decoder(16#c9#)) OR
 					(reg_q1644 AND symb_decoder(16#ff#)) OR
 					(reg_q1644 AND symb_decoder(16#01#)) OR
 					(reg_q1644 AND symb_decoder(16#cd#)) OR
 					(reg_q1644 AND symb_decoder(16#ef#)) OR
 					(reg_q1644 AND symb_decoder(16#b1#)) OR
 					(reg_q1644 AND symb_decoder(16#12#)) OR
 					(reg_q1644 AND symb_decoder(16#8e#)) OR
 					(reg_q1644 AND symb_decoder(16#a1#)) OR
 					(reg_q1644 AND symb_decoder(16#ac#)) OR
 					(reg_q1644 AND symb_decoder(16#cb#)) OR
 					(reg_q1644 AND symb_decoder(16#96#)) OR
 					(reg_q1644 AND symb_decoder(16#af#)) OR
 					(reg_q1644 AND symb_decoder(16#6a#)) OR
 					(reg_q1644 AND symb_decoder(16#54#)) OR
 					(reg_q1644 AND symb_decoder(16#8a#)) OR
 					(reg_q1644 AND symb_decoder(16#d4#)) OR
 					(reg_q1644 AND symb_decoder(16#a3#)) OR
 					(reg_q1644 AND symb_decoder(16#43#)) OR
 					(reg_q1644 AND symb_decoder(16#11#)) OR
 					(reg_q1644 AND symb_decoder(16#3c#)) OR
 					(reg_q1644 AND symb_decoder(16#f1#)) OR
 					(reg_q1644 AND symb_decoder(16#58#)) OR
 					(reg_q1644 AND symb_decoder(16#e3#)) OR
 					(reg_q1644 AND symb_decoder(16#eb#)) OR
 					(reg_q1644 AND symb_decoder(16#c5#)) OR
 					(reg_q1644 AND symb_decoder(16#77#)) OR
 					(reg_q1644 AND symb_decoder(16#48#)) OR
 					(reg_q1644 AND symb_decoder(16#0f#)) OR
 					(reg_q1644 AND symb_decoder(16#16#)) OR
 					(reg_q1644 AND symb_decoder(16#24#)) OR
 					(reg_q1644 AND symb_decoder(16#f3#)) OR
 					(reg_q1644 AND symb_decoder(16#22#)) OR
 					(reg_q1644 AND symb_decoder(16#33#)) OR
 					(reg_q1644 AND symb_decoder(16#3b#)) OR
 					(reg_q1644 AND symb_decoder(16#7d#)) OR
 					(reg_q1644 AND symb_decoder(16#c1#)) OR
 					(reg_q1644 AND symb_decoder(16#13#)) OR
 					(reg_q1644 AND symb_decoder(16#10#)) OR
 					(reg_q1644 AND symb_decoder(16#dc#)) OR
 					(reg_q1644 AND symb_decoder(16#4c#)) OR
 					(reg_q1644 AND symb_decoder(16#fb#)) OR
 					(reg_q1644 AND symb_decoder(16#df#)) OR
 					(reg_q1644 AND symb_decoder(16#7c#)) OR
 					(reg_q1644 AND symb_decoder(16#2e#)) OR
 					(reg_q1644 AND symb_decoder(16#2d#)) OR
 					(reg_q1644 AND symb_decoder(16#a2#)) OR
 					(reg_q1644 AND symb_decoder(16#78#)) OR
 					(reg_q1644 AND symb_decoder(16#e5#)) OR
 					(reg_q1644 AND symb_decoder(16#d6#)) OR
 					(reg_q1644 AND symb_decoder(16#6f#)) OR
 					(reg_q1644 AND symb_decoder(16#d3#)) OR
 					(reg_q1644 AND symb_decoder(16#42#)) OR
 					(reg_q1644 AND symb_decoder(16#8f#)) OR
 					(reg_q1644 AND symb_decoder(16#9e#)) OR
 					(reg_q1644 AND symb_decoder(16#ae#)) OR
 					(reg_q1644 AND symb_decoder(16#23#)) OR
 					(reg_q1644 AND symb_decoder(16#27#)) OR
 					(reg_q1644 AND symb_decoder(16#f5#)) OR
 					(reg_q1644 AND symb_decoder(16#1b#)) OR
 					(reg_q1644 AND symb_decoder(16#f8#)) OR
 					(reg_q1644 AND symb_decoder(16#90#)) OR
 					(reg_q1644 AND symb_decoder(16#ba#)) OR
 					(reg_q1644 AND symb_decoder(16#9f#)) OR
 					(reg_q1644 AND symb_decoder(16#f2#)) OR
 					(reg_q1644 AND symb_decoder(16#e9#)) OR
 					(reg_q1644 AND symb_decoder(16#a5#)) OR
 					(reg_q1644 AND symb_decoder(16#b0#)) OR
 					(reg_q1644 AND symb_decoder(16#0e#)) OR
 					(reg_q1644 AND symb_decoder(16#52#)) OR
 					(reg_q1644 AND symb_decoder(16#fc#)) OR
 					(reg_q1644 AND symb_decoder(16#05#)) OR
 					(reg_q1644 AND symb_decoder(16#e6#)) OR
 					(reg_q1644 AND symb_decoder(16#9b#)) OR
 					(reg_q1644 AND symb_decoder(16#80#)) OR
 					(reg_q1644 AND symb_decoder(16#87#)) OR
 					(reg_q1644 AND symb_decoder(16#c6#)) OR
 					(reg_q1644 AND symb_decoder(16#83#)) OR
 					(reg_q1644 AND symb_decoder(16#8c#)) OR
 					(reg_q1644 AND symb_decoder(16#4b#)) OR
 					(reg_q1644 AND symb_decoder(16#bf#)) OR
 					(reg_q1644 AND symb_decoder(16#a9#)) OR
 					(reg_q1644 AND symb_decoder(16#1d#)) OR
 					(reg_q1644 AND symb_decoder(16#a7#)) OR
 					(reg_q1644 AND symb_decoder(16#18#)) OR
 					(reg_q1644 AND symb_decoder(16#92#)) OR
 					(reg_q1644 AND symb_decoder(16#9a#)) OR
 					(reg_q1644 AND symb_decoder(16#f4#)) OR
 					(reg_q1644 AND symb_decoder(16#5c#)) OR
 					(reg_q1644 AND symb_decoder(16#d8#)) OR
 					(reg_q1644 AND symb_decoder(16#5b#)) OR
 					(reg_q1644 AND symb_decoder(16#2b#)) OR
 					(reg_q1644 AND symb_decoder(16#6c#)) OR
 					(reg_q1644 AND symb_decoder(16#f0#)) OR
 					(reg_q1644 AND symb_decoder(16#39#)) OR
 					(reg_q1644 AND symb_decoder(16#44#)) OR
 					(reg_q1644 AND symb_decoder(16#b6#)) OR
 					(reg_q1644 AND symb_decoder(16#6e#)) OR
 					(reg_q1644 AND symb_decoder(16#6d#)) OR
 					(reg_q1644 AND symb_decoder(16#55#)) OR
 					(reg_q1644 AND symb_decoder(16#1c#)) OR
 					(reg_q1644 AND symb_decoder(16#0a#)) OR
 					(reg_q1644 AND symb_decoder(16#be#)) OR
 					(reg_q1644 AND symb_decoder(16#38#)) OR
 					(reg_q1644 AND symb_decoder(16#2c#)) OR
 					(reg_q1644 AND symb_decoder(16#e8#)) OR
 					(reg_q1644 AND symb_decoder(16#34#)) OR
 					(reg_q1644 AND symb_decoder(16#45#)) OR
 					(reg_q1644 AND symb_decoder(16#91#)) OR
 					(reg_q1644 AND symb_decoder(16#d5#)) OR
 					(reg_q1644 AND symb_decoder(16#2f#)) OR
 					(reg_q1644 AND symb_decoder(16#28#)) OR
 					(reg_q1644 AND symb_decoder(16#97#)) OR
 					(reg_q1644 AND symb_decoder(16#26#)) OR
 					(reg_q1644 AND symb_decoder(16#63#)) OR
 					(reg_q1644 AND symb_decoder(16#c4#)) OR
 					(reg_q1644 AND symb_decoder(16#9d#)) OR
 					(reg_q1644 AND symb_decoder(16#0c#)) OR
 					(reg_q1644 AND symb_decoder(16#e0#)) OR
 					(reg_q1644 AND symb_decoder(16#71#)) OR
 					(reg_q1644 AND symb_decoder(16#3d#)) OR
 					(reg_q1644 AND symb_decoder(16#30#)) OR
 					(reg_q1644 AND symb_decoder(16#bd#)) OR
 					(reg_q1644 AND symb_decoder(16#93#)) OR
 					(reg_q1644 AND symb_decoder(16#68#)) OR
 					(reg_q1644 AND symb_decoder(16#21#)) OR
 					(reg_q1644 AND symb_decoder(16#99#)) OR
 					(reg_q1644 AND symb_decoder(16#5e#)) OR
 					(reg_q1644 AND symb_decoder(16#ce#)) OR
 					(reg_q1644 AND symb_decoder(16#e7#)) OR
 					(reg_q1644 AND symb_decoder(16#d7#)) OR
 					(reg_q1644 AND symb_decoder(16#d2#)) OR
 					(reg_q1644 AND symb_decoder(16#53#)) OR
 					(reg_q1644 AND symb_decoder(16#74#)) OR
 					(reg_q1644 AND symb_decoder(16#b8#)) OR
 					(reg_q1644 AND symb_decoder(16#62#)) OR
 					(reg_q1644 AND symb_decoder(16#67#)) OR
 					(reg_q1644 AND symb_decoder(16#72#)) OR
 					(reg_q1644 AND symb_decoder(16#29#)) OR
 					(reg_q1644 AND symb_decoder(16#f9#)) OR
 					(reg_q1644 AND symb_decoder(16#14#)) OR
 					(reg_q1644 AND symb_decoder(16#1f#)) OR
 					(reg_q1644 AND symb_decoder(16#b9#)) OR
 					(reg_q1644 AND symb_decoder(16#ed#)) OR
 					(reg_q1644 AND symb_decoder(16#49#)) OR
 					(reg_q1644 AND symb_decoder(16#7f#)) OR
 					(reg_q1644 AND symb_decoder(16#7b#)) OR
 					(reg_q1644 AND symb_decoder(16#6b#)) OR
 					(reg_q1644 AND symb_decoder(16#06#)) OR
 					(reg_q1644 AND symb_decoder(16#db#)) OR
 					(reg_q1644 AND symb_decoder(16#bb#)) OR
 					(reg_q1644 AND symb_decoder(16#a6#)) OR
 					(reg_q1644 AND symb_decoder(16#4f#)) OR
 					(reg_q1644 AND symb_decoder(16#5d#)) OR
 					(reg_q1644 AND symb_decoder(16#5a#));
reg_q1644_init <= '0' ;
	p_reg_q1644: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1644 <= reg_q1644_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1644 <= reg_q1644_init;
        else
          reg_q1644 <= reg_q1644_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2249_in <= (reg_q2249 AND symb_decoder(16#34#)) OR
 					(reg_q2249 AND symb_decoder(16#32#)) OR
 					(reg_q2249 AND symb_decoder(16#33#)) OR
 					(reg_q2249 AND symb_decoder(16#35#)) OR
 					(reg_q2249 AND symb_decoder(16#37#)) OR
 					(reg_q2249 AND symb_decoder(16#31#)) OR
 					(reg_q2249 AND symb_decoder(16#36#)) OR
 					(reg_q2249 AND symb_decoder(16#30#)) OR
 					(reg_q2249 AND symb_decoder(16#38#)) OR
 					(reg_q2249 AND symb_decoder(16#39#)) OR
 					(reg_q2247 AND symb_decoder(16#33#)) OR
 					(reg_q2247 AND symb_decoder(16#38#)) OR
 					(reg_q2247 AND symb_decoder(16#32#)) OR
 					(reg_q2247 AND symb_decoder(16#37#)) OR
 					(reg_q2247 AND symb_decoder(16#31#)) OR
 					(reg_q2247 AND symb_decoder(16#34#)) OR
 					(reg_q2247 AND symb_decoder(16#36#)) OR
 					(reg_q2247 AND symb_decoder(16#35#)) OR
 					(reg_q2247 AND symb_decoder(16#39#)) OR
 					(reg_q2247 AND symb_decoder(16#30#));
reg_q2249_init <= '0' ;
	p_reg_q2249: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2249 <= reg_q2249_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2249 <= reg_q2249_init;
        else
          reg_q2249 <= reg_q2249_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q799_in <= (reg_q797 AND symb_decoder(16#2e#));
reg_q799_init <= '0' ;
	p_reg_q799: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q799 <= reg_q799_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q799 <= reg_q799_init;
        else
          reg_q799 <= reg_q799_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q801_in <= (reg_q799 AND symb_decoder(16#38#)) OR
 					(reg_q799 AND symb_decoder(16#34#)) OR
 					(reg_q799 AND symb_decoder(16#33#)) OR
 					(reg_q799 AND symb_decoder(16#36#)) OR
 					(reg_q799 AND symb_decoder(16#30#)) OR
 					(reg_q799 AND symb_decoder(16#31#)) OR
 					(reg_q799 AND symb_decoder(16#35#)) OR
 					(reg_q799 AND symb_decoder(16#39#)) OR
 					(reg_q799 AND symb_decoder(16#32#)) OR
 					(reg_q799 AND symb_decoder(16#37#)) OR
 					(reg_q801 AND symb_decoder(16#37#)) OR
 					(reg_q801 AND symb_decoder(16#34#)) OR
 					(reg_q801 AND symb_decoder(16#38#)) OR
 					(reg_q801 AND symb_decoder(16#33#)) OR
 					(reg_q801 AND symb_decoder(16#35#)) OR
 					(reg_q801 AND symb_decoder(16#31#)) OR
 					(reg_q801 AND symb_decoder(16#39#)) OR
 					(reg_q801 AND symb_decoder(16#30#)) OR
 					(reg_q801 AND symb_decoder(16#36#)) OR
 					(reg_q801 AND symb_decoder(16#32#));
reg_q801_init <= '0' ;
	p_reg_q801: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q801 <= reg_q801_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q801 <= reg_q801_init;
        else
          reg_q801 <= reg_q801_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1195_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1195 AND symb_decoder(16#f0#)) OR
 					(reg_q1195 AND symb_decoder(16#4a#)) OR
 					(reg_q1195 AND symb_decoder(16#15#)) OR
 					(reg_q1195 AND symb_decoder(16#4f#)) OR
 					(reg_q1195 AND symb_decoder(16#a2#)) OR
 					(reg_q1195 AND symb_decoder(16#d2#)) OR
 					(reg_q1195 AND symb_decoder(16#77#)) OR
 					(reg_q1195 AND symb_decoder(16#68#)) OR
 					(reg_q1195 AND symb_decoder(16#55#)) OR
 					(reg_q1195 AND symb_decoder(16#96#)) OR
 					(reg_q1195 AND symb_decoder(16#fc#)) OR
 					(reg_q1195 AND symb_decoder(16#b3#)) OR
 					(reg_q1195 AND symb_decoder(16#35#)) OR
 					(reg_q1195 AND symb_decoder(16#ce#)) OR
 					(reg_q1195 AND symb_decoder(16#c5#)) OR
 					(reg_q1195 AND symb_decoder(16#6a#)) OR
 					(reg_q1195 AND symb_decoder(16#66#)) OR
 					(reg_q1195 AND symb_decoder(16#c4#)) OR
 					(reg_q1195 AND symb_decoder(16#aa#)) OR
 					(reg_q1195 AND symb_decoder(16#70#)) OR
 					(reg_q1195 AND symb_decoder(16#b6#)) OR
 					(reg_q1195 AND symb_decoder(16#8d#)) OR
 					(reg_q1195 AND symb_decoder(16#23#)) OR
 					(reg_q1195 AND symb_decoder(16#64#)) OR
 					(reg_q1195 AND symb_decoder(16#cf#)) OR
 					(reg_q1195 AND symb_decoder(16#f4#)) OR
 					(reg_q1195 AND symb_decoder(16#52#)) OR
 					(reg_q1195 AND symb_decoder(16#d3#)) OR
 					(reg_q1195 AND symb_decoder(16#df#)) OR
 					(reg_q1195 AND symb_decoder(16#ac#)) OR
 					(reg_q1195 AND symb_decoder(16#5a#)) OR
 					(reg_q1195 AND symb_decoder(16#0b#)) OR
 					(reg_q1195 AND symb_decoder(16#40#)) OR
 					(reg_q1195 AND symb_decoder(16#12#)) OR
 					(reg_q1195 AND symb_decoder(16#1d#)) OR
 					(reg_q1195 AND symb_decoder(16#b5#)) OR
 					(reg_q1195 AND symb_decoder(16#11#)) OR
 					(reg_q1195 AND symb_decoder(16#d0#)) OR
 					(reg_q1195 AND symb_decoder(16#34#)) OR
 					(reg_q1195 AND symb_decoder(16#7c#)) OR
 					(reg_q1195 AND symb_decoder(16#e5#)) OR
 					(reg_q1195 AND symb_decoder(16#ee#)) OR
 					(reg_q1195 AND symb_decoder(16#e9#)) OR
 					(reg_q1195 AND symb_decoder(16#bb#)) OR
 					(reg_q1195 AND symb_decoder(16#a1#)) OR
 					(reg_q1195 AND symb_decoder(16#16#)) OR
 					(reg_q1195 AND symb_decoder(16#7e#)) OR
 					(reg_q1195 AND symb_decoder(16#0c#)) OR
 					(reg_q1195 AND symb_decoder(16#d4#)) OR
 					(reg_q1195 AND symb_decoder(16#3c#)) OR
 					(reg_q1195 AND symb_decoder(16#79#)) OR
 					(reg_q1195 AND symb_decoder(16#53#)) OR
 					(reg_q1195 AND symb_decoder(16#e3#)) OR
 					(reg_q1195 AND symb_decoder(16#14#)) OR
 					(reg_q1195 AND symb_decoder(16#d5#)) OR
 					(reg_q1195 AND symb_decoder(16#07#)) OR
 					(reg_q1195 AND symb_decoder(16#39#)) OR
 					(reg_q1195 AND symb_decoder(16#95#)) OR
 					(reg_q1195 AND symb_decoder(16#3e#)) OR
 					(reg_q1195 AND symb_decoder(16#29#)) OR
 					(reg_q1195 AND symb_decoder(16#b1#)) OR
 					(reg_q1195 AND symb_decoder(16#46#)) OR
 					(reg_q1195 AND symb_decoder(16#38#)) OR
 					(reg_q1195 AND symb_decoder(16#2b#)) OR
 					(reg_q1195 AND symb_decoder(16#1e#)) OR
 					(reg_q1195 AND symb_decoder(16#9b#)) OR
 					(reg_q1195 AND symb_decoder(16#89#)) OR
 					(reg_q1195 AND symb_decoder(16#ad#)) OR
 					(reg_q1195 AND symb_decoder(16#09#)) OR
 					(reg_q1195 AND symb_decoder(16#fd#)) OR
 					(reg_q1195 AND symb_decoder(16#bc#)) OR
 					(reg_q1195 AND symb_decoder(16#62#)) OR
 					(reg_q1195 AND symb_decoder(16#67#)) OR
 					(reg_q1195 AND symb_decoder(16#92#)) OR
 					(reg_q1195 AND symb_decoder(16#bd#)) OR
 					(reg_q1195 AND symb_decoder(16#b7#)) OR
 					(reg_q1195 AND symb_decoder(16#bf#)) OR
 					(reg_q1195 AND symb_decoder(16#fa#)) OR
 					(reg_q1195 AND symb_decoder(16#fe#)) OR
 					(reg_q1195 AND symb_decoder(16#c1#)) OR
 					(reg_q1195 AND symb_decoder(16#78#)) OR
 					(reg_q1195 AND symb_decoder(16#59#)) OR
 					(reg_q1195 AND symb_decoder(16#3f#)) OR
 					(reg_q1195 AND symb_decoder(16#1b#)) OR
 					(reg_q1195 AND symb_decoder(16#60#)) OR
 					(reg_q1195 AND symb_decoder(16#cb#)) OR
 					(reg_q1195 AND symb_decoder(16#db#)) OR
 					(reg_q1195 AND symb_decoder(16#f3#)) OR
 					(reg_q1195 AND symb_decoder(16#33#)) OR
 					(reg_q1195 AND symb_decoder(16#8e#)) OR
 					(reg_q1195 AND symb_decoder(16#a4#)) OR
 					(reg_q1195 AND symb_decoder(16#a5#)) OR
 					(reg_q1195 AND symb_decoder(16#17#)) OR
 					(reg_q1195 AND symb_decoder(16#6f#)) OR
 					(reg_q1195 AND symb_decoder(16#d6#)) OR
 					(reg_q1195 AND symb_decoder(16#9f#)) OR
 					(reg_q1195 AND symb_decoder(16#00#)) OR
 					(reg_q1195 AND symb_decoder(16#25#)) OR
 					(reg_q1195 AND symb_decoder(16#f7#)) OR
 					(reg_q1195 AND symb_decoder(16#28#)) OR
 					(reg_q1195 AND symb_decoder(16#98#)) OR
 					(reg_q1195 AND symb_decoder(16#93#)) OR
 					(reg_q1195 AND symb_decoder(16#13#)) OR
 					(reg_q1195 AND symb_decoder(16#26#)) OR
 					(reg_q1195 AND symb_decoder(16#47#)) OR
 					(reg_q1195 AND symb_decoder(16#da#)) OR
 					(reg_q1195 AND symb_decoder(16#a6#)) OR
 					(reg_q1195 AND symb_decoder(16#e0#)) OR
 					(reg_q1195 AND symb_decoder(16#82#)) OR
 					(reg_q1195 AND symb_decoder(16#65#)) OR
 					(reg_q1195 AND symb_decoder(16#a0#)) OR
 					(reg_q1195 AND symb_decoder(16#a7#)) OR
 					(reg_q1195 AND symb_decoder(16#e7#)) OR
 					(reg_q1195 AND symb_decoder(16#d7#)) OR
 					(reg_q1195 AND symb_decoder(16#f6#)) OR
 					(reg_q1195 AND symb_decoder(16#80#)) OR
 					(reg_q1195 AND symb_decoder(16#21#)) OR
 					(reg_q1195 AND symb_decoder(16#7b#)) OR
 					(reg_q1195 AND symb_decoder(16#03#)) OR
 					(reg_q1195 AND symb_decoder(16#0a#)) OR
 					(reg_q1195 AND symb_decoder(16#9a#)) OR
 					(reg_q1195 AND symb_decoder(16#b9#)) OR
 					(reg_q1195 AND symb_decoder(16#c6#)) OR
 					(reg_q1195 AND symb_decoder(16#de#)) OR
 					(reg_q1195 AND symb_decoder(16#7d#)) OR
 					(reg_q1195 AND symb_decoder(16#06#)) OR
 					(reg_q1195 AND symb_decoder(16#45#)) OR
 					(reg_q1195 AND symb_decoder(16#f8#)) OR
 					(reg_q1195 AND symb_decoder(16#b2#)) OR
 					(reg_q1195 AND symb_decoder(16#eb#)) OR
 					(reg_q1195 AND symb_decoder(16#c9#)) OR
 					(reg_q1195 AND symb_decoder(16#2a#)) OR
 					(reg_q1195 AND symb_decoder(16#2d#)) OR
 					(reg_q1195 AND symb_decoder(16#5c#)) OR
 					(reg_q1195 AND symb_decoder(16#f5#)) OR
 					(reg_q1195 AND symb_decoder(16#8f#)) OR
 					(reg_q1195 AND symb_decoder(16#f1#)) OR
 					(reg_q1195 AND symb_decoder(16#49#)) OR
 					(reg_q1195 AND symb_decoder(16#f9#)) OR
 					(reg_q1195 AND symb_decoder(16#18#)) OR
 					(reg_q1195 AND symb_decoder(16#6c#)) OR
 					(reg_q1195 AND symb_decoder(16#42#)) OR
 					(reg_q1195 AND symb_decoder(16#ba#)) OR
 					(reg_q1195 AND symb_decoder(16#97#)) OR
 					(reg_q1195 AND symb_decoder(16#86#)) OR
 					(reg_q1195 AND symb_decoder(16#c8#)) OR
 					(reg_q1195 AND symb_decoder(16#ea#)) OR
 					(reg_q1195 AND symb_decoder(16#1a#)) OR
 					(reg_q1195 AND symb_decoder(16#01#)) OR
 					(reg_q1195 AND symb_decoder(16#5b#)) OR
 					(reg_q1195 AND symb_decoder(16#71#)) OR
 					(reg_q1195 AND symb_decoder(16#61#)) OR
 					(reg_q1195 AND symb_decoder(16#43#)) OR
 					(reg_q1195 AND symb_decoder(16#ec#)) OR
 					(reg_q1195 AND symb_decoder(16#4d#)) OR
 					(reg_q1195 AND symb_decoder(16#94#)) OR
 					(reg_q1195 AND symb_decoder(16#72#)) OR
 					(reg_q1195 AND symb_decoder(16#6e#)) OR
 					(reg_q1195 AND symb_decoder(16#41#)) OR
 					(reg_q1195 AND symb_decoder(16#d8#)) OR
 					(reg_q1195 AND symb_decoder(16#1f#)) OR
 					(reg_q1195 AND symb_decoder(16#4c#)) OR
 					(reg_q1195 AND symb_decoder(16#ef#)) OR
 					(reg_q1195 AND symb_decoder(16#af#)) OR
 					(reg_q1195 AND symb_decoder(16#48#)) OR
 					(reg_q1195 AND symb_decoder(16#c2#)) OR
 					(reg_q1195 AND symb_decoder(16#24#)) OR
 					(reg_q1195 AND symb_decoder(16#51#)) OR
 					(reg_q1195 AND symb_decoder(16#3a#)) OR
 					(reg_q1195 AND symb_decoder(16#90#)) OR
 					(reg_q1195 AND symb_decoder(16#e8#)) OR
 					(reg_q1195 AND symb_decoder(16#4e#)) OR
 					(reg_q1195 AND symb_decoder(16#b4#)) OR
 					(reg_q1195 AND symb_decoder(16#cd#)) OR
 					(reg_q1195 AND symb_decoder(16#a8#)) OR
 					(reg_q1195 AND symb_decoder(16#0f#)) OR
 					(reg_q1195 AND symb_decoder(16#e1#)) OR
 					(reg_q1195 AND symb_decoder(16#ca#)) OR
 					(reg_q1195 AND symb_decoder(16#30#)) OR
 					(reg_q1195 AND symb_decoder(16#36#)) OR
 					(reg_q1195 AND symb_decoder(16#99#)) OR
 					(reg_q1195 AND symb_decoder(16#9e#)) OR
 					(reg_q1195 AND symb_decoder(16#19#)) OR
 					(reg_q1195 AND symb_decoder(16#05#)) OR
 					(reg_q1195 AND symb_decoder(16#08#)) OR
 					(reg_q1195 AND symb_decoder(16#a3#)) OR
 					(reg_q1195 AND symb_decoder(16#dc#)) OR
 					(reg_q1195 AND symb_decoder(16#50#)) OR
 					(reg_q1195 AND symb_decoder(16#91#)) OR
 					(reg_q1195 AND symb_decoder(16#69#)) OR
 					(reg_q1195 AND symb_decoder(16#87#)) OR
 					(reg_q1195 AND symb_decoder(16#20#)) OR
 					(reg_q1195 AND symb_decoder(16#2f#)) OR
 					(reg_q1195 AND symb_decoder(16#84#)) OR
 					(reg_q1195 AND symb_decoder(16#0d#)) OR
 					(reg_q1195 AND symb_decoder(16#44#)) OR
 					(reg_q1195 AND symb_decoder(16#c3#)) OR
 					(reg_q1195 AND symb_decoder(16#22#)) OR
 					(reg_q1195 AND symb_decoder(16#76#)) OR
 					(reg_q1195 AND symb_decoder(16#9c#)) OR
 					(reg_q1195 AND symb_decoder(16#5f#)) OR
 					(reg_q1195 AND symb_decoder(16#7a#)) OR
 					(reg_q1195 AND symb_decoder(16#04#)) OR
 					(reg_q1195 AND symb_decoder(16#e4#)) OR
 					(reg_q1195 AND symb_decoder(16#e2#)) OR
 					(reg_q1195 AND symb_decoder(16#cc#)) OR
 					(reg_q1195 AND symb_decoder(16#5e#)) OR
 					(reg_q1195 AND symb_decoder(16#63#)) OR
 					(reg_q1195 AND symb_decoder(16#75#)) OR
 					(reg_q1195 AND symb_decoder(16#8b#)) OR
 					(reg_q1195 AND symb_decoder(16#ff#)) OR
 					(reg_q1195 AND symb_decoder(16#3d#)) OR
 					(reg_q1195 AND symb_decoder(16#ab#)) OR
 					(reg_q1195 AND symb_decoder(16#d1#)) OR
 					(reg_q1195 AND symb_decoder(16#85#)) OR
 					(reg_q1195 AND symb_decoder(16#dd#)) OR
 					(reg_q1195 AND symb_decoder(16#6b#)) OR
 					(reg_q1195 AND symb_decoder(16#10#)) OR
 					(reg_q1195 AND symb_decoder(16#8c#)) OR
 					(reg_q1195 AND symb_decoder(16#4b#)) OR
 					(reg_q1195 AND symb_decoder(16#58#)) OR
 					(reg_q1195 AND symb_decoder(16#b0#)) OR
 					(reg_q1195 AND symb_decoder(16#9d#)) OR
 					(reg_q1195 AND symb_decoder(16#6d#)) OR
 					(reg_q1195 AND symb_decoder(16#b8#)) OR
 					(reg_q1195 AND symb_decoder(16#73#)) OR
 					(reg_q1195 AND symb_decoder(16#ae#)) OR
 					(reg_q1195 AND symb_decoder(16#31#)) OR
 					(reg_q1195 AND symb_decoder(16#8a#)) OR
 					(reg_q1195 AND symb_decoder(16#57#)) OR
 					(reg_q1195 AND symb_decoder(16#3b#)) OR
 					(reg_q1195 AND symb_decoder(16#32#)) OR
 					(reg_q1195 AND symb_decoder(16#2e#)) OR
 					(reg_q1195 AND symb_decoder(16#1c#)) OR
 					(reg_q1195 AND symb_decoder(16#c0#)) OR
 					(reg_q1195 AND symb_decoder(16#c7#)) OR
 					(reg_q1195 AND symb_decoder(16#74#)) OR
 					(reg_q1195 AND symb_decoder(16#88#)) OR
 					(reg_q1195 AND symb_decoder(16#54#)) OR
 					(reg_q1195 AND symb_decoder(16#ed#)) OR
 					(reg_q1195 AND symb_decoder(16#f2#)) OR
 					(reg_q1195 AND symb_decoder(16#7f#)) OR
 					(reg_q1195 AND symb_decoder(16#0e#)) OR
 					(reg_q1195 AND symb_decoder(16#37#)) OR
 					(reg_q1195 AND symb_decoder(16#a9#)) OR
 					(reg_q1195 AND symb_decoder(16#e6#)) OR
 					(reg_q1195 AND symb_decoder(16#be#)) OR
 					(reg_q1195 AND symb_decoder(16#d9#)) OR
 					(reg_q1195 AND symb_decoder(16#2c#)) OR
 					(reg_q1195 AND symb_decoder(16#27#)) OR
 					(reg_q1195 AND symb_decoder(16#02#)) OR
 					(reg_q1195 AND symb_decoder(16#5d#)) OR
 					(reg_q1195 AND symb_decoder(16#81#)) OR
 					(reg_q1195 AND symb_decoder(16#83#)) OR
 					(reg_q1195 AND symb_decoder(16#fb#)) OR
 					(reg_q1195 AND symb_decoder(16#56#));
reg_q1195_init <= '0' ;
	p_reg_q1195: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1195 <= reg_q1195_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1195 <= reg_q1195_init;
        else
          reg_q1195 <= reg_q1195_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2373_in <= (reg_q2373 AND symb_decoder(16#37#)) OR
 					(reg_q2373 AND symb_decoder(16#35#)) OR
 					(reg_q2373 AND symb_decoder(16#39#)) OR
 					(reg_q2373 AND symb_decoder(16#38#)) OR
 					(reg_q2373 AND symb_decoder(16#34#)) OR
 					(reg_q2373 AND symb_decoder(16#30#)) OR
 					(reg_q2373 AND symb_decoder(16#33#)) OR
 					(reg_q2373 AND symb_decoder(16#36#)) OR
 					(reg_q2373 AND symb_decoder(16#31#)) OR
 					(reg_q2373 AND symb_decoder(16#32#)) OR
 					(reg_q2371 AND symb_decoder(16#32#)) OR
 					(reg_q2371 AND symb_decoder(16#35#)) OR
 					(reg_q2371 AND symb_decoder(16#33#)) OR
 					(reg_q2371 AND symb_decoder(16#39#)) OR
 					(reg_q2371 AND symb_decoder(16#31#)) OR
 					(reg_q2371 AND symb_decoder(16#36#)) OR
 					(reg_q2371 AND symb_decoder(16#34#)) OR
 					(reg_q2371 AND symb_decoder(16#30#)) OR
 					(reg_q2371 AND symb_decoder(16#38#)) OR
 					(reg_q2371 AND symb_decoder(16#37#));
reg_q2373_init <= '0' ;
	p_reg_q2373: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2373 <= reg_q2373_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2373 <= reg_q2373_init;
        else
          reg_q2373 <= reg_q2373_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q91_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q91 AND symb_decoder(16#6e#)) OR
 					(reg_q91 AND symb_decoder(16#07#)) OR
 					(reg_q91 AND symb_decoder(16#f9#)) OR
 					(reg_q91 AND symb_decoder(16#a5#)) OR
 					(reg_q91 AND symb_decoder(16#01#)) OR
 					(reg_q91 AND symb_decoder(16#79#)) OR
 					(reg_q91 AND symb_decoder(16#cf#)) OR
 					(reg_q91 AND symb_decoder(16#5c#)) OR
 					(reg_q91 AND symb_decoder(16#c2#)) OR
 					(reg_q91 AND symb_decoder(16#b1#)) OR
 					(reg_q91 AND symb_decoder(16#4e#)) OR
 					(reg_q91 AND symb_decoder(16#51#)) OR
 					(reg_q91 AND symb_decoder(16#fc#)) OR
 					(reg_q91 AND symb_decoder(16#e9#)) OR
 					(reg_q91 AND symb_decoder(16#71#)) OR
 					(reg_q91 AND symb_decoder(16#e7#)) OR
 					(reg_q91 AND symb_decoder(16#1f#)) OR
 					(reg_q91 AND symb_decoder(16#48#)) OR
 					(reg_q91 AND symb_decoder(16#f0#)) OR
 					(reg_q91 AND symb_decoder(16#9b#)) OR
 					(reg_q91 AND symb_decoder(16#0c#)) OR
 					(reg_q91 AND symb_decoder(16#62#)) OR
 					(reg_q91 AND symb_decoder(16#aa#)) OR
 					(reg_q91 AND symb_decoder(16#bb#)) OR
 					(reg_q91 AND symb_decoder(16#ff#)) OR
 					(reg_q91 AND symb_decoder(16#2e#)) OR
 					(reg_q91 AND symb_decoder(16#ec#)) OR
 					(reg_q91 AND symb_decoder(16#f3#)) OR
 					(reg_q91 AND symb_decoder(16#eb#)) OR
 					(reg_q91 AND symb_decoder(16#d6#)) OR
 					(reg_q91 AND symb_decoder(16#6b#)) OR
 					(reg_q91 AND symb_decoder(16#ae#)) OR
 					(reg_q91 AND symb_decoder(16#1b#)) OR
 					(reg_q91 AND symb_decoder(16#93#)) OR
 					(reg_q91 AND symb_decoder(16#53#)) OR
 					(reg_q91 AND symb_decoder(16#50#)) OR
 					(reg_q91 AND symb_decoder(16#0a#)) OR
 					(reg_q91 AND symb_decoder(16#77#)) OR
 					(reg_q91 AND symb_decoder(16#99#)) OR
 					(reg_q91 AND symb_decoder(16#69#)) OR
 					(reg_q91 AND symb_decoder(16#54#)) OR
 					(reg_q91 AND symb_decoder(16#f6#)) OR
 					(reg_q91 AND symb_decoder(16#6c#)) OR
 					(reg_q91 AND symb_decoder(16#b6#)) OR
 					(reg_q91 AND symb_decoder(16#e5#)) OR
 					(reg_q91 AND symb_decoder(16#a3#)) OR
 					(reg_q91 AND symb_decoder(16#9e#)) OR
 					(reg_q91 AND symb_decoder(16#2d#)) OR
 					(reg_q91 AND symb_decoder(16#38#)) OR
 					(reg_q91 AND symb_decoder(16#9c#)) OR
 					(reg_q91 AND symb_decoder(16#94#)) OR
 					(reg_q91 AND symb_decoder(16#b0#)) OR
 					(reg_q91 AND symb_decoder(16#df#)) OR
 					(reg_q91 AND symb_decoder(16#57#)) OR
 					(reg_q91 AND symb_decoder(16#3b#)) OR
 					(reg_q91 AND symb_decoder(16#a7#)) OR
 					(reg_q91 AND symb_decoder(16#55#)) OR
 					(reg_q91 AND symb_decoder(16#b4#)) OR
 					(reg_q91 AND symb_decoder(16#1c#)) OR
 					(reg_q91 AND symb_decoder(16#68#)) OR
 					(reg_q91 AND symb_decoder(16#e3#)) OR
 					(reg_q91 AND symb_decoder(16#8b#)) OR
 					(reg_q91 AND symb_decoder(16#c3#)) OR
 					(reg_q91 AND symb_decoder(16#1a#)) OR
 					(reg_q91 AND symb_decoder(16#36#)) OR
 					(reg_q91 AND symb_decoder(16#4b#)) OR
 					(reg_q91 AND symb_decoder(16#23#)) OR
 					(reg_q91 AND symb_decoder(16#76#)) OR
 					(reg_q91 AND symb_decoder(16#c9#)) OR
 					(reg_q91 AND symb_decoder(16#81#)) OR
 					(reg_q91 AND symb_decoder(16#83#)) OR
 					(reg_q91 AND symb_decoder(16#c6#)) OR
 					(reg_q91 AND symb_decoder(16#86#)) OR
 					(reg_q91 AND symb_decoder(16#a1#)) OR
 					(reg_q91 AND symb_decoder(16#d2#)) OR
 					(reg_q91 AND symb_decoder(16#8c#)) OR
 					(reg_q91 AND symb_decoder(16#49#)) OR
 					(reg_q91 AND symb_decoder(16#e1#)) OR
 					(reg_q91 AND symb_decoder(16#ef#)) OR
 					(reg_q91 AND symb_decoder(16#87#)) OR
 					(reg_q91 AND symb_decoder(16#98#)) OR
 					(reg_q91 AND symb_decoder(16#0d#)) OR
 					(reg_q91 AND symb_decoder(16#be#)) OR
 					(reg_q91 AND symb_decoder(16#f1#)) OR
 					(reg_q91 AND symb_decoder(16#fa#)) OR
 					(reg_q91 AND symb_decoder(16#42#)) OR
 					(reg_q91 AND symb_decoder(16#46#)) OR
 					(reg_q91 AND symb_decoder(16#dc#)) OR
 					(reg_q91 AND symb_decoder(16#ab#)) OR
 					(reg_q91 AND symb_decoder(16#96#)) OR
 					(reg_q91 AND symb_decoder(16#52#)) OR
 					(reg_q91 AND symb_decoder(16#15#)) OR
 					(reg_q91 AND symb_decoder(16#63#)) OR
 					(reg_q91 AND symb_decoder(16#e2#)) OR
 					(reg_q91 AND symb_decoder(16#91#)) OR
 					(reg_q91 AND symb_decoder(16#f5#)) OR
 					(reg_q91 AND symb_decoder(16#e0#)) OR
 					(reg_q91 AND symb_decoder(16#24#)) OR
 					(reg_q91 AND symb_decoder(16#37#)) OR
 					(reg_q91 AND symb_decoder(16#92#)) OR
 					(reg_q91 AND symb_decoder(16#bf#)) OR
 					(reg_q91 AND symb_decoder(16#8f#)) OR
 					(reg_q91 AND symb_decoder(16#7a#)) OR
 					(reg_q91 AND symb_decoder(16#a0#)) OR
 					(reg_q91 AND symb_decoder(16#a8#)) OR
 					(reg_q91 AND symb_decoder(16#75#)) OR
 					(reg_q91 AND symb_decoder(16#64#)) OR
 					(reg_q91 AND symb_decoder(16#7b#)) OR
 					(reg_q91 AND symb_decoder(16#f4#)) OR
 					(reg_q91 AND symb_decoder(16#ca#)) OR
 					(reg_q91 AND symb_decoder(16#73#)) OR
 					(reg_q91 AND symb_decoder(16#89#)) OR
 					(reg_q91 AND symb_decoder(16#ea#)) OR
 					(reg_q91 AND symb_decoder(16#a2#)) OR
 					(reg_q91 AND symb_decoder(16#58#)) OR
 					(reg_q91 AND symb_decoder(16#b3#)) OR
 					(reg_q91 AND symb_decoder(16#5e#)) OR
 					(reg_q91 AND symb_decoder(16#40#)) OR
 					(reg_q91 AND symb_decoder(16#d8#)) OR
 					(reg_q91 AND symb_decoder(16#da#)) OR
 					(reg_q91 AND symb_decoder(16#3a#)) OR
 					(reg_q91 AND symb_decoder(16#ba#)) OR
 					(reg_q91 AND symb_decoder(16#ad#)) OR
 					(reg_q91 AND symb_decoder(16#19#)) OR
 					(reg_q91 AND symb_decoder(16#67#)) OR
 					(reg_q91 AND symb_decoder(16#00#)) OR
 					(reg_q91 AND symb_decoder(16#6f#)) OR
 					(reg_q91 AND symb_decoder(16#d1#)) OR
 					(reg_q91 AND symb_decoder(16#5b#)) OR
 					(reg_q91 AND symb_decoder(16#59#)) OR
 					(reg_q91 AND symb_decoder(16#35#)) OR
 					(reg_q91 AND symb_decoder(16#82#)) OR
 					(reg_q91 AND symb_decoder(16#2b#)) OR
 					(reg_q91 AND symb_decoder(16#ed#)) OR
 					(reg_q91 AND symb_decoder(16#22#)) OR
 					(reg_q91 AND symb_decoder(16#02#)) OR
 					(reg_q91 AND symb_decoder(16#a9#)) OR
 					(reg_q91 AND symb_decoder(16#11#)) OR
 					(reg_q91 AND symb_decoder(16#13#)) OR
 					(reg_q91 AND symb_decoder(16#ee#)) OR
 					(reg_q91 AND symb_decoder(16#e6#)) OR
 					(reg_q91 AND symb_decoder(16#d4#)) OR
 					(reg_q91 AND symb_decoder(16#33#)) OR
 					(reg_q91 AND symb_decoder(16#c7#)) OR
 					(reg_q91 AND symb_decoder(16#d0#)) OR
 					(reg_q91 AND symb_decoder(16#78#)) OR
 					(reg_q91 AND symb_decoder(16#2c#)) OR
 					(reg_q91 AND symb_decoder(16#03#)) OR
 					(reg_q91 AND symb_decoder(16#ce#)) OR
 					(reg_q91 AND symb_decoder(16#18#)) OR
 					(reg_q91 AND symb_decoder(16#29#)) OR
 					(reg_q91 AND symb_decoder(16#5d#)) OR
 					(reg_q91 AND symb_decoder(16#14#)) OR
 					(reg_q91 AND symb_decoder(16#2f#)) OR
 					(reg_q91 AND symb_decoder(16#28#)) OR
 					(reg_q91 AND symb_decoder(16#c4#)) OR
 					(reg_q91 AND symb_decoder(16#4a#)) OR
 					(reg_q91 AND symb_decoder(16#47#)) OR
 					(reg_q91 AND symb_decoder(16#cc#)) OR
 					(reg_q91 AND symb_decoder(16#af#)) OR
 					(reg_q91 AND symb_decoder(16#d5#)) OR
 					(reg_q91 AND symb_decoder(16#2a#)) OR
 					(reg_q91 AND symb_decoder(16#6d#)) OR
 					(reg_q91 AND symb_decoder(16#c1#)) OR
 					(reg_q91 AND symb_decoder(16#1e#)) OR
 					(reg_q91 AND symb_decoder(16#e8#)) OR
 					(reg_q91 AND symb_decoder(16#dd#)) OR
 					(reg_q91 AND symb_decoder(16#09#)) OR
 					(reg_q91 AND symb_decoder(16#bc#)) OR
 					(reg_q91 AND symb_decoder(16#b5#)) OR
 					(reg_q91 AND symb_decoder(16#db#)) OR
 					(reg_q91 AND symb_decoder(16#f7#)) OR
 					(reg_q91 AND symb_decoder(16#56#)) OR
 					(reg_q91 AND symb_decoder(16#e4#)) OR
 					(reg_q91 AND symb_decoder(16#61#)) OR
 					(reg_q91 AND symb_decoder(16#25#)) OR
 					(reg_q91 AND symb_decoder(16#fd#)) OR
 					(reg_q91 AND symb_decoder(16#80#)) OR
 					(reg_q91 AND symb_decoder(16#12#)) OR
 					(reg_q91 AND symb_decoder(16#06#)) OR
 					(reg_q91 AND symb_decoder(16#4f#)) OR
 					(reg_q91 AND symb_decoder(16#7f#)) OR
 					(reg_q91 AND symb_decoder(16#85#)) OR
 					(reg_q91 AND symb_decoder(16#39#)) OR
 					(reg_q91 AND symb_decoder(16#a4#)) OR
 					(reg_q91 AND symb_decoder(16#f8#)) OR
 					(reg_q91 AND symb_decoder(16#95#)) OR
 					(reg_q91 AND symb_decoder(16#34#)) OR
 					(reg_q91 AND symb_decoder(16#3f#)) OR
 					(reg_q91 AND symb_decoder(16#b7#)) OR
 					(reg_q91 AND symb_decoder(16#10#)) OR
 					(reg_q91 AND symb_decoder(16#cd#)) OR
 					(reg_q91 AND symb_decoder(16#1d#)) OR
 					(reg_q91 AND symb_decoder(16#fe#)) OR
 					(reg_q91 AND symb_decoder(16#31#)) OR
 					(reg_q91 AND symb_decoder(16#16#)) OR
 					(reg_q91 AND symb_decoder(16#20#)) OR
 					(reg_q91 AND symb_decoder(16#b9#)) OR
 					(reg_q91 AND symb_decoder(16#3e#)) OR
 					(reg_q91 AND symb_decoder(16#cb#)) OR
 					(reg_q91 AND symb_decoder(16#de#)) OR
 					(reg_q91 AND symb_decoder(16#d3#)) OR
 					(reg_q91 AND symb_decoder(16#43#)) OR
 					(reg_q91 AND symb_decoder(16#3d#)) OR
 					(reg_q91 AND symb_decoder(16#44#)) OR
 					(reg_q91 AND symb_decoder(16#97#)) OR
 					(reg_q91 AND symb_decoder(16#f2#)) OR
 					(reg_q91 AND symb_decoder(16#5f#)) OR
 					(reg_q91 AND symb_decoder(16#26#)) OR
 					(reg_q91 AND symb_decoder(16#08#)) OR
 					(reg_q91 AND symb_decoder(16#9a#)) OR
 					(reg_q91 AND symb_decoder(16#32#)) OR
 					(reg_q91 AND symb_decoder(16#21#)) OR
 					(reg_q91 AND symb_decoder(16#6a#)) OR
 					(reg_q91 AND symb_decoder(16#ac#)) OR
 					(reg_q91 AND symb_decoder(16#41#)) OR
 					(reg_q91 AND symb_decoder(16#c5#)) OR
 					(reg_q91 AND symb_decoder(16#0f#)) OR
 					(reg_q91 AND symb_decoder(16#74#)) OR
 					(reg_q91 AND symb_decoder(16#8d#)) OR
 					(reg_q91 AND symb_decoder(16#a6#)) OR
 					(reg_q91 AND symb_decoder(16#04#)) OR
 					(reg_q91 AND symb_decoder(16#45#)) OR
 					(reg_q91 AND symb_decoder(16#fb#)) OR
 					(reg_q91 AND symb_decoder(16#0b#)) OR
 					(reg_q91 AND symb_decoder(16#72#)) OR
 					(reg_q91 AND symb_decoder(16#8e#)) OR
 					(reg_q91 AND symb_decoder(16#5a#)) OR
 					(reg_q91 AND symb_decoder(16#60#)) OR
 					(reg_q91 AND symb_decoder(16#84#)) OR
 					(reg_q91 AND symb_decoder(16#27#)) OR
 					(reg_q91 AND symb_decoder(16#d7#)) OR
 					(reg_q91 AND symb_decoder(16#17#)) OR
 					(reg_q91 AND symb_decoder(16#7d#)) OR
 					(reg_q91 AND symb_decoder(16#bd#)) OR
 					(reg_q91 AND symb_decoder(16#4c#)) OR
 					(reg_q91 AND symb_decoder(16#9f#)) OR
 					(reg_q91 AND symb_decoder(16#9d#)) OR
 					(reg_q91 AND symb_decoder(16#0e#)) OR
 					(reg_q91 AND symb_decoder(16#d9#)) OR
 					(reg_q91 AND symb_decoder(16#90#)) OR
 					(reg_q91 AND symb_decoder(16#7c#)) OR
 					(reg_q91 AND symb_decoder(16#65#)) OR
 					(reg_q91 AND symb_decoder(16#3c#)) OR
 					(reg_q91 AND symb_decoder(16#30#)) OR
 					(reg_q91 AND symb_decoder(16#7e#)) OR
 					(reg_q91 AND symb_decoder(16#b8#)) OR
 					(reg_q91 AND symb_decoder(16#70#)) OR
 					(reg_q91 AND symb_decoder(16#b2#)) OR
 					(reg_q91 AND symb_decoder(16#4d#)) OR
 					(reg_q91 AND symb_decoder(16#66#)) OR
 					(reg_q91 AND symb_decoder(16#88#)) OR
 					(reg_q91 AND symb_decoder(16#05#)) OR
 					(reg_q91 AND symb_decoder(16#8a#)) OR
 					(reg_q91 AND symb_decoder(16#c8#)) OR
 					(reg_q91 AND symb_decoder(16#c0#));
reg_q91_init <= '0' ;
	p_reg_q91: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q91 <= reg_q91_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q91 <= reg_q91_init;
        else
          reg_q91 <= reg_q91_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q125_in <= (reg_q123 AND symb_decoder(16#2e#));
reg_q125_init <= '0' ;
	p_reg_q125: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q125 <= reg_q125_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q125 <= reg_q125_init;
        else
          reg_q125 <= reg_q125_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q127_in <= (reg_q125 AND symb_decoder(16#34#)) OR
 					(reg_q125 AND symb_decoder(16#37#)) OR
 					(reg_q125 AND symb_decoder(16#35#)) OR
 					(reg_q125 AND symb_decoder(16#31#)) OR
 					(reg_q125 AND symb_decoder(16#36#)) OR
 					(reg_q125 AND symb_decoder(16#38#)) OR
 					(reg_q125 AND symb_decoder(16#33#)) OR
 					(reg_q125 AND symb_decoder(16#39#)) OR
 					(reg_q125 AND symb_decoder(16#32#)) OR
 					(reg_q125 AND symb_decoder(16#30#)) OR
 					(reg_q127 AND symb_decoder(16#31#)) OR
 					(reg_q127 AND symb_decoder(16#39#)) OR
 					(reg_q127 AND symb_decoder(16#30#)) OR
 					(reg_q127 AND symb_decoder(16#32#)) OR
 					(reg_q127 AND symb_decoder(16#36#)) OR
 					(reg_q127 AND symb_decoder(16#35#)) OR
 					(reg_q127 AND symb_decoder(16#33#)) OR
 					(reg_q127 AND symb_decoder(16#38#)) OR
 					(reg_q127 AND symb_decoder(16#34#)) OR
 					(reg_q127 AND symb_decoder(16#37#));
reg_q127_init <= '0' ;
	p_reg_q127: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q127 <= reg_q127_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q127 <= reg_q127_init;
        else
          reg_q127 <= reg_q127_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q714_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q714 AND symb_decoder(16#a9#)) OR
 					(reg_q714 AND symb_decoder(16#21#)) OR
 					(reg_q714 AND symb_decoder(16#e2#)) OR
 					(reg_q714 AND symb_decoder(16#c9#)) OR
 					(reg_q714 AND symb_decoder(16#ba#)) OR
 					(reg_q714 AND symb_decoder(16#e4#)) OR
 					(reg_q714 AND symb_decoder(16#48#)) OR
 					(reg_q714 AND symb_decoder(16#3f#)) OR
 					(reg_q714 AND symb_decoder(16#d2#)) OR
 					(reg_q714 AND symb_decoder(16#ff#)) OR
 					(reg_q714 AND symb_decoder(16#02#)) OR
 					(reg_q714 AND symb_decoder(16#fd#)) OR
 					(reg_q714 AND symb_decoder(16#60#)) OR
 					(reg_q714 AND symb_decoder(16#ee#)) OR
 					(reg_q714 AND symb_decoder(16#c5#)) OR
 					(reg_q714 AND symb_decoder(16#ae#)) OR
 					(reg_q714 AND symb_decoder(16#97#)) OR
 					(reg_q714 AND symb_decoder(16#16#)) OR
 					(reg_q714 AND symb_decoder(16#fb#)) OR
 					(reg_q714 AND symb_decoder(16#f6#)) OR
 					(reg_q714 AND symb_decoder(16#3c#)) OR
 					(reg_q714 AND symb_decoder(16#bb#)) OR
 					(reg_q714 AND symb_decoder(16#81#)) OR
 					(reg_q714 AND symb_decoder(16#bc#)) OR
 					(reg_q714 AND symb_decoder(16#6a#)) OR
 					(reg_q714 AND symb_decoder(16#04#)) OR
 					(reg_q714 AND symb_decoder(16#8f#)) OR
 					(reg_q714 AND symb_decoder(16#2f#)) OR
 					(reg_q714 AND symb_decoder(16#a8#)) OR
 					(reg_q714 AND symb_decoder(16#fa#)) OR
 					(reg_q714 AND symb_decoder(16#77#)) OR
 					(reg_q714 AND symb_decoder(16#0b#)) OR
 					(reg_q714 AND symb_decoder(16#01#)) OR
 					(reg_q714 AND symb_decoder(16#2c#)) OR
 					(reg_q714 AND symb_decoder(16#f8#)) OR
 					(reg_q714 AND symb_decoder(16#20#)) OR
 					(reg_q714 AND symb_decoder(16#d7#)) OR
 					(reg_q714 AND symb_decoder(16#3b#)) OR
 					(reg_q714 AND symb_decoder(16#33#)) OR
 					(reg_q714 AND symb_decoder(16#de#)) OR
 					(reg_q714 AND symb_decoder(16#43#)) OR
 					(reg_q714 AND symb_decoder(16#f5#)) OR
 					(reg_q714 AND symb_decoder(16#ce#)) OR
 					(reg_q714 AND symb_decoder(16#38#)) OR
 					(reg_q714 AND symb_decoder(16#e8#)) OR
 					(reg_q714 AND symb_decoder(16#89#)) OR
 					(reg_q714 AND symb_decoder(16#e0#)) OR
 					(reg_q714 AND symb_decoder(16#b1#)) OR
 					(reg_q714 AND symb_decoder(16#13#)) OR
 					(reg_q714 AND symb_decoder(16#e7#)) OR
 					(reg_q714 AND symb_decoder(16#dc#)) OR
 					(reg_q714 AND symb_decoder(16#05#)) OR
 					(reg_q714 AND symb_decoder(16#b6#)) OR
 					(reg_q714 AND symb_decoder(16#e3#)) OR
 					(reg_q714 AND symb_decoder(16#39#)) OR
 					(reg_q714 AND symb_decoder(16#df#)) OR
 					(reg_q714 AND symb_decoder(16#a3#)) OR
 					(reg_q714 AND symb_decoder(16#95#)) OR
 					(reg_q714 AND symb_decoder(16#23#)) OR
 					(reg_q714 AND symb_decoder(16#40#)) OR
 					(reg_q714 AND symb_decoder(16#3e#)) OR
 					(reg_q714 AND symb_decoder(16#9b#)) OR
 					(reg_q714 AND symb_decoder(16#fe#)) OR
 					(reg_q714 AND symb_decoder(16#65#)) OR
 					(reg_q714 AND symb_decoder(16#8e#)) OR
 					(reg_q714 AND symb_decoder(16#1b#)) OR
 					(reg_q714 AND symb_decoder(16#4f#)) OR
 					(reg_q714 AND symb_decoder(16#36#)) OR
 					(reg_q714 AND symb_decoder(16#87#)) OR
 					(reg_q714 AND symb_decoder(16#2b#)) OR
 					(reg_q714 AND symb_decoder(16#c7#)) OR
 					(reg_q714 AND symb_decoder(16#32#)) OR
 					(reg_q714 AND symb_decoder(16#19#)) OR
 					(reg_q714 AND symb_decoder(16#4e#)) OR
 					(reg_q714 AND symb_decoder(16#18#)) OR
 					(reg_q714 AND symb_decoder(16#9e#)) OR
 					(reg_q714 AND symb_decoder(16#73#)) OR
 					(reg_q714 AND symb_decoder(16#ea#)) OR
 					(reg_q714 AND symb_decoder(16#42#)) OR
 					(reg_q714 AND symb_decoder(16#0e#)) OR
 					(reg_q714 AND symb_decoder(16#0c#)) OR
 					(reg_q714 AND symb_decoder(16#5a#)) OR
 					(reg_q714 AND symb_decoder(16#08#)) OR
 					(reg_q714 AND symb_decoder(16#98#)) OR
 					(reg_q714 AND symb_decoder(16#5e#)) OR
 					(reg_q714 AND symb_decoder(16#29#)) OR
 					(reg_q714 AND symb_decoder(16#f1#)) OR
 					(reg_q714 AND symb_decoder(16#72#)) OR
 					(reg_q714 AND symb_decoder(16#e1#)) OR
 					(reg_q714 AND symb_decoder(16#d6#)) OR
 					(reg_q714 AND symb_decoder(16#79#)) OR
 					(reg_q714 AND symb_decoder(16#f7#)) OR
 					(reg_q714 AND symb_decoder(16#3d#)) OR
 					(reg_q714 AND symb_decoder(16#db#)) OR
 					(reg_q714 AND symb_decoder(16#ad#)) OR
 					(reg_q714 AND symb_decoder(16#59#)) OR
 					(reg_q714 AND symb_decoder(16#ca#)) OR
 					(reg_q714 AND symb_decoder(16#a0#)) OR
 					(reg_q714 AND symb_decoder(16#58#)) OR
 					(reg_q714 AND symb_decoder(16#0d#)) OR
 					(reg_q714 AND symb_decoder(16#55#)) OR
 					(reg_q714 AND symb_decoder(16#d8#)) OR
 					(reg_q714 AND symb_decoder(16#24#)) OR
 					(reg_q714 AND symb_decoder(16#6d#)) OR
 					(reg_q714 AND symb_decoder(16#4d#)) OR
 					(reg_q714 AND symb_decoder(16#b3#)) OR
 					(reg_q714 AND symb_decoder(16#8c#)) OR
 					(reg_q714 AND symb_decoder(16#7b#)) OR
 					(reg_q714 AND symb_decoder(16#a2#)) OR
 					(reg_q714 AND symb_decoder(16#26#)) OR
 					(reg_q714 AND symb_decoder(16#ef#)) OR
 					(reg_q714 AND symb_decoder(16#4a#)) OR
 					(reg_q714 AND symb_decoder(16#76#)) OR
 					(reg_q714 AND symb_decoder(16#86#)) OR
 					(reg_q714 AND symb_decoder(16#b5#)) OR
 					(reg_q714 AND symb_decoder(16#a5#)) OR
 					(reg_q714 AND symb_decoder(16#2d#)) OR
 					(reg_q714 AND symb_decoder(16#7a#)) OR
 					(reg_q714 AND symb_decoder(16#d1#)) OR
 					(reg_q714 AND symb_decoder(16#d9#)) OR
 					(reg_q714 AND symb_decoder(16#7c#)) OR
 					(reg_q714 AND symb_decoder(16#d3#)) OR
 					(reg_q714 AND symb_decoder(16#e9#)) OR
 					(reg_q714 AND symb_decoder(16#1a#)) OR
 					(reg_q714 AND symb_decoder(16#1d#)) OR
 					(reg_q714 AND symb_decoder(16#4b#)) OR
 					(reg_q714 AND symb_decoder(16#15#)) OR
 					(reg_q714 AND symb_decoder(16#9f#)) OR
 					(reg_q714 AND symb_decoder(16#4c#)) OR
 					(reg_q714 AND symb_decoder(16#c1#)) OR
 					(reg_q714 AND symb_decoder(16#a6#)) OR
 					(reg_q714 AND symb_decoder(16#f9#)) OR
 					(reg_q714 AND symb_decoder(16#61#)) OR
 					(reg_q714 AND symb_decoder(16#c0#)) OR
 					(reg_q714 AND symb_decoder(16#14#)) OR
 					(reg_q714 AND symb_decoder(16#74#)) OR
 					(reg_q714 AND symb_decoder(16#bf#)) OR
 					(reg_q714 AND symb_decoder(16#6c#)) OR
 					(reg_q714 AND symb_decoder(16#cb#)) OR
 					(reg_q714 AND symb_decoder(16#67#)) OR
 					(reg_q714 AND symb_decoder(16#5d#)) OR
 					(reg_q714 AND symb_decoder(16#0a#)) OR
 					(reg_q714 AND symb_decoder(16#66#)) OR
 					(reg_q714 AND symb_decoder(16#2e#)) OR
 					(reg_q714 AND symb_decoder(16#03#)) OR
 					(reg_q714 AND symb_decoder(16#52#)) OR
 					(reg_q714 AND symb_decoder(16#d0#)) OR
 					(reg_q714 AND symb_decoder(16#f2#)) OR
 					(reg_q714 AND symb_decoder(16#9c#)) OR
 					(reg_q714 AND symb_decoder(16#cc#)) OR
 					(reg_q714 AND symb_decoder(16#f0#)) OR
 					(reg_q714 AND symb_decoder(16#5f#)) OR
 					(reg_q714 AND symb_decoder(16#84#)) OR
 					(reg_q714 AND symb_decoder(16#a7#)) OR
 					(reg_q714 AND symb_decoder(16#ab#)) OR
 					(reg_q714 AND symb_decoder(16#da#)) OR
 					(reg_q714 AND symb_decoder(16#c3#)) OR
 					(reg_q714 AND symb_decoder(16#85#)) OR
 					(reg_q714 AND symb_decoder(16#46#)) OR
 					(reg_q714 AND symb_decoder(16#37#)) OR
 					(reg_q714 AND symb_decoder(16#d5#)) OR
 					(reg_q714 AND symb_decoder(16#cf#)) OR
 					(reg_q714 AND symb_decoder(16#b2#)) OR
 					(reg_q714 AND symb_decoder(16#8a#)) OR
 					(reg_q714 AND symb_decoder(16#54#)) OR
 					(reg_q714 AND symb_decoder(16#9d#)) OR
 					(reg_q714 AND symb_decoder(16#e6#)) OR
 					(reg_q714 AND symb_decoder(16#fc#)) OR
 					(reg_q714 AND symb_decoder(16#27#)) OR
 					(reg_q714 AND symb_decoder(16#1c#)) OR
 					(reg_q714 AND symb_decoder(16#99#)) OR
 					(reg_q714 AND symb_decoder(16#22#)) OR
 					(reg_q714 AND symb_decoder(16#ed#)) OR
 					(reg_q714 AND symb_decoder(16#68#)) OR
 					(reg_q714 AND symb_decoder(16#6e#)) OR
 					(reg_q714 AND symb_decoder(16#9a#)) OR
 					(reg_q714 AND symb_decoder(16#dd#)) OR
 					(reg_q714 AND symb_decoder(16#25#)) OR
 					(reg_q714 AND symb_decoder(16#53#)) OR
 					(reg_q714 AND symb_decoder(16#91#)) OR
 					(reg_q714 AND symb_decoder(16#7d#)) OR
 					(reg_q714 AND symb_decoder(16#6f#)) OR
 					(reg_q714 AND symb_decoder(16#f4#)) OR
 					(reg_q714 AND symb_decoder(16#d4#)) OR
 					(reg_q714 AND symb_decoder(16#34#)) OR
 					(reg_q714 AND symb_decoder(16#71#)) OR
 					(reg_q714 AND symb_decoder(16#5c#)) OR
 					(reg_q714 AND symb_decoder(16#10#)) OR
 					(reg_q714 AND symb_decoder(16#82#)) OR
 					(reg_q714 AND symb_decoder(16#a4#)) OR
 					(reg_q714 AND symb_decoder(16#5b#)) OR
 					(reg_q714 AND symb_decoder(16#bd#)) OR
 					(reg_q714 AND symb_decoder(16#8b#)) OR
 					(reg_q714 AND symb_decoder(16#30#)) OR
 					(reg_q714 AND symb_decoder(16#2a#)) OR
 					(reg_q714 AND symb_decoder(16#7f#)) OR
 					(reg_q714 AND symb_decoder(16#75#)) OR
 					(reg_q714 AND symb_decoder(16#eb#)) OR
 					(reg_q714 AND symb_decoder(16#3a#)) OR
 					(reg_q714 AND symb_decoder(16#69#)) OR
 					(reg_q714 AND symb_decoder(16#00#)) OR
 					(reg_q714 AND symb_decoder(16#17#)) OR
 					(reg_q714 AND symb_decoder(16#35#)) OR
 					(reg_q714 AND symb_decoder(16#b9#)) OR
 					(reg_q714 AND symb_decoder(16#6b#)) OR
 					(reg_q714 AND symb_decoder(16#e5#)) OR
 					(reg_q714 AND symb_decoder(16#0f#)) OR
 					(reg_q714 AND symb_decoder(16#63#)) OR
 					(reg_q714 AND symb_decoder(16#78#)) OR
 					(reg_q714 AND symb_decoder(16#90#)) OR
 					(reg_q714 AND symb_decoder(16#c6#)) OR
 					(reg_q714 AND symb_decoder(16#b8#)) OR
 					(reg_q714 AND symb_decoder(16#88#)) OR
 					(reg_q714 AND symb_decoder(16#92#)) OR
 					(reg_q714 AND symb_decoder(16#aa#)) OR
 					(reg_q714 AND symb_decoder(16#12#)) OR
 					(reg_q714 AND symb_decoder(16#70#)) OR
 					(reg_q714 AND symb_decoder(16#80#)) OR
 					(reg_q714 AND symb_decoder(16#b0#)) OR
 					(reg_q714 AND symb_decoder(16#51#)) OR
 					(reg_q714 AND symb_decoder(16#83#)) OR
 					(reg_q714 AND symb_decoder(16#7e#)) OR
 					(reg_q714 AND symb_decoder(16#09#)) OR
 					(reg_q714 AND symb_decoder(16#f3#)) OR
 					(reg_q714 AND symb_decoder(16#b4#)) OR
 					(reg_q714 AND symb_decoder(16#1f#)) OR
 					(reg_q714 AND symb_decoder(16#44#)) OR
 					(reg_q714 AND symb_decoder(16#62#)) OR
 					(reg_q714 AND symb_decoder(16#af#)) OR
 					(reg_q714 AND symb_decoder(16#49#)) OR
 					(reg_q714 AND symb_decoder(16#94#)) OR
 					(reg_q714 AND symb_decoder(16#be#)) OR
 					(reg_q714 AND symb_decoder(16#a1#)) OR
 					(reg_q714 AND symb_decoder(16#06#)) OR
 					(reg_q714 AND symb_decoder(16#31#)) OR
 					(reg_q714 AND symb_decoder(16#45#)) OR
 					(reg_q714 AND symb_decoder(16#c8#)) OR
 					(reg_q714 AND symb_decoder(16#11#)) OR
 					(reg_q714 AND symb_decoder(16#cd#)) OR
 					(reg_q714 AND symb_decoder(16#41#)) OR
 					(reg_q714 AND symb_decoder(16#8d#)) OR
 					(reg_q714 AND symb_decoder(16#96#)) OR
 					(reg_q714 AND symb_decoder(16#28#)) OR
 					(reg_q714 AND symb_decoder(16#64#)) OR
 					(reg_q714 AND symb_decoder(16#56#)) OR
 					(reg_q714 AND symb_decoder(16#50#)) OR
 					(reg_q714 AND symb_decoder(16#ac#)) OR
 					(reg_q714 AND symb_decoder(16#1e#)) OR
 					(reg_q714 AND symb_decoder(16#c4#)) OR
 					(reg_q714 AND symb_decoder(16#47#)) OR
 					(reg_q714 AND symb_decoder(16#07#)) OR
 					(reg_q714 AND symb_decoder(16#57#)) OR
 					(reg_q714 AND symb_decoder(16#c2#)) OR
 					(reg_q714 AND symb_decoder(16#b7#)) OR
 					(reg_q714 AND symb_decoder(16#ec#)) OR
 					(reg_q714 AND symb_decoder(16#93#));
reg_q714_init <= '0' ;
	p_reg_q714: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q714 <= reg_q714_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q714 <= reg_q714_init;
        else
          reg_q714 <= reg_q714_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1544_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1544 AND symb_decoder(16#3e#)) OR
 					(reg_q1544 AND symb_decoder(16#c5#)) OR
 					(reg_q1544 AND symb_decoder(16#f0#)) OR
 					(reg_q1544 AND symb_decoder(16#5d#)) OR
 					(reg_q1544 AND symb_decoder(16#cc#)) OR
 					(reg_q1544 AND symb_decoder(16#51#)) OR
 					(reg_q1544 AND symb_decoder(16#f5#)) OR
 					(reg_q1544 AND symb_decoder(16#b1#)) OR
 					(reg_q1544 AND symb_decoder(16#f8#)) OR
 					(reg_q1544 AND symb_decoder(16#04#)) OR
 					(reg_q1544 AND symb_decoder(16#34#)) OR
 					(reg_q1544 AND symb_decoder(16#35#)) OR
 					(reg_q1544 AND symb_decoder(16#37#)) OR
 					(reg_q1544 AND symb_decoder(16#6c#)) OR
 					(reg_q1544 AND symb_decoder(16#7d#)) OR
 					(reg_q1544 AND symb_decoder(16#30#)) OR
 					(reg_q1544 AND symb_decoder(16#66#)) OR
 					(reg_q1544 AND symb_decoder(16#a6#)) OR
 					(reg_q1544 AND symb_decoder(16#a3#)) OR
 					(reg_q1544 AND symb_decoder(16#2a#)) OR
 					(reg_q1544 AND symb_decoder(16#8d#)) OR
 					(reg_q1544 AND symb_decoder(16#60#)) OR
 					(reg_q1544 AND symb_decoder(16#6a#)) OR
 					(reg_q1544 AND symb_decoder(16#86#)) OR
 					(reg_q1544 AND symb_decoder(16#ad#)) OR
 					(reg_q1544 AND symb_decoder(16#62#)) OR
 					(reg_q1544 AND symb_decoder(16#f1#)) OR
 					(reg_q1544 AND symb_decoder(16#07#)) OR
 					(reg_q1544 AND symb_decoder(16#ed#)) OR
 					(reg_q1544 AND symb_decoder(16#58#)) OR
 					(reg_q1544 AND symb_decoder(16#f4#)) OR
 					(reg_q1544 AND symb_decoder(16#f3#)) OR
 					(reg_q1544 AND symb_decoder(16#e9#)) OR
 					(reg_q1544 AND symb_decoder(16#83#)) OR
 					(reg_q1544 AND symb_decoder(16#8e#)) OR
 					(reg_q1544 AND symb_decoder(16#bc#)) OR
 					(reg_q1544 AND symb_decoder(16#72#)) OR
 					(reg_q1544 AND symb_decoder(16#87#)) OR
 					(reg_q1544 AND symb_decoder(16#7e#)) OR
 					(reg_q1544 AND symb_decoder(16#c2#)) OR
 					(reg_q1544 AND symb_decoder(16#45#)) OR
 					(reg_q1544 AND symb_decoder(16#96#)) OR
 					(reg_q1544 AND symb_decoder(16#2d#)) OR
 					(reg_q1544 AND symb_decoder(16#47#)) OR
 					(reg_q1544 AND symb_decoder(16#1d#)) OR
 					(reg_q1544 AND symb_decoder(16#95#)) OR
 					(reg_q1544 AND symb_decoder(16#52#)) OR
 					(reg_q1544 AND symb_decoder(16#20#)) OR
 					(reg_q1544 AND symb_decoder(16#9f#)) OR
 					(reg_q1544 AND symb_decoder(16#0b#)) OR
 					(reg_q1544 AND symb_decoder(16#cb#)) OR
 					(reg_q1544 AND symb_decoder(16#59#)) OR
 					(reg_q1544 AND symb_decoder(16#6f#)) OR
 					(reg_q1544 AND symb_decoder(16#7c#)) OR
 					(reg_q1544 AND symb_decoder(16#1f#)) OR
 					(reg_q1544 AND symb_decoder(16#4e#)) OR
 					(reg_q1544 AND symb_decoder(16#3d#)) OR
 					(reg_q1544 AND symb_decoder(16#e3#)) OR
 					(reg_q1544 AND symb_decoder(16#94#)) OR
 					(reg_q1544 AND symb_decoder(16#0c#)) OR
 					(reg_q1544 AND symb_decoder(16#64#)) OR
 					(reg_q1544 AND symb_decoder(16#dc#)) OR
 					(reg_q1544 AND symb_decoder(16#fe#)) OR
 					(reg_q1544 AND symb_decoder(16#d9#)) OR
 					(reg_q1544 AND symb_decoder(16#db#)) OR
 					(reg_q1544 AND symb_decoder(16#e4#)) OR
 					(reg_q1544 AND symb_decoder(16#d8#)) OR
 					(reg_q1544 AND symb_decoder(16#e8#)) OR
 					(reg_q1544 AND symb_decoder(16#49#)) OR
 					(reg_q1544 AND symb_decoder(16#11#)) OR
 					(reg_q1544 AND symb_decoder(16#39#)) OR
 					(reg_q1544 AND symb_decoder(16#c9#)) OR
 					(reg_q1544 AND symb_decoder(16#c7#)) OR
 					(reg_q1544 AND symb_decoder(16#f9#)) OR
 					(reg_q1544 AND symb_decoder(16#d0#)) OR
 					(reg_q1544 AND symb_decoder(16#0a#)) OR
 					(reg_q1544 AND symb_decoder(16#68#)) OR
 					(reg_q1544 AND symb_decoder(16#32#)) OR
 					(reg_q1544 AND symb_decoder(16#fa#)) OR
 					(reg_q1544 AND symb_decoder(16#6b#)) OR
 					(reg_q1544 AND symb_decoder(16#0e#)) OR
 					(reg_q1544 AND symb_decoder(16#16#)) OR
 					(reg_q1544 AND symb_decoder(16#14#)) OR
 					(reg_q1544 AND symb_decoder(16#84#)) OR
 					(reg_q1544 AND symb_decoder(16#df#)) OR
 					(reg_q1544 AND symb_decoder(16#2b#)) OR
 					(reg_q1544 AND symb_decoder(16#70#)) OR
 					(reg_q1544 AND symb_decoder(16#0f#)) OR
 					(reg_q1544 AND symb_decoder(16#ea#)) OR
 					(reg_q1544 AND symb_decoder(16#e7#)) OR
 					(reg_q1544 AND symb_decoder(16#63#)) OR
 					(reg_q1544 AND symb_decoder(16#57#)) OR
 					(reg_q1544 AND symb_decoder(16#8c#)) OR
 					(reg_q1544 AND symb_decoder(16#79#)) OR
 					(reg_q1544 AND symb_decoder(16#f7#)) OR
 					(reg_q1544 AND symb_decoder(16#69#)) OR
 					(reg_q1544 AND symb_decoder(16#15#)) OR
 					(reg_q1544 AND symb_decoder(16#c3#)) OR
 					(reg_q1544 AND symb_decoder(16#ac#)) OR
 					(reg_q1544 AND symb_decoder(16#e1#)) OR
 					(reg_q1544 AND symb_decoder(16#ff#)) OR
 					(reg_q1544 AND symb_decoder(16#42#)) OR
 					(reg_q1544 AND symb_decoder(16#12#)) OR
 					(reg_q1544 AND symb_decoder(16#08#)) OR
 					(reg_q1544 AND symb_decoder(16#61#)) OR
 					(reg_q1544 AND symb_decoder(16#e5#)) OR
 					(reg_q1544 AND symb_decoder(16#28#)) OR
 					(reg_q1544 AND symb_decoder(16#5a#)) OR
 					(reg_q1544 AND symb_decoder(16#2c#)) OR
 					(reg_q1544 AND symb_decoder(16#c4#)) OR
 					(reg_q1544 AND symb_decoder(16#75#)) OR
 					(reg_q1544 AND symb_decoder(16#d2#)) OR
 					(reg_q1544 AND symb_decoder(16#55#)) OR
 					(reg_q1544 AND symb_decoder(16#c8#)) OR
 					(reg_q1544 AND symb_decoder(16#89#)) OR
 					(reg_q1544 AND symb_decoder(16#25#)) OR
 					(reg_q1544 AND symb_decoder(16#43#)) OR
 					(reg_q1544 AND symb_decoder(16#4f#)) OR
 					(reg_q1544 AND symb_decoder(16#02#)) OR
 					(reg_q1544 AND symb_decoder(16#c0#)) OR
 					(reg_q1544 AND symb_decoder(16#b5#)) OR
 					(reg_q1544 AND symb_decoder(16#71#)) OR
 					(reg_q1544 AND symb_decoder(16#ce#)) OR
 					(reg_q1544 AND symb_decoder(16#74#)) OR
 					(reg_q1544 AND symb_decoder(16#8a#)) OR
 					(reg_q1544 AND symb_decoder(16#2f#)) OR
 					(reg_q1544 AND symb_decoder(16#f2#)) OR
 					(reg_q1544 AND symb_decoder(16#d4#)) OR
 					(reg_q1544 AND symb_decoder(16#03#)) OR
 					(reg_q1544 AND symb_decoder(16#26#)) OR
 					(reg_q1544 AND symb_decoder(16#01#)) OR
 					(reg_q1544 AND symb_decoder(16#8f#)) OR
 					(reg_q1544 AND symb_decoder(16#3b#)) OR
 					(reg_q1544 AND symb_decoder(16#1a#)) OR
 					(reg_q1544 AND symb_decoder(16#ae#)) OR
 					(reg_q1544 AND symb_decoder(16#e0#)) OR
 					(reg_q1544 AND symb_decoder(16#5e#)) OR
 					(reg_q1544 AND symb_decoder(16#d1#)) OR
 					(reg_q1544 AND symb_decoder(16#ba#)) OR
 					(reg_q1544 AND symb_decoder(16#48#)) OR
 					(reg_q1544 AND symb_decoder(16#fb#)) OR
 					(reg_q1544 AND symb_decoder(16#23#)) OR
 					(reg_q1544 AND symb_decoder(16#31#)) OR
 					(reg_q1544 AND symb_decoder(16#50#)) OR
 					(reg_q1544 AND symb_decoder(16#33#)) OR
 					(reg_q1544 AND symb_decoder(16#73#)) OR
 					(reg_q1544 AND symb_decoder(16#1c#)) OR
 					(reg_q1544 AND symb_decoder(16#5f#)) OR
 					(reg_q1544 AND symb_decoder(16#81#)) OR
 					(reg_q1544 AND symb_decoder(16#56#)) OR
 					(reg_q1544 AND symb_decoder(16#3f#)) OR
 					(reg_q1544 AND symb_decoder(16#dd#)) OR
 					(reg_q1544 AND symb_decoder(16#88#)) OR
 					(reg_q1544 AND symb_decoder(16#ee#)) OR
 					(reg_q1544 AND symb_decoder(16#a4#)) OR
 					(reg_q1544 AND symb_decoder(16#b2#)) OR
 					(reg_q1544 AND symb_decoder(16#c6#)) OR
 					(reg_q1544 AND symb_decoder(16#e6#)) OR
 					(reg_q1544 AND symb_decoder(16#a7#)) OR
 					(reg_q1544 AND symb_decoder(16#6d#)) OR
 					(reg_q1544 AND symb_decoder(16#7b#)) OR
 					(reg_q1544 AND symb_decoder(16#7a#)) OR
 					(reg_q1544 AND symb_decoder(16#cf#)) OR
 					(reg_q1544 AND symb_decoder(16#65#)) OR
 					(reg_q1544 AND symb_decoder(16#91#)) OR
 					(reg_q1544 AND symb_decoder(16#76#)) OR
 					(reg_q1544 AND symb_decoder(16#3c#)) OR
 					(reg_q1544 AND symb_decoder(16#bf#)) OR
 					(reg_q1544 AND symb_decoder(16#be#)) OR
 					(reg_q1544 AND symb_decoder(16#53#)) OR
 					(reg_q1544 AND symb_decoder(16#36#)) OR
 					(reg_q1544 AND symb_decoder(16#78#)) OR
 					(reg_q1544 AND symb_decoder(16#00#)) OR
 					(reg_q1544 AND symb_decoder(16#1e#)) OR
 					(reg_q1544 AND symb_decoder(16#0d#)) OR
 					(reg_q1544 AND symb_decoder(16#ab#)) OR
 					(reg_q1544 AND symb_decoder(16#09#)) OR
 					(reg_q1544 AND symb_decoder(16#80#)) OR
 					(reg_q1544 AND symb_decoder(16#3a#)) OR
 					(reg_q1544 AND symb_decoder(16#9d#)) OR
 					(reg_q1544 AND symb_decoder(16#98#)) OR
 					(reg_q1544 AND symb_decoder(16#ef#)) OR
 					(reg_q1544 AND symb_decoder(16#f6#)) OR
 					(reg_q1544 AND symb_decoder(16#ec#)) OR
 					(reg_q1544 AND symb_decoder(16#de#)) OR
 					(reg_q1544 AND symb_decoder(16#d5#)) OR
 					(reg_q1544 AND symb_decoder(16#b8#)) OR
 					(reg_q1544 AND symb_decoder(16#13#)) OR
 					(reg_q1544 AND symb_decoder(16#5c#)) OR
 					(reg_q1544 AND symb_decoder(16#d6#)) OR
 					(reg_q1544 AND symb_decoder(16#c1#)) OR
 					(reg_q1544 AND symb_decoder(16#85#)) OR
 					(reg_q1544 AND symb_decoder(16#67#)) OR
 					(reg_q1544 AND symb_decoder(16#fc#)) OR
 					(reg_q1544 AND symb_decoder(16#17#)) OR
 					(reg_q1544 AND symb_decoder(16#27#)) OR
 					(reg_q1544 AND symb_decoder(16#5b#)) OR
 					(reg_q1544 AND symb_decoder(16#d7#)) OR
 					(reg_q1544 AND symb_decoder(16#a0#)) OR
 					(reg_q1544 AND symb_decoder(16#b9#)) OR
 					(reg_q1544 AND symb_decoder(16#54#)) OR
 					(reg_q1544 AND symb_decoder(16#90#)) OR
 					(reg_q1544 AND symb_decoder(16#41#)) OR
 					(reg_q1544 AND symb_decoder(16#a5#)) OR
 					(reg_q1544 AND symb_decoder(16#b4#)) OR
 					(reg_q1544 AND symb_decoder(16#38#)) OR
 					(reg_q1544 AND symb_decoder(16#21#)) OR
 					(reg_q1544 AND symb_decoder(16#bb#)) OR
 					(reg_q1544 AND symb_decoder(16#9a#)) OR
 					(reg_q1544 AND symb_decoder(16#b0#)) OR
 					(reg_q1544 AND symb_decoder(16#05#)) OR
 					(reg_q1544 AND symb_decoder(16#eb#)) OR
 					(reg_q1544 AND symb_decoder(16#8b#)) OR
 					(reg_q1544 AND symb_decoder(16#97#)) OR
 					(reg_q1544 AND symb_decoder(16#da#)) OR
 					(reg_q1544 AND symb_decoder(16#aa#)) OR
 					(reg_q1544 AND symb_decoder(16#a9#)) OR
 					(reg_q1544 AND symb_decoder(16#af#)) OR
 					(reg_q1544 AND symb_decoder(16#24#)) OR
 					(reg_q1544 AND symb_decoder(16#fd#)) OR
 					(reg_q1544 AND symb_decoder(16#a2#)) OR
 					(reg_q1544 AND symb_decoder(16#19#)) OR
 					(reg_q1544 AND symb_decoder(16#44#)) OR
 					(reg_q1544 AND symb_decoder(16#9b#)) OR
 					(reg_q1544 AND symb_decoder(16#6e#)) OR
 					(reg_q1544 AND symb_decoder(16#4d#)) OR
 					(reg_q1544 AND symb_decoder(16#cd#)) OR
 					(reg_q1544 AND symb_decoder(16#b6#)) OR
 					(reg_q1544 AND symb_decoder(16#40#)) OR
 					(reg_q1544 AND symb_decoder(16#b7#)) OR
 					(reg_q1544 AND symb_decoder(16#22#)) OR
 					(reg_q1544 AND symb_decoder(16#99#)) OR
 					(reg_q1544 AND symb_decoder(16#b3#)) OR
 					(reg_q1544 AND symb_decoder(16#4b#)) OR
 					(reg_q1544 AND symb_decoder(16#bd#)) OR
 					(reg_q1544 AND symb_decoder(16#2e#)) OR
 					(reg_q1544 AND symb_decoder(16#9e#)) OR
 					(reg_q1544 AND symb_decoder(16#4c#)) OR
 					(reg_q1544 AND symb_decoder(16#4a#)) OR
 					(reg_q1544 AND symb_decoder(16#82#)) OR
 					(reg_q1544 AND symb_decoder(16#92#)) OR
 					(reg_q1544 AND symb_decoder(16#ca#)) OR
 					(reg_q1544 AND symb_decoder(16#46#)) OR
 					(reg_q1544 AND symb_decoder(16#7f#)) OR
 					(reg_q1544 AND symb_decoder(16#9c#)) OR
 					(reg_q1544 AND symb_decoder(16#d3#)) OR
 					(reg_q1544 AND symb_decoder(16#10#)) OR
 					(reg_q1544 AND symb_decoder(16#e2#)) OR
 					(reg_q1544 AND symb_decoder(16#93#)) OR
 					(reg_q1544 AND symb_decoder(16#a8#)) OR
 					(reg_q1544 AND symb_decoder(16#1b#)) OR
 					(reg_q1544 AND symb_decoder(16#29#)) OR
 					(reg_q1544 AND symb_decoder(16#77#)) OR
 					(reg_q1544 AND symb_decoder(16#06#)) OR
 					(reg_q1544 AND symb_decoder(16#a1#)) OR
 					(reg_q1544 AND symb_decoder(16#18#));
reg_q1544_init <= '0' ;
	p_reg_q1544: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1544 <= reg_q1544_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1544 <= reg_q1544_init;
        else
          reg_q1544 <= reg_q1544_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1928_in <= (reg_q1926 AND symb_decoder(16#62#)) OR
 					(reg_q1926 AND symb_decoder(16#42#));
reg_q1928_init <= '0' ;
	p_reg_q1928: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1928 <= reg_q1928_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1928 <= reg_q1928_init;
        else
          reg_q1928 <= reg_q1928_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1930_in <= (reg_q1928 AND symb_decoder(16#61#)) OR
 					(reg_q1928 AND symb_decoder(16#41#));
reg_q1930_init <= '0' ;
	p_reg_q1930: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1930 <= reg_q1930_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1930 <= reg_q1930_init;
        else
          reg_q1930 <= reg_q1930_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2533_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2533 AND symb_decoder(16#68#)) OR
 					(reg_q2533 AND symb_decoder(16#b0#)) OR
 					(reg_q2533 AND symb_decoder(16#29#)) OR
 					(reg_q2533 AND symb_decoder(16#f9#)) OR
 					(reg_q2533 AND symb_decoder(16#41#)) OR
 					(reg_q2533 AND symb_decoder(16#3a#)) OR
 					(reg_q2533 AND symb_decoder(16#d7#)) OR
 					(reg_q2533 AND symb_decoder(16#b4#)) OR
 					(reg_q2533 AND symb_decoder(16#2b#)) OR
 					(reg_q2533 AND symb_decoder(16#ac#)) OR
 					(reg_q2533 AND symb_decoder(16#fb#)) OR
 					(reg_q2533 AND symb_decoder(16#5e#)) OR
 					(reg_q2533 AND symb_decoder(16#db#)) OR
 					(reg_q2533 AND symb_decoder(16#cb#)) OR
 					(reg_q2533 AND symb_decoder(16#12#)) OR
 					(reg_q2533 AND symb_decoder(16#72#)) OR
 					(reg_q2533 AND symb_decoder(16#f4#)) OR
 					(reg_q2533 AND symb_decoder(16#1f#)) OR
 					(reg_q2533 AND symb_decoder(16#76#)) OR
 					(reg_q2533 AND symb_decoder(16#01#)) OR
 					(reg_q2533 AND symb_decoder(16#75#)) OR
 					(reg_q2533 AND symb_decoder(16#a3#)) OR
 					(reg_q2533 AND symb_decoder(16#44#)) OR
 					(reg_q2533 AND symb_decoder(16#70#)) OR
 					(reg_q2533 AND symb_decoder(16#a2#)) OR
 					(reg_q2533 AND symb_decoder(16#9d#)) OR
 					(reg_q2533 AND symb_decoder(16#c7#)) OR
 					(reg_q2533 AND symb_decoder(16#50#)) OR
 					(reg_q2533 AND symb_decoder(16#81#)) OR
 					(reg_q2533 AND symb_decoder(16#d5#)) OR
 					(reg_q2533 AND symb_decoder(16#bc#)) OR
 					(reg_q2533 AND symb_decoder(16#b9#)) OR
 					(reg_q2533 AND symb_decoder(16#e8#)) OR
 					(reg_q2533 AND symb_decoder(16#88#)) OR
 					(reg_q2533 AND symb_decoder(16#2a#)) OR
 					(reg_q2533 AND symb_decoder(16#de#)) OR
 					(reg_q2533 AND symb_decoder(16#cc#)) OR
 					(reg_q2533 AND symb_decoder(16#1e#)) OR
 					(reg_q2533 AND symb_decoder(16#8e#)) OR
 					(reg_q2533 AND symb_decoder(16#11#)) OR
 					(reg_q2533 AND symb_decoder(16#1a#)) OR
 					(reg_q2533 AND symb_decoder(16#fc#)) OR
 					(reg_q2533 AND symb_decoder(16#74#)) OR
 					(reg_q2533 AND symb_decoder(16#24#)) OR
 					(reg_q2533 AND symb_decoder(16#55#)) OR
 					(reg_q2533 AND symb_decoder(16#64#)) OR
 					(reg_q2533 AND symb_decoder(16#8d#)) OR
 					(reg_q2533 AND symb_decoder(16#91#)) OR
 					(reg_q2533 AND symb_decoder(16#b8#)) OR
 					(reg_q2533 AND symb_decoder(16#0e#)) OR
 					(reg_q2533 AND symb_decoder(16#d3#)) OR
 					(reg_q2533 AND symb_decoder(16#c0#)) OR
 					(reg_q2533 AND symb_decoder(16#5b#)) OR
 					(reg_q2533 AND symb_decoder(16#a9#)) OR
 					(reg_q2533 AND symb_decoder(16#27#)) OR
 					(reg_q2533 AND symb_decoder(16#49#)) OR
 					(reg_q2533 AND symb_decoder(16#84#)) OR
 					(reg_q2533 AND symb_decoder(16#6c#)) OR
 					(reg_q2533 AND symb_decoder(16#59#)) OR
 					(reg_q2533 AND symb_decoder(16#f5#)) OR
 					(reg_q2533 AND symb_decoder(16#3d#)) OR
 					(reg_q2533 AND symb_decoder(16#10#)) OR
 					(reg_q2533 AND symb_decoder(16#a8#)) OR
 					(reg_q2533 AND symb_decoder(16#04#)) OR
 					(reg_q2533 AND symb_decoder(16#0a#)) OR
 					(reg_q2533 AND symb_decoder(16#9a#)) OR
 					(reg_q2533 AND symb_decoder(16#85#)) OR
 					(reg_q2533 AND symb_decoder(16#2f#)) OR
 					(reg_q2533 AND symb_decoder(16#05#)) OR
 					(reg_q2533 AND symb_decoder(16#39#)) OR
 					(reg_q2533 AND symb_decoder(16#e5#)) OR
 					(reg_q2533 AND symb_decoder(16#0c#)) OR
 					(reg_q2533 AND symb_decoder(16#4f#)) OR
 					(reg_q2533 AND symb_decoder(16#ba#)) OR
 					(reg_q2533 AND symb_decoder(16#dd#)) OR
 					(reg_q2533 AND symb_decoder(16#ec#)) OR
 					(reg_q2533 AND symb_decoder(16#0b#)) OR
 					(reg_q2533 AND symb_decoder(16#52#)) OR
 					(reg_q2533 AND symb_decoder(16#cd#)) OR
 					(reg_q2533 AND symb_decoder(16#02#)) OR
 					(reg_q2533 AND symb_decoder(16#2e#)) OR
 					(reg_q2533 AND symb_decoder(16#fa#)) OR
 					(reg_q2533 AND symb_decoder(16#fe#)) OR
 					(reg_q2533 AND symb_decoder(16#40#)) OR
 					(reg_q2533 AND symb_decoder(16#a6#)) OR
 					(reg_q2533 AND symb_decoder(16#6d#)) OR
 					(reg_q2533 AND symb_decoder(16#7f#)) OR
 					(reg_q2533 AND symb_decoder(16#ce#)) OR
 					(reg_q2533 AND symb_decoder(16#e6#)) OR
 					(reg_q2533 AND symb_decoder(16#da#)) OR
 					(reg_q2533 AND symb_decoder(16#08#)) OR
 					(reg_q2533 AND symb_decoder(16#45#)) OR
 					(reg_q2533 AND symb_decoder(16#c9#)) OR
 					(reg_q2533 AND symb_decoder(16#a0#)) OR
 					(reg_q2533 AND symb_decoder(16#f8#)) OR
 					(reg_q2533 AND symb_decoder(16#eb#)) OR
 					(reg_q2533 AND symb_decoder(16#e1#)) OR
 					(reg_q2533 AND symb_decoder(16#4a#)) OR
 					(reg_q2533 AND symb_decoder(16#0f#)) OR
 					(reg_q2533 AND symb_decoder(16#f6#)) OR
 					(reg_q2533 AND symb_decoder(16#b3#)) OR
 					(reg_q2533 AND symb_decoder(16#d6#)) OR
 					(reg_q2533 AND symb_decoder(16#7c#)) OR
 					(reg_q2533 AND symb_decoder(16#c6#)) OR
 					(reg_q2533 AND symb_decoder(16#c2#)) OR
 					(reg_q2533 AND symb_decoder(16#b1#)) OR
 					(reg_q2533 AND symb_decoder(16#58#)) OR
 					(reg_q2533 AND symb_decoder(16#3b#)) OR
 					(reg_q2533 AND symb_decoder(16#53#)) OR
 					(reg_q2533 AND symb_decoder(16#54#)) OR
 					(reg_q2533 AND symb_decoder(16#92#)) OR
 					(reg_q2533 AND symb_decoder(16#03#)) OR
 					(reg_q2533 AND symb_decoder(16#51#)) OR
 					(reg_q2533 AND symb_decoder(16#c3#)) OR
 					(reg_q2533 AND symb_decoder(16#5a#)) OR
 					(reg_q2533 AND symb_decoder(16#83#)) OR
 					(reg_q2533 AND symb_decoder(16#20#)) OR
 					(reg_q2533 AND symb_decoder(16#19#)) OR
 					(reg_q2533 AND symb_decoder(16#e0#)) OR
 					(reg_q2533 AND symb_decoder(16#13#)) OR
 					(reg_q2533 AND symb_decoder(16#6e#)) OR
 					(reg_q2533 AND symb_decoder(16#96#)) OR
 					(reg_q2533 AND symb_decoder(16#a7#)) OR
 					(reg_q2533 AND symb_decoder(16#18#)) OR
 					(reg_q2533 AND symb_decoder(16#aa#)) OR
 					(reg_q2533 AND symb_decoder(16#78#)) OR
 					(reg_q2533 AND symb_decoder(16#8f#)) OR
 					(reg_q2533 AND symb_decoder(16#bd#)) OR
 					(reg_q2533 AND symb_decoder(16#32#)) OR
 					(reg_q2533 AND symb_decoder(16#4e#)) OR
 					(reg_q2533 AND symb_decoder(16#86#)) OR
 					(reg_q2533 AND symb_decoder(16#d2#)) OR
 					(reg_q2533 AND symb_decoder(16#43#)) OR
 					(reg_q2533 AND symb_decoder(16#fd#)) OR
 					(reg_q2533 AND symb_decoder(16#2d#)) OR
 					(reg_q2533 AND symb_decoder(16#a4#)) OR
 					(reg_q2533 AND symb_decoder(16#a1#)) OR
 					(reg_q2533 AND symb_decoder(16#46#)) OR
 					(reg_q2533 AND symb_decoder(16#57#)) OR
 					(reg_q2533 AND symb_decoder(16#b7#)) OR
 					(reg_q2533 AND symb_decoder(16#7e#)) OR
 					(reg_q2533 AND symb_decoder(16#65#)) OR
 					(reg_q2533 AND symb_decoder(16#e3#)) OR
 					(reg_q2533 AND symb_decoder(16#cf#)) OR
 					(reg_q2533 AND symb_decoder(16#9e#)) OR
 					(reg_q2533 AND symb_decoder(16#80#)) OR
 					(reg_q2533 AND symb_decoder(16#93#)) OR
 					(reg_q2533 AND symb_decoder(16#31#)) OR
 					(reg_q2533 AND symb_decoder(16#98#)) OR
 					(reg_q2533 AND symb_decoder(16#e7#)) OR
 					(reg_q2533 AND symb_decoder(16#d9#)) OR
 					(reg_q2533 AND symb_decoder(16#73#)) OR
 					(reg_q2533 AND symb_decoder(16#48#)) OR
 					(reg_q2533 AND symb_decoder(16#c8#)) OR
 					(reg_q2533 AND symb_decoder(16#9f#)) OR
 					(reg_q2533 AND symb_decoder(16#f1#)) OR
 					(reg_q2533 AND symb_decoder(16#b2#)) OR
 					(reg_q2533 AND symb_decoder(16#17#)) OR
 					(reg_q2533 AND symb_decoder(16#90#)) OR
 					(reg_q2533 AND symb_decoder(16#b5#)) OR
 					(reg_q2533 AND symb_decoder(16#06#)) OR
 					(reg_q2533 AND symb_decoder(16#8b#)) OR
 					(reg_q2533 AND symb_decoder(16#ff#)) OR
 					(reg_q2533 AND symb_decoder(16#4c#)) OR
 					(reg_q2533 AND symb_decoder(16#0d#)) OR
 					(reg_q2533 AND symb_decoder(16#dc#)) OR
 					(reg_q2533 AND symb_decoder(16#47#)) OR
 					(reg_q2533 AND symb_decoder(16#28#)) OR
 					(reg_q2533 AND symb_decoder(16#1b#)) OR
 					(reg_q2533 AND symb_decoder(16#af#)) OR
 					(reg_q2533 AND symb_decoder(16#99#)) OR
 					(reg_q2533 AND symb_decoder(16#f0#)) OR
 					(reg_q2533 AND symb_decoder(16#25#)) OR
 					(reg_q2533 AND symb_decoder(16#35#)) OR
 					(reg_q2533 AND symb_decoder(16#a5#)) OR
 					(reg_q2533 AND symb_decoder(16#71#)) OR
 					(reg_q2533 AND symb_decoder(16#5f#)) OR
 					(reg_q2533 AND symb_decoder(16#d4#)) OR
 					(reg_q2533 AND symb_decoder(16#82#)) OR
 					(reg_q2533 AND symb_decoder(16#00#)) OR
 					(reg_q2533 AND symb_decoder(16#60#)) OR
 					(reg_q2533 AND symb_decoder(16#97#)) OR
 					(reg_q2533 AND symb_decoder(16#33#)) OR
 					(reg_q2533 AND symb_decoder(16#ae#)) OR
 					(reg_q2533 AND symb_decoder(16#16#)) OR
 					(reg_q2533 AND symb_decoder(16#21#)) OR
 					(reg_q2533 AND symb_decoder(16#9c#)) OR
 					(reg_q2533 AND symb_decoder(16#6a#)) OR
 					(reg_q2533 AND symb_decoder(16#4d#)) OR
 					(reg_q2533 AND symb_decoder(16#34#)) OR
 					(reg_q2533 AND symb_decoder(16#36#)) OR
 					(reg_q2533 AND symb_decoder(16#94#)) OR
 					(reg_q2533 AND symb_decoder(16#c1#)) OR
 					(reg_q2533 AND symb_decoder(16#62#)) OR
 					(reg_q2533 AND symb_decoder(16#b6#)) OR
 					(reg_q2533 AND symb_decoder(16#ef#)) OR
 					(reg_q2533 AND symb_decoder(16#ca#)) OR
 					(reg_q2533 AND symb_decoder(16#2c#)) OR
 					(reg_q2533 AND symb_decoder(16#07#)) OR
 					(reg_q2533 AND symb_decoder(16#d1#)) OR
 					(reg_q2533 AND symb_decoder(16#77#)) OR
 					(reg_q2533 AND symb_decoder(16#7a#)) OR
 					(reg_q2533 AND symb_decoder(16#5d#)) OR
 					(reg_q2533 AND symb_decoder(16#42#)) OR
 					(reg_q2533 AND symb_decoder(16#f7#)) OR
 					(reg_q2533 AND symb_decoder(16#c4#)) OR
 					(reg_q2533 AND symb_decoder(16#bb#)) OR
 					(reg_q2533 AND symb_decoder(16#c5#)) OR
 					(reg_q2533 AND symb_decoder(16#1d#)) OR
 					(reg_q2533 AND symb_decoder(16#79#)) OR
 					(reg_q2533 AND symb_decoder(16#7d#)) OR
 					(reg_q2533 AND symb_decoder(16#9b#)) OR
 					(reg_q2533 AND symb_decoder(16#df#)) OR
 					(reg_q2533 AND symb_decoder(16#ed#)) OR
 					(reg_q2533 AND symb_decoder(16#89#)) OR
 					(reg_q2533 AND symb_decoder(16#5c#)) OR
 					(reg_q2533 AND symb_decoder(16#14#)) OR
 					(reg_q2533 AND symb_decoder(16#f3#)) OR
 					(reg_q2533 AND symb_decoder(16#8c#)) OR
 					(reg_q2533 AND symb_decoder(16#95#)) OR
 					(reg_q2533 AND symb_decoder(16#4b#)) OR
 					(reg_q2533 AND symb_decoder(16#26#)) OR
 					(reg_q2533 AND symb_decoder(16#67#)) OR
 					(reg_q2533 AND symb_decoder(16#ea#)) OR
 					(reg_q2533 AND symb_decoder(16#d0#)) OR
 					(reg_q2533 AND symb_decoder(16#6b#)) OR
 					(reg_q2533 AND symb_decoder(16#3c#)) OR
 					(reg_q2533 AND symb_decoder(16#e9#)) OR
 					(reg_q2533 AND symb_decoder(16#7b#)) OR
 					(reg_q2533 AND symb_decoder(16#3e#)) OR
 					(reg_q2533 AND symb_decoder(16#e2#)) OR
 					(reg_q2533 AND symb_decoder(16#56#)) OR
 					(reg_q2533 AND symb_decoder(16#e4#)) OR
 					(reg_q2533 AND symb_decoder(16#87#)) OR
 					(reg_q2533 AND symb_decoder(16#37#)) OR
 					(reg_q2533 AND symb_decoder(16#38#)) OR
 					(reg_q2533 AND symb_decoder(16#15#)) OR
 					(reg_q2533 AND symb_decoder(16#30#)) OR
 					(reg_q2533 AND symb_decoder(16#d8#)) OR
 					(reg_q2533 AND symb_decoder(16#be#)) OR
 					(reg_q2533 AND symb_decoder(16#61#)) OR
 					(reg_q2533 AND symb_decoder(16#ee#)) OR
 					(reg_q2533 AND symb_decoder(16#3f#)) OR
 					(reg_q2533 AND symb_decoder(16#8a#)) OR
 					(reg_q2533 AND symb_decoder(16#63#)) OR
 					(reg_q2533 AND symb_decoder(16#ad#)) OR
 					(reg_q2533 AND symb_decoder(16#ab#)) OR
 					(reg_q2533 AND symb_decoder(16#69#)) OR
 					(reg_q2533 AND symb_decoder(16#23#)) OR
 					(reg_q2533 AND symb_decoder(16#66#)) OR
 					(reg_q2533 AND symb_decoder(16#6f#)) OR
 					(reg_q2533 AND symb_decoder(16#22#)) OR
 					(reg_q2533 AND symb_decoder(16#1c#)) OR
 					(reg_q2533 AND symb_decoder(16#bf#)) OR
 					(reg_q2533 AND symb_decoder(16#f2#)) OR
 					(reg_q2533 AND symb_decoder(16#09#));
reg_q2533_init <= '0' ;
	p_reg_q2533: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2533 <= reg_q2533_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2533 <= reg_q2533_init;
        else
          reg_q2533 <= reg_q2533_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1742_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1742 AND symb_decoder(16#b8#)) OR
 					(reg_q1742 AND symb_decoder(16#00#)) OR
 					(reg_q1742 AND symb_decoder(16#42#)) OR
 					(reg_q1742 AND symb_decoder(16#a5#)) OR
 					(reg_q1742 AND symb_decoder(16#54#)) OR
 					(reg_q1742 AND symb_decoder(16#b3#)) OR
 					(reg_q1742 AND symb_decoder(16#da#)) OR
 					(reg_q1742 AND symb_decoder(16#d9#)) OR
 					(reg_q1742 AND symb_decoder(16#de#)) OR
 					(reg_q1742 AND symb_decoder(16#21#)) OR
 					(reg_q1742 AND symb_decoder(16#d1#)) OR
 					(reg_q1742 AND symb_decoder(16#0b#)) OR
 					(reg_q1742 AND symb_decoder(16#8d#)) OR
 					(reg_q1742 AND symb_decoder(16#62#)) OR
 					(reg_q1742 AND symb_decoder(16#f4#)) OR
 					(reg_q1742 AND symb_decoder(16#c7#)) OR
 					(reg_q1742 AND symb_decoder(16#f5#)) OR
 					(reg_q1742 AND symb_decoder(16#51#)) OR
 					(reg_q1742 AND symb_decoder(16#94#)) OR
 					(reg_q1742 AND symb_decoder(16#2a#)) OR
 					(reg_q1742 AND symb_decoder(16#eb#)) OR
 					(reg_q1742 AND symb_decoder(16#96#)) OR
 					(reg_q1742 AND symb_decoder(16#27#)) OR
 					(reg_q1742 AND symb_decoder(16#ed#)) OR
 					(reg_q1742 AND symb_decoder(16#7a#)) OR
 					(reg_q1742 AND symb_decoder(16#09#)) OR
 					(reg_q1742 AND symb_decoder(16#e5#)) OR
 					(reg_q1742 AND symb_decoder(16#66#)) OR
 					(reg_q1742 AND symb_decoder(16#aa#)) OR
 					(reg_q1742 AND symb_decoder(16#82#)) OR
 					(reg_q1742 AND symb_decoder(16#d3#)) OR
 					(reg_q1742 AND symb_decoder(16#ae#)) OR
 					(reg_q1742 AND symb_decoder(16#98#)) OR
 					(reg_q1742 AND symb_decoder(16#0e#)) OR
 					(reg_q1742 AND symb_decoder(16#30#)) OR
 					(reg_q1742 AND symb_decoder(16#46#)) OR
 					(reg_q1742 AND symb_decoder(16#0f#)) OR
 					(reg_q1742 AND symb_decoder(16#1c#)) OR
 					(reg_q1742 AND symb_decoder(16#97#)) OR
 					(reg_q1742 AND symb_decoder(16#ef#)) OR
 					(reg_q1742 AND symb_decoder(16#a1#)) OR
 					(reg_q1742 AND symb_decoder(16#e1#)) OR
 					(reg_q1742 AND symb_decoder(16#5d#)) OR
 					(reg_q1742 AND symb_decoder(16#9d#)) OR
 					(reg_q1742 AND symb_decoder(16#45#)) OR
 					(reg_q1742 AND symb_decoder(16#4b#)) OR
 					(reg_q1742 AND symb_decoder(16#cd#)) OR
 					(reg_q1742 AND symb_decoder(16#20#)) OR
 					(reg_q1742 AND symb_decoder(16#93#)) OR
 					(reg_q1742 AND symb_decoder(16#f0#)) OR
 					(reg_q1742 AND symb_decoder(16#fe#)) OR
 					(reg_q1742 AND symb_decoder(16#11#)) OR
 					(reg_q1742 AND symb_decoder(16#63#)) OR
 					(reg_q1742 AND symb_decoder(16#e7#)) OR
 					(reg_q1742 AND symb_decoder(16#c1#)) OR
 					(reg_q1742 AND symb_decoder(16#d6#)) OR
 					(reg_q1742 AND symb_decoder(16#06#)) OR
 					(reg_q1742 AND symb_decoder(16#e9#)) OR
 					(reg_q1742 AND symb_decoder(16#47#)) OR
 					(reg_q1742 AND symb_decoder(16#80#)) OR
 					(reg_q1742 AND symb_decoder(16#d2#)) OR
 					(reg_q1742 AND symb_decoder(16#f8#)) OR
 					(reg_q1742 AND symb_decoder(16#ce#)) OR
 					(reg_q1742 AND symb_decoder(16#48#)) OR
 					(reg_q1742 AND symb_decoder(16#75#)) OR
 					(reg_q1742 AND symb_decoder(16#d5#)) OR
 					(reg_q1742 AND symb_decoder(16#3d#)) OR
 					(reg_q1742 AND symb_decoder(16#76#)) OR
 					(reg_q1742 AND symb_decoder(16#9f#)) OR
 					(reg_q1742 AND symb_decoder(16#9a#)) OR
 					(reg_q1742 AND symb_decoder(16#7c#)) OR
 					(reg_q1742 AND symb_decoder(16#1a#)) OR
 					(reg_q1742 AND symb_decoder(16#b0#)) OR
 					(reg_q1742 AND symb_decoder(16#65#)) OR
 					(reg_q1742 AND symb_decoder(16#33#)) OR
 					(reg_q1742 AND symb_decoder(16#18#)) OR
 					(reg_q1742 AND symb_decoder(16#43#)) OR
 					(reg_q1742 AND symb_decoder(16#d0#)) OR
 					(reg_q1742 AND symb_decoder(16#77#)) OR
 					(reg_q1742 AND symb_decoder(16#c6#)) OR
 					(reg_q1742 AND symb_decoder(16#0d#)) OR
 					(reg_q1742 AND symb_decoder(16#5a#)) OR
 					(reg_q1742 AND symb_decoder(16#dd#)) OR
 					(reg_q1742 AND symb_decoder(16#bd#)) OR
 					(reg_q1742 AND symb_decoder(16#67#)) OR
 					(reg_q1742 AND symb_decoder(16#83#)) OR
 					(reg_q1742 AND symb_decoder(16#b6#)) OR
 					(reg_q1742 AND symb_decoder(16#8b#)) OR
 					(reg_q1742 AND symb_decoder(16#87#)) OR
 					(reg_q1742 AND symb_decoder(16#02#)) OR
 					(reg_q1742 AND symb_decoder(16#d4#)) OR
 					(reg_q1742 AND symb_decoder(16#ff#)) OR
 					(reg_q1742 AND symb_decoder(16#40#)) OR
 					(reg_q1742 AND symb_decoder(16#74#)) OR
 					(reg_q1742 AND symb_decoder(16#8f#)) OR
 					(reg_q1742 AND symb_decoder(16#6d#)) OR
 					(reg_q1742 AND symb_decoder(16#ab#)) OR
 					(reg_q1742 AND symb_decoder(16#10#)) OR
 					(reg_q1742 AND symb_decoder(16#4f#)) OR
 					(reg_q1742 AND symb_decoder(16#19#)) OR
 					(reg_q1742 AND symb_decoder(16#69#)) OR
 					(reg_q1742 AND symb_decoder(16#4e#)) OR
 					(reg_q1742 AND symb_decoder(16#58#)) OR
 					(reg_q1742 AND symb_decoder(16#68#)) OR
 					(reg_q1742 AND symb_decoder(16#ea#)) OR
 					(reg_q1742 AND symb_decoder(16#64#)) OR
 					(reg_q1742 AND symb_decoder(16#39#)) OR
 					(reg_q1742 AND symb_decoder(16#c9#)) OR
 					(reg_q1742 AND symb_decoder(16#0a#)) OR
 					(reg_q1742 AND symb_decoder(16#2b#)) OR
 					(reg_q1742 AND symb_decoder(16#56#)) OR
 					(reg_q1742 AND symb_decoder(16#72#)) OR
 					(reg_q1742 AND symb_decoder(16#2e#)) OR
 					(reg_q1742 AND symb_decoder(16#4d#)) OR
 					(reg_q1742 AND symb_decoder(16#6a#)) OR
 					(reg_q1742 AND symb_decoder(16#bc#)) OR
 					(reg_q1742 AND symb_decoder(16#57#)) OR
 					(reg_q1742 AND symb_decoder(16#9e#)) OR
 					(reg_q1742 AND symb_decoder(16#0c#)) OR
 					(reg_q1742 AND symb_decoder(16#3b#)) OR
 					(reg_q1742 AND symb_decoder(16#ba#)) OR
 					(reg_q1742 AND symb_decoder(16#fd#)) OR
 					(reg_q1742 AND symb_decoder(16#95#)) OR
 					(reg_q1742 AND symb_decoder(16#a0#)) OR
 					(reg_q1742 AND symb_decoder(16#b1#)) OR
 					(reg_q1742 AND symb_decoder(16#7e#)) OR
 					(reg_q1742 AND symb_decoder(16#e8#)) OR
 					(reg_q1742 AND symb_decoder(16#23#)) OR
 					(reg_q1742 AND symb_decoder(16#37#)) OR
 					(reg_q1742 AND symb_decoder(16#84#)) OR
 					(reg_q1742 AND symb_decoder(16#73#)) OR
 					(reg_q1742 AND symb_decoder(16#b2#)) OR
 					(reg_q1742 AND symb_decoder(16#5c#)) OR
 					(reg_q1742 AND symb_decoder(16#16#)) OR
 					(reg_q1742 AND symb_decoder(16#5b#)) OR
 					(reg_q1742 AND symb_decoder(16#a3#)) OR
 					(reg_q1742 AND symb_decoder(16#fb#)) OR
 					(reg_q1742 AND symb_decoder(16#cb#)) OR
 					(reg_q1742 AND symb_decoder(16#ee#)) OR
 					(reg_q1742 AND symb_decoder(16#81#)) OR
 					(reg_q1742 AND symb_decoder(16#a7#)) OR
 					(reg_q1742 AND symb_decoder(16#b4#)) OR
 					(reg_q1742 AND symb_decoder(16#c5#)) OR
 					(reg_q1742 AND symb_decoder(16#f6#)) OR
 					(reg_q1742 AND symb_decoder(16#e6#)) OR
 					(reg_q1742 AND symb_decoder(16#c4#)) OR
 					(reg_q1742 AND symb_decoder(16#22#)) OR
 					(reg_q1742 AND symb_decoder(16#13#)) OR
 					(reg_q1742 AND symb_decoder(16#df#)) OR
 					(reg_q1742 AND symb_decoder(16#24#)) OR
 					(reg_q1742 AND symb_decoder(16#d7#)) OR
 					(reg_q1742 AND symb_decoder(16#c8#)) OR
 					(reg_q1742 AND symb_decoder(16#c0#)) OR
 					(reg_q1742 AND symb_decoder(16#ca#)) OR
 					(reg_q1742 AND symb_decoder(16#79#)) OR
 					(reg_q1742 AND symb_decoder(16#36#)) OR
 					(reg_q1742 AND symb_decoder(16#4a#)) OR
 					(reg_q1742 AND symb_decoder(16#99#)) OR
 					(reg_q1742 AND symb_decoder(16#f3#)) OR
 					(reg_q1742 AND symb_decoder(16#85#)) OR
 					(reg_q1742 AND symb_decoder(16#2c#)) OR
 					(reg_q1742 AND symb_decoder(16#53#)) OR
 					(reg_q1742 AND symb_decoder(16#a4#)) OR
 					(reg_q1742 AND symb_decoder(16#b5#)) OR
 					(reg_q1742 AND symb_decoder(16#32#)) OR
 					(reg_q1742 AND symb_decoder(16#01#)) OR
 					(reg_q1742 AND symb_decoder(16#41#)) OR
 					(reg_q1742 AND symb_decoder(16#a8#)) OR
 					(reg_q1742 AND symb_decoder(16#50#)) OR
 					(reg_q1742 AND symb_decoder(16#dc#)) OR
 					(reg_q1742 AND symb_decoder(16#7f#)) OR
 					(reg_q1742 AND symb_decoder(16#14#)) OR
 					(reg_q1742 AND symb_decoder(16#fa#)) OR
 					(reg_q1742 AND symb_decoder(16#90#)) OR
 					(reg_q1742 AND symb_decoder(16#38#)) OR
 					(reg_q1742 AND symb_decoder(16#29#)) OR
 					(reg_q1742 AND symb_decoder(16#71#)) OR
 					(reg_q1742 AND symb_decoder(16#5e#)) OR
 					(reg_q1742 AND symb_decoder(16#3a#)) OR
 					(reg_q1742 AND symb_decoder(16#3f#)) OR
 					(reg_q1742 AND symb_decoder(16#b7#)) OR
 					(reg_q1742 AND symb_decoder(16#55#)) OR
 					(reg_q1742 AND symb_decoder(16#9b#)) OR
 					(reg_q1742 AND symb_decoder(16#6c#)) OR
 					(reg_q1742 AND symb_decoder(16#9c#)) OR
 					(reg_q1742 AND symb_decoder(16#52#)) OR
 					(reg_q1742 AND symb_decoder(16#f1#)) OR
 					(reg_q1742 AND symb_decoder(16#c2#)) OR
 					(reg_q1742 AND symb_decoder(16#25#)) OR
 					(reg_q1742 AND symb_decoder(16#a9#)) OR
 					(reg_q1742 AND symb_decoder(16#d8#)) OR
 					(reg_q1742 AND symb_decoder(16#70#)) OR
 					(reg_q1742 AND symb_decoder(16#e0#)) OR
 					(reg_q1742 AND symb_decoder(16#fc#)) OR
 					(reg_q1742 AND symb_decoder(16#7d#)) OR
 					(reg_q1742 AND symb_decoder(16#28#)) OR
 					(reg_q1742 AND symb_decoder(16#e2#)) OR
 					(reg_q1742 AND symb_decoder(16#8c#)) OR
 					(reg_q1742 AND symb_decoder(16#8e#)) OR
 					(reg_q1742 AND symb_decoder(16#b9#)) OR
 					(reg_q1742 AND symb_decoder(16#08#)) OR
 					(reg_q1742 AND symb_decoder(16#5f#)) OR
 					(reg_q1742 AND symb_decoder(16#c3#)) OR
 					(reg_q1742 AND symb_decoder(16#3e#)) OR
 					(reg_q1742 AND symb_decoder(16#cc#)) OR
 					(reg_q1742 AND symb_decoder(16#ad#)) OR
 					(reg_q1742 AND symb_decoder(16#2d#)) OR
 					(reg_q1742 AND symb_decoder(16#34#)) OR
 					(reg_q1742 AND symb_decoder(16#78#)) OR
 					(reg_q1742 AND symb_decoder(16#92#)) OR
 					(reg_q1742 AND symb_decoder(16#af#)) OR
 					(reg_q1742 AND symb_decoder(16#6b#)) OR
 					(reg_q1742 AND symb_decoder(16#ac#)) OR
 					(reg_q1742 AND symb_decoder(16#35#)) OR
 					(reg_q1742 AND symb_decoder(16#f7#)) OR
 					(reg_q1742 AND symb_decoder(16#6f#)) OR
 					(reg_q1742 AND symb_decoder(16#12#)) OR
 					(reg_q1742 AND symb_decoder(16#1d#)) OR
 					(reg_q1742 AND symb_decoder(16#bb#)) OR
 					(reg_q1742 AND symb_decoder(16#4c#)) OR
 					(reg_q1742 AND symb_decoder(16#31#)) OR
 					(reg_q1742 AND symb_decoder(16#17#)) OR
 					(reg_q1742 AND symb_decoder(16#f2#)) OR
 					(reg_q1742 AND symb_decoder(16#3c#)) OR
 					(reg_q1742 AND symb_decoder(16#ec#)) OR
 					(reg_q1742 AND symb_decoder(16#26#)) OR
 					(reg_q1742 AND symb_decoder(16#44#)) OR
 					(reg_q1742 AND symb_decoder(16#1f#)) OR
 					(reg_q1742 AND symb_decoder(16#cf#)) OR
 					(reg_q1742 AND symb_decoder(16#bf#)) OR
 					(reg_q1742 AND symb_decoder(16#a6#)) OR
 					(reg_q1742 AND symb_decoder(16#db#)) OR
 					(reg_q1742 AND symb_decoder(16#7b#)) OR
 					(reg_q1742 AND symb_decoder(16#89#)) OR
 					(reg_q1742 AND symb_decoder(16#e4#)) OR
 					(reg_q1742 AND symb_decoder(16#8a#)) OR
 					(reg_q1742 AND symb_decoder(16#88#)) OR
 					(reg_q1742 AND symb_decoder(16#be#)) OR
 					(reg_q1742 AND symb_decoder(16#a2#)) OR
 					(reg_q1742 AND symb_decoder(16#61#)) OR
 					(reg_q1742 AND symb_decoder(16#1b#)) OR
 					(reg_q1742 AND symb_decoder(16#60#)) OR
 					(reg_q1742 AND symb_decoder(16#03#)) OR
 					(reg_q1742 AND symb_decoder(16#07#)) OR
 					(reg_q1742 AND symb_decoder(16#59#)) OR
 					(reg_q1742 AND symb_decoder(16#91#)) OR
 					(reg_q1742 AND symb_decoder(16#f9#)) OR
 					(reg_q1742 AND symb_decoder(16#15#)) OR
 					(reg_q1742 AND symb_decoder(16#e3#)) OR
 					(reg_q1742 AND symb_decoder(16#04#)) OR
 					(reg_q1742 AND symb_decoder(16#1e#)) OR
 					(reg_q1742 AND symb_decoder(16#86#)) OR
 					(reg_q1742 AND symb_decoder(16#6e#)) OR
 					(reg_q1742 AND symb_decoder(16#2f#)) OR
 					(reg_q1742 AND symb_decoder(16#05#)) OR
 					(reg_q1742 AND symb_decoder(16#49#));
reg_q1742_init <= '0' ;
	p_reg_q1742: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1742 <= reg_q1742_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1742 <= reg_q1742_init;
        else
          reg_q1742 <= reg_q1742_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1668_in <= (reg_q1666 AND symb_decoder(16#2e#));
reg_q1668_init <= '0' ;
	p_reg_q1668: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1668 <= reg_q1668_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1668 <= reg_q1668_init;
        else
          reg_q1668 <= reg_q1668_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1670_in <= (reg_q1668 AND symb_decoder(16#34#)) OR
 					(reg_q1668 AND symb_decoder(16#39#)) OR
 					(reg_q1668 AND symb_decoder(16#36#)) OR
 					(reg_q1668 AND symb_decoder(16#35#)) OR
 					(reg_q1668 AND symb_decoder(16#37#)) OR
 					(reg_q1668 AND symb_decoder(16#32#)) OR
 					(reg_q1668 AND symb_decoder(16#31#)) OR
 					(reg_q1668 AND symb_decoder(16#38#)) OR
 					(reg_q1668 AND symb_decoder(16#33#)) OR
 					(reg_q1668 AND symb_decoder(16#30#)) OR
 					(reg_q1670 AND symb_decoder(16#34#)) OR
 					(reg_q1670 AND symb_decoder(16#39#)) OR
 					(reg_q1670 AND symb_decoder(16#36#)) OR
 					(reg_q1670 AND symb_decoder(16#33#)) OR
 					(reg_q1670 AND symb_decoder(16#31#)) OR
 					(reg_q1670 AND symb_decoder(16#38#)) OR
 					(reg_q1670 AND symb_decoder(16#32#)) OR
 					(reg_q1670 AND symb_decoder(16#35#)) OR
 					(reg_q1670 AND symb_decoder(16#37#)) OR
 					(reg_q1670 AND symb_decoder(16#30#));
reg_q1670_init <= '0' ;
	p_reg_q1670: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1670 <= reg_q1670_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1670 <= reg_q1670_init;
        else
          reg_q1670 <= reg_q1670_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1050_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1050 AND symb_decoder(16#4d#)) OR
 					(reg_q1050 AND symb_decoder(16#06#)) OR
 					(reg_q1050 AND symb_decoder(16#8c#)) OR
 					(reg_q1050 AND symb_decoder(16#82#)) OR
 					(reg_q1050 AND symb_decoder(16#2a#)) OR
 					(reg_q1050 AND symb_decoder(16#1d#)) OR
 					(reg_q1050 AND symb_decoder(16#7a#)) OR
 					(reg_q1050 AND symb_decoder(16#42#)) OR
 					(reg_q1050 AND symb_decoder(16#72#)) OR
 					(reg_q1050 AND symb_decoder(16#ac#)) OR
 					(reg_q1050 AND symb_decoder(16#39#)) OR
 					(reg_q1050 AND symb_decoder(16#b6#)) OR
 					(reg_q1050 AND symb_decoder(16#8d#)) OR
 					(reg_q1050 AND symb_decoder(16#3e#)) OR
 					(reg_q1050 AND symb_decoder(16#ec#)) OR
 					(reg_q1050 AND symb_decoder(16#e4#)) OR
 					(reg_q1050 AND symb_decoder(16#1f#)) OR
 					(reg_q1050 AND symb_decoder(16#14#)) OR
 					(reg_q1050 AND symb_decoder(16#ef#)) OR
 					(reg_q1050 AND symb_decoder(16#d7#)) OR
 					(reg_q1050 AND symb_decoder(16#ee#)) OR
 					(reg_q1050 AND symb_decoder(16#92#)) OR
 					(reg_q1050 AND symb_decoder(16#01#)) OR
 					(reg_q1050 AND symb_decoder(16#17#)) OR
 					(reg_q1050 AND symb_decoder(16#f7#)) OR
 					(reg_q1050 AND symb_decoder(16#28#)) OR
 					(reg_q1050 AND symb_decoder(16#35#)) OR
 					(reg_q1050 AND symb_decoder(16#9d#)) OR
 					(reg_q1050 AND symb_decoder(16#b0#)) OR
 					(reg_q1050 AND symb_decoder(16#80#)) OR
 					(reg_q1050 AND symb_decoder(16#b4#)) OR
 					(reg_q1050 AND symb_decoder(16#2b#)) OR
 					(reg_q1050 AND symb_decoder(16#a3#)) OR
 					(reg_q1050 AND symb_decoder(16#3b#)) OR
 					(reg_q1050 AND symb_decoder(16#10#)) OR
 					(reg_q1050 AND symb_decoder(16#68#)) OR
 					(reg_q1050 AND symb_decoder(16#0d#)) OR
 					(reg_q1050 AND symb_decoder(16#dc#)) OR
 					(reg_q1050 AND symb_decoder(16#f2#)) OR
 					(reg_q1050 AND symb_decoder(16#5b#)) OR
 					(reg_q1050 AND symb_decoder(16#43#)) OR
 					(reg_q1050 AND symb_decoder(16#33#)) OR
 					(reg_q1050 AND symb_decoder(16#1e#)) OR
 					(reg_q1050 AND symb_decoder(16#bd#)) OR
 					(reg_q1050 AND symb_decoder(16#47#)) OR
 					(reg_q1050 AND symb_decoder(16#f1#)) OR
 					(reg_q1050 AND symb_decoder(16#ce#)) OR
 					(reg_q1050 AND symb_decoder(16#5f#)) OR
 					(reg_q1050 AND symb_decoder(16#de#)) OR
 					(reg_q1050 AND symb_decoder(16#61#)) OR
 					(reg_q1050 AND symb_decoder(16#7f#)) OR
 					(reg_q1050 AND symb_decoder(16#a9#)) OR
 					(reg_q1050 AND symb_decoder(16#ba#)) OR
 					(reg_q1050 AND symb_decoder(16#fd#)) OR
 					(reg_q1050 AND symb_decoder(16#e2#)) OR
 					(reg_q1050 AND symb_decoder(16#0a#)) OR
 					(reg_q1050 AND symb_decoder(16#b3#)) OR
 					(reg_q1050 AND symb_decoder(16#8e#)) OR
 					(reg_q1050 AND symb_decoder(16#bc#)) OR
 					(reg_q1050 AND symb_decoder(16#d0#)) OR
 					(reg_q1050 AND symb_decoder(16#ff#)) OR
 					(reg_q1050 AND symb_decoder(16#3c#)) OR
 					(reg_q1050 AND symb_decoder(16#24#)) OR
 					(reg_q1050 AND symb_decoder(16#5a#)) OR
 					(reg_q1050 AND symb_decoder(16#58#)) OR
 					(reg_q1050 AND symb_decoder(16#e9#)) OR
 					(reg_q1050 AND symb_decoder(16#f4#)) OR
 					(reg_q1050 AND symb_decoder(16#55#)) OR
 					(reg_q1050 AND symb_decoder(16#73#)) OR
 					(reg_q1050 AND symb_decoder(16#63#)) OR
 					(reg_q1050 AND symb_decoder(16#be#)) OR
 					(reg_q1050 AND symb_decoder(16#a7#)) OR
 					(reg_q1050 AND symb_decoder(16#20#)) OR
 					(reg_q1050 AND symb_decoder(16#27#)) OR
 					(reg_q1050 AND symb_decoder(16#8b#)) OR
 					(reg_q1050 AND symb_decoder(16#52#)) OR
 					(reg_q1050 AND symb_decoder(16#ea#)) OR
 					(reg_q1050 AND symb_decoder(16#c9#)) OR
 					(reg_q1050 AND symb_decoder(16#09#)) OR
 					(reg_q1050 AND symb_decoder(16#75#)) OR
 					(reg_q1050 AND symb_decoder(16#81#)) OR
 					(reg_q1050 AND symb_decoder(16#49#)) OR
 					(reg_q1050 AND symb_decoder(16#d1#)) OR
 					(reg_q1050 AND symb_decoder(16#31#)) OR
 					(reg_q1050 AND symb_decoder(16#a0#)) OR
 					(reg_q1050 AND symb_decoder(16#46#)) OR
 					(reg_q1050 AND symb_decoder(16#4f#)) OR
 					(reg_q1050 AND symb_decoder(16#2f#)) OR
 					(reg_q1050 AND symb_decoder(16#1b#)) OR
 					(reg_q1050 AND symb_decoder(16#05#)) OR
 					(reg_q1050 AND symb_decoder(16#f5#)) OR
 					(reg_q1050 AND symb_decoder(16#c5#)) OR
 					(reg_q1050 AND symb_decoder(16#6a#)) OR
 					(reg_q1050 AND symb_decoder(16#a5#)) OR
 					(reg_q1050 AND symb_decoder(16#16#)) OR
 					(reg_q1050 AND symb_decoder(16#4a#)) OR
 					(reg_q1050 AND symb_decoder(16#76#)) OR
 					(reg_q1050 AND symb_decoder(16#38#)) OR
 					(reg_q1050 AND symb_decoder(16#78#)) OR
 					(reg_q1050 AND symb_decoder(16#bf#)) OR
 					(reg_q1050 AND symb_decoder(16#8a#)) OR
 					(reg_q1050 AND symb_decoder(16#23#)) OR
 					(reg_q1050 AND symb_decoder(16#90#)) OR
 					(reg_q1050 AND symb_decoder(16#d5#)) OR
 					(reg_q1050 AND symb_decoder(16#3d#)) OR
 					(reg_q1050 AND symb_decoder(16#e5#)) OR
 					(reg_q1050 AND symb_decoder(16#03#)) OR
 					(reg_q1050 AND symb_decoder(16#a4#)) OR
 					(reg_q1050 AND symb_decoder(16#04#)) OR
 					(reg_q1050 AND symb_decoder(16#4b#)) OR
 					(reg_q1050 AND symb_decoder(16#93#)) OR
 					(reg_q1050 AND symb_decoder(16#0c#)) OR
 					(reg_q1050 AND symb_decoder(16#21#)) OR
 					(reg_q1050 AND symb_decoder(16#12#)) OR
 					(reg_q1050 AND symb_decoder(16#a1#)) OR
 					(reg_q1050 AND symb_decoder(16#66#)) OR
 					(reg_q1050 AND symb_decoder(16#d9#)) OR
 					(reg_q1050 AND symb_decoder(16#cd#)) OR
 					(reg_q1050 AND symb_decoder(16#74#)) OR
 					(reg_q1050 AND symb_decoder(16#84#)) OR
 					(reg_q1050 AND symb_decoder(16#4c#)) OR
 					(reg_q1050 AND symb_decoder(16#c2#)) OR
 					(reg_q1050 AND symb_decoder(16#96#)) OR
 					(reg_q1050 AND symb_decoder(16#57#)) OR
 					(reg_q1050 AND symb_decoder(16#3f#)) OR
 					(reg_q1050 AND symb_decoder(16#88#)) OR
 					(reg_q1050 AND symb_decoder(16#19#)) OR
 					(reg_q1050 AND symb_decoder(16#7e#)) OR
 					(reg_q1050 AND symb_decoder(16#4e#)) OR
 					(reg_q1050 AND symb_decoder(16#e1#)) OR
 					(reg_q1050 AND symb_decoder(16#ed#)) OR
 					(reg_q1050 AND symb_decoder(16#dd#)) OR
 					(reg_q1050 AND symb_decoder(16#fc#)) OR
 					(reg_q1050 AND symb_decoder(16#af#)) OR
 					(reg_q1050 AND symb_decoder(16#3a#)) OR
 					(reg_q1050 AND symb_decoder(16#a2#)) OR
 					(reg_q1050 AND symb_decoder(16#30#)) OR
 					(reg_q1050 AND symb_decoder(16#aa#)) OR
 					(reg_q1050 AND symb_decoder(16#50#)) OR
 					(reg_q1050 AND symb_decoder(16#fb#)) OR
 					(reg_q1050 AND symb_decoder(16#94#)) OR
 					(reg_q1050 AND symb_decoder(16#11#)) OR
 					(reg_q1050 AND symb_decoder(16#d6#)) OR
 					(reg_q1050 AND symb_decoder(16#9f#)) OR
 					(reg_q1050 AND symb_decoder(16#e7#)) OR
 					(reg_q1050 AND symb_decoder(16#45#)) OR
 					(reg_q1050 AND symb_decoder(16#c4#)) OR
 					(reg_q1050 AND symb_decoder(16#6f#)) OR
 					(reg_q1050 AND symb_decoder(16#b2#)) OR
 					(reg_q1050 AND symb_decoder(16#ab#)) OR
 					(reg_q1050 AND symb_decoder(16#cf#)) OR
 					(reg_q1050 AND symb_decoder(16#d2#)) OR
 					(reg_q1050 AND symb_decoder(16#51#)) OR
 					(reg_q1050 AND symb_decoder(16#48#)) OR
 					(reg_q1050 AND symb_decoder(16#f8#)) OR
 					(reg_q1050 AND symb_decoder(16#5d#)) OR
 					(reg_q1050 AND symb_decoder(16#36#)) OR
 					(reg_q1050 AND symb_decoder(16#c0#)) OR
 					(reg_q1050 AND symb_decoder(16#b7#)) OR
 					(reg_q1050 AND symb_decoder(16#99#)) OR
 					(reg_q1050 AND symb_decoder(16#9b#)) OR
 					(reg_q1050 AND symb_decoder(16#c3#)) OR
 					(reg_q1050 AND symb_decoder(16#f9#)) OR
 					(reg_q1050 AND symb_decoder(16#69#)) OR
 					(reg_q1050 AND symb_decoder(16#41#)) OR
 					(reg_q1050 AND symb_decoder(16#53#)) OR
 					(reg_q1050 AND symb_decoder(16#86#)) OR
 					(reg_q1050 AND symb_decoder(16#d3#)) OR
 					(reg_q1050 AND symb_decoder(16#83#)) OR
 					(reg_q1050 AND symb_decoder(16#8f#)) OR
 					(reg_q1050 AND symb_decoder(16#f6#)) OR
 					(reg_q1050 AND symb_decoder(16#ae#)) OR
 					(reg_q1050 AND symb_decoder(16#5e#)) OR
 					(reg_q1050 AND symb_decoder(16#d4#)) OR
 					(reg_q1050 AND symb_decoder(16#26#)) OR
 					(reg_q1050 AND symb_decoder(16#fe#)) OR
 					(reg_q1050 AND symb_decoder(16#db#)) OR
 					(reg_q1050 AND symb_decoder(16#1a#)) OR
 					(reg_q1050 AND symb_decoder(16#08#)) OR
 					(reg_q1050 AND symb_decoder(16#a6#)) OR
 					(reg_q1050 AND symb_decoder(16#da#)) OR
 					(reg_q1050 AND symb_decoder(16#b1#)) OR
 					(reg_q1050 AND symb_decoder(16#71#)) OR
 					(reg_q1050 AND symb_decoder(16#bb#)) OR
 					(reg_q1050 AND symb_decoder(16#0e#)) OR
 					(reg_q1050 AND symb_decoder(16#25#)) OR
 					(reg_q1050 AND symb_decoder(16#60#)) OR
 					(reg_q1050 AND symb_decoder(16#cb#)) OR
 					(reg_q1050 AND symb_decoder(16#18#)) OR
 					(reg_q1050 AND symb_decoder(16#2e#)) OR
 					(reg_q1050 AND symb_decoder(16#13#)) OR
 					(reg_q1050 AND symb_decoder(16#40#)) OR
 					(reg_q1050 AND symb_decoder(16#98#)) OR
 					(reg_q1050 AND symb_decoder(16#e8#)) OR
 					(reg_q1050 AND symb_decoder(16#f3#)) OR
 					(reg_q1050 AND symb_decoder(16#c7#)) OR
 					(reg_q1050 AND symb_decoder(16#7b#)) OR
 					(reg_q1050 AND symb_decoder(16#a8#)) OR
 					(reg_q1050 AND symb_decoder(16#54#)) OR
 					(reg_q1050 AND symb_decoder(16#22#)) OR
 					(reg_q1050 AND symb_decoder(16#1c#)) OR
 					(reg_q1050 AND symb_decoder(16#15#)) OR
 					(reg_q1050 AND symb_decoder(16#32#)) OR
 					(reg_q1050 AND symb_decoder(16#79#)) OR
 					(reg_q1050 AND symb_decoder(16#b5#)) OR
 					(reg_q1050 AND symb_decoder(16#02#)) OR
 					(reg_q1050 AND symb_decoder(16#c8#)) OR
 					(reg_q1050 AND symb_decoder(16#77#)) OR
 					(reg_q1050 AND symb_decoder(16#c6#)) OR
 					(reg_q1050 AND symb_decoder(16#7d#)) OR
 					(reg_q1050 AND symb_decoder(16#df#)) OR
 					(reg_q1050 AND symb_decoder(16#70#)) OR
 					(reg_q1050 AND symb_decoder(16#e0#)) OR
 					(reg_q1050 AND symb_decoder(16#87#)) OR
 					(reg_q1050 AND symb_decoder(16#cc#)) OR
 					(reg_q1050 AND symb_decoder(16#67#)) OR
 					(reg_q1050 AND symb_decoder(16#29#)) OR
 					(reg_q1050 AND symb_decoder(16#ad#)) OR
 					(reg_q1050 AND symb_decoder(16#97#)) OR
 					(reg_q1050 AND symb_decoder(16#e3#)) OR
 					(reg_q1050 AND symb_decoder(16#6b#)) OR
 					(reg_q1050 AND symb_decoder(16#0f#)) OR
 					(reg_q1050 AND symb_decoder(16#ca#)) OR
 					(reg_q1050 AND symb_decoder(16#0b#)) OR
 					(reg_q1050 AND symb_decoder(16#85#)) OR
 					(reg_q1050 AND symb_decoder(16#c1#)) OR
 					(reg_q1050 AND symb_decoder(16#2c#)) OR
 					(reg_q1050 AND symb_decoder(16#37#)) OR
 					(reg_q1050 AND symb_decoder(16#b9#)) OR
 					(reg_q1050 AND symb_decoder(16#9e#)) OR
 					(reg_q1050 AND symb_decoder(16#e6#)) OR
 					(reg_q1050 AND symb_decoder(16#44#)) OR
 					(reg_q1050 AND symb_decoder(16#d8#)) OR
 					(reg_q1050 AND symb_decoder(16#fa#)) OR
 					(reg_q1050 AND symb_decoder(16#07#)) OR
 					(reg_q1050 AND symb_decoder(16#89#)) OR
 					(reg_q1050 AND symb_decoder(16#00#)) OR
 					(reg_q1050 AND symb_decoder(16#65#)) OR
 					(reg_q1050 AND symb_decoder(16#9c#)) OR
 					(reg_q1050 AND symb_decoder(16#34#)) OR
 					(reg_q1050 AND symb_decoder(16#2d#)) OR
 					(reg_q1050 AND symb_decoder(16#7c#)) OR
 					(reg_q1050 AND symb_decoder(16#5c#)) OR
 					(reg_q1050 AND symb_decoder(16#6c#)) OR
 					(reg_q1050 AND symb_decoder(16#95#)) OR
 					(reg_q1050 AND symb_decoder(16#6e#)) OR
 					(reg_q1050 AND symb_decoder(16#91#)) OR
 					(reg_q1050 AND symb_decoder(16#f0#)) OR
 					(reg_q1050 AND symb_decoder(16#64#)) OR
 					(reg_q1050 AND symb_decoder(16#b8#)) OR
 					(reg_q1050 AND symb_decoder(16#56#)) OR
 					(reg_q1050 AND symb_decoder(16#6d#)) OR
 					(reg_q1050 AND symb_decoder(16#eb#)) OR
 					(reg_q1050 AND symb_decoder(16#62#)) OR
 					(reg_q1050 AND symb_decoder(16#59#)) OR
 					(reg_q1050 AND symb_decoder(16#9a#));
reg_q1050_init <= '0' ;
	p_reg_q1050: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1050 <= reg_q1050_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1050 <= reg_q1050_init;
        else
          reg_q1050 <= reg_q1050_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q780_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q779 AND symb_decoder(16#0d#)) OR
 					(reg_q779 AND symb_decoder(16#0a#));
reg_q780_init <= '0' ;
	p_reg_q780: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q780 <= reg_q780_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q780 <= reg_q780_init;
        else
          reg_q780 <= reg_q780_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2156_in <= (reg_q2154 AND symb_decoder(16#61#)) OR
 					(reg_q2154 AND symb_decoder(16#41#));
reg_q2156_init <= '0' ;
	p_reg_q2156: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2156 <= reg_q2156_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2156 <= reg_q2156_init;
        else
          reg_q2156 <= reg_q2156_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2158_in <= (reg_q2156 AND symb_decoder(16#54#)) OR
 					(reg_q2156 AND symb_decoder(16#74#));
reg_q2158_init <= '0' ;
	p_reg_q2158: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2158 <= reg_q2158_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2158 <= reg_q2158_init;
        else
          reg_q2158 <= reg_q2158_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1521_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1521 AND symb_decoder(16#35#)) OR
 					(reg_q1521 AND symb_decoder(16#4b#)) OR
 					(reg_q1521 AND symb_decoder(16#41#)) OR
 					(reg_q1521 AND symb_decoder(16#3a#)) OR
 					(reg_q1521 AND symb_decoder(16#0e#)) OR
 					(reg_q1521 AND symb_decoder(16#df#)) OR
 					(reg_q1521 AND symb_decoder(16#dd#)) OR
 					(reg_q1521 AND symb_decoder(16#a5#)) OR
 					(reg_q1521 AND symb_decoder(16#9a#)) OR
 					(reg_q1521 AND symb_decoder(16#59#)) OR
 					(reg_q1521 AND symb_decoder(16#0f#)) OR
 					(reg_q1521 AND symb_decoder(16#62#)) OR
 					(reg_q1521 AND symb_decoder(16#d5#)) OR
 					(reg_q1521 AND symb_decoder(16#50#)) OR
 					(reg_q1521 AND symb_decoder(16#56#)) OR
 					(reg_q1521 AND symb_decoder(16#24#)) OR
 					(reg_q1521 AND symb_decoder(16#84#)) OR
 					(reg_q1521 AND symb_decoder(16#8c#)) OR
 					(reg_q1521 AND symb_decoder(16#09#)) OR
 					(reg_q1521 AND symb_decoder(16#4e#)) OR
 					(reg_q1521 AND symb_decoder(16#b7#)) OR
 					(reg_q1521 AND symb_decoder(16#a0#)) OR
 					(reg_q1521 AND symb_decoder(16#2d#)) OR
 					(reg_q1521 AND symb_decoder(16#ce#)) OR
 					(reg_q1521 AND symb_decoder(16#7d#)) OR
 					(reg_q1521 AND symb_decoder(16#c1#)) OR
 					(reg_q1521 AND symb_decoder(16#63#)) OR
 					(reg_q1521 AND symb_decoder(16#65#)) OR
 					(reg_q1521 AND symb_decoder(16#67#)) OR
 					(reg_q1521 AND symb_decoder(16#29#)) OR
 					(reg_q1521 AND symb_decoder(16#11#)) OR
 					(reg_q1521 AND symb_decoder(16#81#)) OR
 					(reg_q1521 AND symb_decoder(16#07#)) OR
 					(reg_q1521 AND symb_decoder(16#91#)) OR
 					(reg_q1521 AND symb_decoder(16#68#)) OR
 					(reg_q1521 AND symb_decoder(16#1e#)) OR
 					(reg_q1521 AND symb_decoder(16#fc#)) OR
 					(reg_q1521 AND symb_decoder(16#1b#)) OR
 					(reg_q1521 AND symb_decoder(16#c0#)) OR
 					(reg_q1521 AND symb_decoder(16#c8#)) OR
 					(reg_q1521 AND symb_decoder(16#96#)) OR
 					(reg_q1521 AND symb_decoder(16#8f#)) OR
 					(reg_q1521 AND symb_decoder(16#6a#)) OR
 					(reg_q1521 AND symb_decoder(16#2b#)) OR
 					(reg_q1521 AND symb_decoder(16#cb#)) OR
 					(reg_q1521 AND symb_decoder(16#6e#)) OR
 					(reg_q1521 AND symb_decoder(16#b1#)) OR
 					(reg_q1521 AND symb_decoder(16#14#)) OR
 					(reg_q1521 AND symb_decoder(16#f8#)) OR
 					(reg_q1521 AND symb_decoder(16#5e#)) OR
 					(reg_q1521 AND symb_decoder(16#10#)) OR
 					(reg_q1521 AND symb_decoder(16#a6#)) OR
 					(reg_q1521 AND symb_decoder(16#37#)) OR
 					(reg_q1521 AND symb_decoder(16#f4#)) OR
 					(reg_q1521 AND symb_decoder(16#1a#)) OR
 					(reg_q1521 AND symb_decoder(16#f1#)) OR
 					(reg_q1521 AND symb_decoder(16#be#)) OR
 					(reg_q1521 AND symb_decoder(16#f3#)) OR
 					(reg_q1521 AND symb_decoder(16#46#)) OR
 					(reg_q1521 AND symb_decoder(16#38#)) OR
 					(reg_q1521 AND symb_decoder(16#06#)) OR
 					(reg_q1521 AND symb_decoder(16#39#)) OR
 					(reg_q1521 AND symb_decoder(16#0d#)) OR
 					(reg_q1521 AND symb_decoder(16#40#)) OR
 					(reg_q1521 AND symb_decoder(16#b0#)) OR
 					(reg_q1521 AND symb_decoder(16#b6#)) OR
 					(reg_q1521 AND symb_decoder(16#0a#)) OR
 					(reg_q1521 AND symb_decoder(16#ec#)) OR
 					(reg_q1521 AND symb_decoder(16#53#)) OR
 					(reg_q1521 AND symb_decoder(16#20#)) OR
 					(reg_q1521 AND symb_decoder(16#86#)) OR
 					(reg_q1521 AND symb_decoder(16#98#)) OR
 					(reg_q1521 AND symb_decoder(16#ab#)) OR
 					(reg_q1521 AND symb_decoder(16#a9#)) OR
 					(reg_q1521 AND symb_decoder(16#75#)) OR
 					(reg_q1521 AND symb_decoder(16#e2#)) OR
 					(reg_q1521 AND symb_decoder(16#47#)) OR
 					(reg_q1521 AND symb_decoder(16#e4#)) OR
 					(reg_q1521 AND symb_decoder(16#4d#)) OR
 					(reg_q1521 AND symb_decoder(16#9f#)) OR
 					(reg_q1521 AND symb_decoder(16#12#)) OR
 					(reg_q1521 AND symb_decoder(16#49#)) OR
 					(reg_q1521 AND symb_decoder(16#c5#)) OR
 					(reg_q1521 AND symb_decoder(16#73#)) OR
 					(reg_q1521 AND symb_decoder(16#2c#)) OR
 					(reg_q1521 AND symb_decoder(16#42#)) OR
 					(reg_q1521 AND symb_decoder(16#cf#)) OR
 					(reg_q1521 AND symb_decoder(16#c6#)) OR
 					(reg_q1521 AND symb_decoder(16#93#)) OR
 					(reg_q1521 AND symb_decoder(16#33#)) OR
 					(reg_q1521 AND symb_decoder(16#74#)) OR
 					(reg_q1521 AND symb_decoder(16#f9#)) OR
 					(reg_q1521 AND symb_decoder(16#64#)) OR
 					(reg_q1521 AND symb_decoder(16#92#)) OR
 					(reg_q1521 AND symb_decoder(16#18#)) OR
 					(reg_q1521 AND symb_decoder(16#97#)) OR
 					(reg_q1521 AND symb_decoder(16#6d#)) OR
 					(reg_q1521 AND symb_decoder(16#17#)) OR
 					(reg_q1521 AND symb_decoder(16#2a#)) OR
 					(reg_q1521 AND symb_decoder(16#ee#)) OR
 					(reg_q1521 AND symb_decoder(16#de#)) OR
 					(reg_q1521 AND symb_decoder(16#a3#)) OR
 					(reg_q1521 AND symb_decoder(16#5b#)) OR
 					(reg_q1521 AND symb_decoder(16#b3#)) OR
 					(reg_q1521 AND symb_decoder(16#89#)) OR
 					(reg_q1521 AND symb_decoder(16#4a#)) OR
 					(reg_q1521 AND symb_decoder(16#61#)) OR
 					(reg_q1521 AND symb_decoder(16#36#)) OR
 					(reg_q1521 AND symb_decoder(16#7e#)) OR
 					(reg_q1521 AND symb_decoder(16#28#)) OR
 					(reg_q1521 AND symb_decoder(16#72#)) OR
 					(reg_q1521 AND symb_decoder(16#c4#)) OR
 					(reg_q1521 AND symb_decoder(16#9c#)) OR
 					(reg_q1521 AND symb_decoder(16#77#)) OR
 					(reg_q1521 AND symb_decoder(16#44#)) OR
 					(reg_q1521 AND symb_decoder(16#cd#)) OR
 					(reg_q1521 AND symb_decoder(16#f5#)) OR
 					(reg_q1521 AND symb_decoder(16#2f#)) OR
 					(reg_q1521 AND symb_decoder(16#c2#)) OR
 					(reg_q1521 AND symb_decoder(16#31#)) OR
 					(reg_q1521 AND symb_decoder(16#d7#)) OR
 					(reg_q1521 AND symb_decoder(16#db#)) OR
 					(reg_q1521 AND symb_decoder(16#dc#)) OR
 					(reg_q1521 AND symb_decoder(16#04#)) OR
 					(reg_q1521 AND symb_decoder(16#51#)) OR
 					(reg_q1521 AND symb_decoder(16#7b#)) OR
 					(reg_q1521 AND symb_decoder(16#e0#)) OR
 					(reg_q1521 AND symb_decoder(16#76#)) OR
 					(reg_q1521 AND symb_decoder(16#1f#)) OR
 					(reg_q1521 AND symb_decoder(16#88#)) OR
 					(reg_q1521 AND symb_decoder(16#bf#)) OR
 					(reg_q1521 AND symb_decoder(16#95#)) OR
 					(reg_q1521 AND symb_decoder(16#ed#)) OR
 					(reg_q1521 AND symb_decoder(16#ea#)) OR
 					(reg_q1521 AND symb_decoder(16#0b#)) OR
 					(reg_q1521 AND symb_decoder(16#22#)) OR
 					(reg_q1521 AND symb_decoder(16#8e#)) OR
 					(reg_q1521 AND symb_decoder(16#0c#)) OR
 					(reg_q1521 AND symb_decoder(16#66#)) OR
 					(reg_q1521 AND symb_decoder(16#6f#)) OR
 					(reg_q1521 AND symb_decoder(16#c7#)) OR
 					(reg_q1521 AND symb_decoder(16#e8#)) OR
 					(reg_q1521 AND symb_decoder(16#6b#)) OR
 					(reg_q1521 AND symb_decoder(16#fe#)) OR
 					(reg_q1521 AND symb_decoder(16#bd#)) OR
 					(reg_q1521 AND symb_decoder(16#a7#)) OR
 					(reg_q1521 AND symb_decoder(16#f2#)) OR
 					(reg_q1521 AND symb_decoder(16#d6#)) OR
 					(reg_q1521 AND symb_decoder(16#52#)) OR
 					(reg_q1521 AND symb_decoder(16#4c#)) OR
 					(reg_q1521 AND symb_decoder(16#b5#)) OR
 					(reg_q1521 AND symb_decoder(16#8a#)) OR
 					(reg_q1521 AND symb_decoder(16#54#)) OR
 					(reg_q1521 AND symb_decoder(16#30#)) OR
 					(reg_q1521 AND symb_decoder(16#d3#)) OR
 					(reg_q1521 AND symb_decoder(16#8b#)) OR
 					(reg_q1521 AND symb_decoder(16#3c#)) OR
 					(reg_q1521 AND symb_decoder(16#d2#)) OR
 					(reg_q1521 AND symb_decoder(16#cc#)) OR
 					(reg_q1521 AND symb_decoder(16#78#)) OR
 					(reg_q1521 AND symb_decoder(16#2e#)) OR
 					(reg_q1521 AND symb_decoder(16#5d#)) OR
 					(reg_q1521 AND symb_decoder(16#aa#)) OR
 					(reg_q1521 AND symb_decoder(16#3f#)) OR
 					(reg_q1521 AND symb_decoder(16#34#)) OR
 					(reg_q1521 AND symb_decoder(16#83#)) OR
 					(reg_q1521 AND symb_decoder(16#ac#)) OR
 					(reg_q1521 AND symb_decoder(16#9b#)) OR
 					(reg_q1521 AND symb_decoder(16#af#)) OR
 					(reg_q1521 AND symb_decoder(16#a8#)) OR
 					(reg_q1521 AND symb_decoder(16#b2#)) OR
 					(reg_q1521 AND symb_decoder(16#9d#)) OR
 					(reg_q1521 AND symb_decoder(16#a2#)) OR
 					(reg_q1521 AND symb_decoder(16#d9#)) OR
 					(reg_q1521 AND symb_decoder(16#f6#)) OR
 					(reg_q1521 AND symb_decoder(16#e6#)) OR
 					(reg_q1521 AND symb_decoder(16#3e#)) OR
 					(reg_q1521 AND symb_decoder(16#45#)) OR
 					(reg_q1521 AND symb_decoder(16#1d#)) OR
 					(reg_q1521 AND symb_decoder(16#90#)) OR
 					(reg_q1521 AND symb_decoder(16#87#)) OR
 					(reg_q1521 AND symb_decoder(16#7a#)) OR
 					(reg_q1521 AND symb_decoder(16#9e#)) OR
 					(reg_q1521 AND symb_decoder(16#55#)) OR
 					(reg_q1521 AND symb_decoder(16#00#)) OR
 					(reg_q1521 AND symb_decoder(16#fd#)) OR
 					(reg_q1521 AND symb_decoder(16#13#)) OR
 					(reg_q1521 AND symb_decoder(16#16#)) OR
 					(reg_q1521 AND symb_decoder(16#69#)) OR
 					(reg_q1521 AND symb_decoder(16#02#)) OR
 					(reg_q1521 AND symb_decoder(16#ca#)) OR
 					(reg_q1521 AND symb_decoder(16#58#)) OR
 					(reg_q1521 AND symb_decoder(16#80#)) OR
 					(reg_q1521 AND symb_decoder(16#fa#)) OR
 					(reg_q1521 AND symb_decoder(16#ad#)) OR
 					(reg_q1521 AND symb_decoder(16#3b#)) OR
 					(reg_q1521 AND symb_decoder(16#99#)) OR
 					(reg_q1521 AND symb_decoder(16#a4#)) OR
 					(reg_q1521 AND symb_decoder(16#05#)) OR
 					(reg_q1521 AND symb_decoder(16#60#)) OR
 					(reg_q1521 AND symb_decoder(16#e7#)) OR
 					(reg_q1521 AND symb_decoder(16#5a#)) OR
 					(reg_q1521 AND symb_decoder(16#01#)) OR
 					(reg_q1521 AND symb_decoder(16#d1#)) OR
 					(reg_q1521 AND symb_decoder(16#ae#)) OR
 					(reg_q1521 AND symb_decoder(16#ff#)) OR
 					(reg_q1521 AND symb_decoder(16#32#)) OR
 					(reg_q1521 AND symb_decoder(16#e5#)) OR
 					(reg_q1521 AND symb_decoder(16#5f#)) OR
 					(reg_q1521 AND symb_decoder(16#27#)) OR
 					(reg_q1521 AND symb_decoder(16#5c#)) OR
 					(reg_q1521 AND symb_decoder(16#43#)) OR
 					(reg_q1521 AND symb_decoder(16#b8#)) OR
 					(reg_q1521 AND symb_decoder(16#08#)) OR
 					(reg_q1521 AND symb_decoder(16#03#)) OR
 					(reg_q1521 AND symb_decoder(16#d4#)) OR
 					(reg_q1521 AND symb_decoder(16#da#)) OR
 					(reg_q1521 AND symb_decoder(16#48#)) OR
 					(reg_q1521 AND symb_decoder(16#94#)) OR
 					(reg_q1521 AND symb_decoder(16#26#)) OR
 					(reg_q1521 AND symb_decoder(16#b9#)) OR
 					(reg_q1521 AND symb_decoder(16#bc#)) OR
 					(reg_q1521 AND symb_decoder(16#d0#)) OR
 					(reg_q1521 AND symb_decoder(16#71#)) OR
 					(reg_q1521 AND symb_decoder(16#a1#)) OR
 					(reg_q1521 AND symb_decoder(16#c3#)) OR
 					(reg_q1521 AND symb_decoder(16#fb#)) OR
 					(reg_q1521 AND symb_decoder(16#82#)) OR
 					(reg_q1521 AND symb_decoder(16#f7#)) OR
 					(reg_q1521 AND symb_decoder(16#7c#)) OR
 					(reg_q1521 AND symb_decoder(16#57#)) OR
 					(reg_q1521 AND symb_decoder(16#e9#)) OR
 					(reg_q1521 AND symb_decoder(16#8d#)) OR
 					(reg_q1521 AND symb_decoder(16#19#)) OR
 					(reg_q1521 AND symb_decoder(16#bb#)) OR
 					(reg_q1521 AND symb_decoder(16#70#)) OR
 					(reg_q1521 AND symb_decoder(16#85#)) OR
 					(reg_q1521 AND symb_decoder(16#e1#)) OR
 					(reg_q1521 AND symb_decoder(16#1c#)) OR
 					(reg_q1521 AND symb_decoder(16#e3#)) OR
 					(reg_q1521 AND symb_decoder(16#21#)) OR
 					(reg_q1521 AND symb_decoder(16#eb#)) OR
 					(reg_q1521 AND symb_decoder(16#7f#)) OR
 					(reg_q1521 AND symb_decoder(16#23#)) OR
 					(reg_q1521 AND symb_decoder(16#3d#)) OR
 					(reg_q1521 AND symb_decoder(16#79#)) OR
 					(reg_q1521 AND symb_decoder(16#ef#)) OR
 					(reg_q1521 AND symb_decoder(16#c9#)) OR
 					(reg_q1521 AND symb_decoder(16#25#)) OR
 					(reg_q1521 AND symb_decoder(16#d8#)) OR
 					(reg_q1521 AND symb_decoder(16#b4#)) OR
 					(reg_q1521 AND symb_decoder(16#4f#)) OR
 					(reg_q1521 AND symb_decoder(16#15#)) OR
 					(reg_q1521 AND symb_decoder(16#f0#)) OR
 					(reg_q1521 AND symb_decoder(16#6c#)) OR
 					(reg_q1521 AND symb_decoder(16#ba#));
reg_q1521_init <= '0' ;
	p_reg_q1521: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1521 <= reg_q1521_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1521 <= reg_q1521_init;
        else
          reg_q1521 <= reg_q1521_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1377_in <= (reg_q1375 AND symb_decoder(16#69#)) OR
 					(reg_q1375 AND symb_decoder(16#49#));
reg_q1377_init <= '0' ;
	p_reg_q1377: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1377 <= reg_q1377_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1377 <= reg_q1377_init;
        else
          reg_q1377 <= reg_q1377_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1379_in <= (reg_q1377 AND symb_decoder(16#4c#)) OR
 					(reg_q1377 AND symb_decoder(16#6c#));
reg_q1379_init <= '0' ;
	p_reg_q1379: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1379 <= reg_q1379_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1379 <= reg_q1379_init;
        else
          reg_q1379 <= reg_q1379_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q688_in <= (reg_q688 AND symb_decoder(16#37#)) OR
 					(reg_q688 AND symb_decoder(16#36#)) OR
 					(reg_q688 AND symb_decoder(16#31#)) OR
 					(reg_q688 AND symb_decoder(16#33#)) OR
 					(reg_q688 AND symb_decoder(16#39#)) OR
 					(reg_q688 AND symb_decoder(16#30#)) OR
 					(reg_q688 AND symb_decoder(16#35#)) OR
 					(reg_q688 AND symb_decoder(16#38#)) OR
 					(reg_q688 AND symb_decoder(16#32#)) OR
 					(reg_q688 AND symb_decoder(16#34#)) OR
 					(reg_q686 AND symb_decoder(16#38#)) OR
 					(reg_q686 AND symb_decoder(16#30#)) OR
 					(reg_q686 AND symb_decoder(16#35#)) OR
 					(reg_q686 AND symb_decoder(16#32#)) OR
 					(reg_q686 AND symb_decoder(16#34#)) OR
 					(reg_q686 AND symb_decoder(16#31#)) OR
 					(reg_q686 AND symb_decoder(16#37#)) OR
 					(reg_q686 AND symb_decoder(16#33#)) OR
 					(reg_q686 AND symb_decoder(16#39#)) OR
 					(reg_q686 AND symb_decoder(16#36#));
reg_q688_init <= '0' ;
	p_reg_q688: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q688 <= reg_q688_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q688 <= reg_q688_init;
        else
          reg_q688 <= reg_q688_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q690_in <= (reg_q688 AND symb_decoder(16#2e#));
reg_q690_init <= '0' ;
	p_reg_q690: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q690 <= reg_q690_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q690 <= reg_q690_init;
        else
          reg_q690 <= reg_q690_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q644_in <= (reg_q642 AND symb_decoder(16#45#)) OR
 					(reg_q642 AND symb_decoder(16#65#));
reg_q644_init <= '0' ;
	p_reg_q644: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q644 <= reg_q644_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q644 <= reg_q644_init;
        else
          reg_q644 <= reg_q644_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q646_in <= (reg_q644 AND symb_decoder(16#25#));
reg_q646_init <= '0' ;
	p_reg_q646: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q646 <= reg_q646_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q646 <= reg_q646_init;
        else
          reg_q646 <= reg_q646_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1955_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1955 AND symb_decoder(16#54#)) OR
 					(reg_q1955 AND symb_decoder(16#b7#)) OR
 					(reg_q1955 AND symb_decoder(16#20#)) OR
 					(reg_q1955 AND symb_decoder(16#c3#)) OR
 					(reg_q1955 AND symb_decoder(16#c6#)) OR
 					(reg_q1955 AND symb_decoder(16#10#)) OR
 					(reg_q1955 AND symb_decoder(16#ed#)) OR
 					(reg_q1955 AND symb_decoder(16#61#)) OR
 					(reg_q1955 AND symb_decoder(16#3b#)) OR
 					(reg_q1955 AND symb_decoder(16#43#)) OR
 					(reg_q1955 AND symb_decoder(16#0f#)) OR
 					(reg_q1955 AND symb_decoder(16#6b#)) OR
 					(reg_q1955 AND symb_decoder(16#b3#)) OR
 					(reg_q1955 AND symb_decoder(16#9d#)) OR
 					(reg_q1955 AND symb_decoder(16#a6#)) OR
 					(reg_q1955 AND symb_decoder(16#79#)) OR
 					(reg_q1955 AND symb_decoder(16#65#)) OR
 					(reg_q1955 AND symb_decoder(16#9e#)) OR
 					(reg_q1955 AND symb_decoder(16#d0#)) OR
 					(reg_q1955 AND symb_decoder(16#d5#)) OR
 					(reg_q1955 AND symb_decoder(16#c7#)) OR
 					(reg_q1955 AND symb_decoder(16#63#)) OR
 					(reg_q1955 AND symb_decoder(16#56#)) OR
 					(reg_q1955 AND symb_decoder(16#27#)) OR
 					(reg_q1955 AND symb_decoder(16#97#)) OR
 					(reg_q1955 AND symb_decoder(16#ab#)) OR
 					(reg_q1955 AND symb_decoder(16#ff#)) OR
 					(reg_q1955 AND symb_decoder(16#34#)) OR
 					(reg_q1955 AND symb_decoder(16#4f#)) OR
 					(reg_q1955 AND symb_decoder(16#19#)) OR
 					(reg_q1955 AND symb_decoder(16#5f#)) OR
 					(reg_q1955 AND symb_decoder(16#3e#)) OR
 					(reg_q1955 AND symb_decoder(16#7c#)) OR
 					(reg_q1955 AND symb_decoder(16#82#)) OR
 					(reg_q1955 AND symb_decoder(16#cc#)) OR
 					(reg_q1955 AND symb_decoder(16#dc#)) OR
 					(reg_q1955 AND symb_decoder(16#59#)) OR
 					(reg_q1955 AND symb_decoder(16#f8#)) OR
 					(reg_q1955 AND symb_decoder(16#72#)) OR
 					(reg_q1955 AND symb_decoder(16#cb#)) OR
 					(reg_q1955 AND symb_decoder(16#0a#)) OR
 					(reg_q1955 AND symb_decoder(16#38#)) OR
 					(reg_q1955 AND symb_decoder(16#b9#)) OR
 					(reg_q1955 AND symb_decoder(16#69#)) OR
 					(reg_q1955 AND symb_decoder(16#52#)) OR
 					(reg_q1955 AND symb_decoder(16#c4#)) OR
 					(reg_q1955 AND symb_decoder(16#78#)) OR
 					(reg_q1955 AND symb_decoder(16#6f#)) OR
 					(reg_q1955 AND symb_decoder(16#cd#)) OR
 					(reg_q1955 AND symb_decoder(16#ba#)) OR
 					(reg_q1955 AND symb_decoder(16#c8#)) OR
 					(reg_q1955 AND symb_decoder(16#f9#)) OR
 					(reg_q1955 AND symb_decoder(16#be#)) OR
 					(reg_q1955 AND symb_decoder(16#2a#)) OR
 					(reg_q1955 AND symb_decoder(16#8e#)) OR
 					(reg_q1955 AND symb_decoder(16#b1#)) OR
 					(reg_q1955 AND symb_decoder(16#aa#)) OR
 					(reg_q1955 AND symb_decoder(16#81#)) OR
 					(reg_q1955 AND symb_decoder(16#51#)) OR
 					(reg_q1955 AND symb_decoder(16#4b#)) OR
 					(reg_q1955 AND symb_decoder(16#ae#)) OR
 					(reg_q1955 AND symb_decoder(16#3d#)) OR
 					(reg_q1955 AND symb_decoder(16#8c#)) OR
 					(reg_q1955 AND symb_decoder(16#87#)) OR
 					(reg_q1955 AND symb_decoder(16#95#)) OR
 					(reg_q1955 AND symb_decoder(16#c1#)) OR
 					(reg_q1955 AND symb_decoder(16#d3#)) OR
 					(reg_q1955 AND symb_decoder(16#29#)) OR
 					(reg_q1955 AND symb_decoder(16#9b#)) OR
 					(reg_q1955 AND symb_decoder(16#33#)) OR
 					(reg_q1955 AND symb_decoder(16#fc#)) OR
 					(reg_q1955 AND symb_decoder(16#f0#)) OR
 					(reg_q1955 AND symb_decoder(16#7b#)) OR
 					(reg_q1955 AND symb_decoder(16#6c#)) OR
 					(reg_q1955 AND symb_decoder(16#37#)) OR
 					(reg_q1955 AND symb_decoder(16#2f#)) OR
 					(reg_q1955 AND symb_decoder(16#e6#)) OR
 					(reg_q1955 AND symb_decoder(16#86#)) OR
 					(reg_q1955 AND symb_decoder(16#1e#)) OR
 					(reg_q1955 AND symb_decoder(16#e2#)) OR
 					(reg_q1955 AND symb_decoder(16#f7#)) OR
 					(reg_q1955 AND symb_decoder(16#fd#)) OR
 					(reg_q1955 AND symb_decoder(16#04#)) OR
 					(reg_q1955 AND symb_decoder(16#dd#)) OR
 					(reg_q1955 AND symb_decoder(16#e0#)) OR
 					(reg_q1955 AND symb_decoder(16#12#)) OR
 					(reg_q1955 AND symb_decoder(16#7d#)) OR
 					(reg_q1955 AND symb_decoder(16#ec#)) OR
 					(reg_q1955 AND symb_decoder(16#03#)) OR
 					(reg_q1955 AND symb_decoder(16#f1#)) OR
 					(reg_q1955 AND symb_decoder(16#f5#)) OR
 					(reg_q1955 AND symb_decoder(16#b5#)) OR
 					(reg_q1955 AND symb_decoder(16#a0#)) OR
 					(reg_q1955 AND symb_decoder(16#73#)) OR
 					(reg_q1955 AND symb_decoder(16#5c#)) OR
 					(reg_q1955 AND symb_decoder(16#90#)) OR
 					(reg_q1955 AND symb_decoder(16#42#)) OR
 					(reg_q1955 AND symb_decoder(16#b6#)) OR
 					(reg_q1955 AND symb_decoder(16#05#)) OR
 					(reg_q1955 AND symb_decoder(16#93#)) OR
 					(reg_q1955 AND symb_decoder(16#83#)) OR
 					(reg_q1955 AND symb_decoder(16#e3#)) OR
 					(reg_q1955 AND symb_decoder(16#f2#)) OR
 					(reg_q1955 AND symb_decoder(16#57#)) OR
 					(reg_q1955 AND symb_decoder(16#4a#)) OR
 					(reg_q1955 AND symb_decoder(16#01#)) OR
 					(reg_q1955 AND symb_decoder(16#23#)) OR
 					(reg_q1955 AND symb_decoder(16#6d#)) OR
 					(reg_q1955 AND symb_decoder(16#2d#)) OR
 					(reg_q1955 AND symb_decoder(16#94#)) OR
 					(reg_q1955 AND symb_decoder(16#16#)) OR
 					(reg_q1955 AND symb_decoder(16#2b#)) OR
 					(reg_q1955 AND symb_decoder(16#74#)) OR
 					(reg_q1955 AND symb_decoder(16#49#)) OR
 					(reg_q1955 AND symb_decoder(16#66#)) OR
 					(reg_q1955 AND symb_decoder(16#5a#)) OR
 					(reg_q1955 AND symb_decoder(16#5e#)) OR
 					(reg_q1955 AND symb_decoder(16#8b#)) OR
 					(reg_q1955 AND symb_decoder(16#00#)) OR
 					(reg_q1955 AND symb_decoder(16#7f#)) OR
 					(reg_q1955 AND symb_decoder(16#e4#)) OR
 					(reg_q1955 AND symb_decoder(16#ac#)) OR
 					(reg_q1955 AND symb_decoder(16#3a#)) OR
 					(reg_q1955 AND symb_decoder(16#91#)) OR
 					(reg_q1955 AND symb_decoder(16#df#)) OR
 					(reg_q1955 AND symb_decoder(16#3c#)) OR
 					(reg_q1955 AND symb_decoder(16#8f#)) OR
 					(reg_q1955 AND symb_decoder(16#8a#)) OR
 					(reg_q1955 AND symb_decoder(16#50#)) OR
 					(reg_q1955 AND symb_decoder(16#e7#)) OR
 					(reg_q1955 AND symb_decoder(16#48#)) OR
 					(reg_q1955 AND symb_decoder(16#47#)) OR
 					(reg_q1955 AND symb_decoder(16#eb#)) OR
 					(reg_q1955 AND symb_decoder(16#13#)) OR
 					(reg_q1955 AND symb_decoder(16#a7#)) OR
 					(reg_q1955 AND symb_decoder(16#31#)) OR
 					(reg_q1955 AND symb_decoder(16#4d#)) OR
 					(reg_q1955 AND symb_decoder(16#0b#)) OR
 					(reg_q1955 AND symb_decoder(16#0e#)) OR
 					(reg_q1955 AND symb_decoder(16#71#)) OR
 					(reg_q1955 AND symb_decoder(16#06#)) OR
 					(reg_q1955 AND symb_decoder(16#17#)) OR
 					(reg_q1955 AND symb_decoder(16#7e#)) OR
 					(reg_q1955 AND symb_decoder(16#1a#)) OR
 					(reg_q1955 AND symb_decoder(16#15#)) OR
 					(reg_q1955 AND symb_decoder(16#41#)) OR
 					(reg_q1955 AND symb_decoder(16#30#)) OR
 					(reg_q1955 AND symb_decoder(16#bb#)) OR
 					(reg_q1955 AND symb_decoder(16#76#)) OR
 					(reg_q1955 AND symb_decoder(16#c9#)) OR
 					(reg_q1955 AND symb_decoder(16#58#)) OR
 					(reg_q1955 AND symb_decoder(16#68#)) OR
 					(reg_q1955 AND symb_decoder(16#f6#)) OR
 					(reg_q1955 AND symb_decoder(16#fe#)) OR
 					(reg_q1955 AND symb_decoder(16#cf#)) OR
 					(reg_q1955 AND symb_decoder(16#53#)) OR
 					(reg_q1955 AND symb_decoder(16#a4#)) OR
 					(reg_q1955 AND symb_decoder(16#b8#)) OR
 					(reg_q1955 AND symb_decoder(16#f3#)) OR
 					(reg_q1955 AND symb_decoder(16#a1#)) OR
 					(reg_q1955 AND symb_decoder(16#d4#)) OR
 					(reg_q1955 AND symb_decoder(16#11#)) OR
 					(reg_q1955 AND symb_decoder(16#45#)) OR
 					(reg_q1955 AND symb_decoder(16#44#)) OR
 					(reg_q1955 AND symb_decoder(16#ef#)) OR
 					(reg_q1955 AND symb_decoder(16#25#)) OR
 					(reg_q1955 AND symb_decoder(16#4e#)) OR
 					(reg_q1955 AND symb_decoder(16#c2#)) OR
 					(reg_q1955 AND symb_decoder(16#d6#)) OR
 					(reg_q1955 AND symb_decoder(16#6e#)) OR
 					(reg_q1955 AND symb_decoder(16#18#)) OR
 					(reg_q1955 AND symb_decoder(16#6a#)) OR
 					(reg_q1955 AND symb_decoder(16#99#)) OR
 					(reg_q1955 AND symb_decoder(16#21#)) OR
 					(reg_q1955 AND symb_decoder(16#02#)) OR
 					(reg_q1955 AND symb_decoder(16#fa#)) OR
 					(reg_q1955 AND symb_decoder(16#0d#)) OR
 					(reg_q1955 AND symb_decoder(16#46#)) OR
 					(reg_q1955 AND symb_decoder(16#a9#)) OR
 					(reg_q1955 AND symb_decoder(16#64#)) OR
 					(reg_q1955 AND symb_decoder(16#b0#)) OR
 					(reg_q1955 AND symb_decoder(16#e5#)) OR
 					(reg_q1955 AND symb_decoder(16#c0#)) OR
 					(reg_q1955 AND symb_decoder(16#8d#)) OR
 					(reg_q1955 AND symb_decoder(16#1c#)) OR
 					(reg_q1955 AND symb_decoder(16#f4#)) OR
 					(reg_q1955 AND symb_decoder(16#2c#)) OR
 					(reg_q1955 AND symb_decoder(16#d8#)) OR
 					(reg_q1955 AND symb_decoder(16#1d#)) OR
 					(reg_q1955 AND symb_decoder(16#36#)) OR
 					(reg_q1955 AND symb_decoder(16#3f#)) OR
 					(reg_q1955 AND symb_decoder(16#60#)) OR
 					(reg_q1955 AND symb_decoder(16#ca#)) OR
 					(reg_q1955 AND symb_decoder(16#1f#)) OR
 					(reg_q1955 AND symb_decoder(16#92#)) OR
 					(reg_q1955 AND symb_decoder(16#bd#)) OR
 					(reg_q1955 AND symb_decoder(16#08#)) OR
 					(reg_q1955 AND symb_decoder(16#5d#)) OR
 					(reg_q1955 AND symb_decoder(16#fb#)) OR
 					(reg_q1955 AND symb_decoder(16#db#)) OR
 					(reg_q1955 AND symb_decoder(16#a3#)) OR
 					(reg_q1955 AND symb_decoder(16#d1#)) OR
 					(reg_q1955 AND symb_decoder(16#e8#)) OR
 					(reg_q1955 AND symb_decoder(16#88#)) OR
 					(reg_q1955 AND symb_decoder(16#85#)) OR
 					(reg_q1955 AND symb_decoder(16#b4#)) OR
 					(reg_q1955 AND symb_decoder(16#4c#)) OR
 					(reg_q1955 AND symb_decoder(16#2e#)) OR
 					(reg_q1955 AND symb_decoder(16#55#)) OR
 					(reg_q1955 AND symb_decoder(16#a8#)) OR
 					(reg_q1955 AND symb_decoder(16#a2#)) OR
 					(reg_q1955 AND symb_decoder(16#7a#)) OR
 					(reg_q1955 AND symb_decoder(16#0c#)) OR
 					(reg_q1955 AND symb_decoder(16#5b#)) OR
 					(reg_q1955 AND symb_decoder(16#14#)) OR
 					(reg_q1955 AND symb_decoder(16#de#)) OR
 					(reg_q1955 AND symb_decoder(16#9a#)) OR
 					(reg_q1955 AND symb_decoder(16#28#)) OR
 					(reg_q1955 AND symb_decoder(16#a5#)) OR
 					(reg_q1955 AND symb_decoder(16#d2#)) OR
 					(reg_q1955 AND symb_decoder(16#62#)) OR
 					(reg_q1955 AND symb_decoder(16#e9#)) OR
 					(reg_q1955 AND symb_decoder(16#35#)) OR
 					(reg_q1955 AND symb_decoder(16#9f#)) OR
 					(reg_q1955 AND symb_decoder(16#09#)) OR
 					(reg_q1955 AND symb_decoder(16#e1#)) OR
 					(reg_q1955 AND symb_decoder(16#ea#)) OR
 					(reg_q1955 AND symb_decoder(16#da#)) OR
 					(reg_q1955 AND symb_decoder(16#98#)) OR
 					(reg_q1955 AND symb_decoder(16#24#)) OR
 					(reg_q1955 AND symb_decoder(16#67#)) OR
 					(reg_q1955 AND symb_decoder(16#d9#)) OR
 					(reg_q1955 AND symb_decoder(16#32#)) OR
 					(reg_q1955 AND symb_decoder(16#bc#)) OR
 					(reg_q1955 AND symb_decoder(16#84#)) OR
 					(reg_q1955 AND symb_decoder(16#70#)) OR
 					(reg_q1955 AND symb_decoder(16#39#)) OR
 					(reg_q1955 AND symb_decoder(16#d7#)) OR
 					(reg_q1955 AND symb_decoder(16#89#)) OR
 					(reg_q1955 AND symb_decoder(16#40#)) OR
 					(reg_q1955 AND symb_decoder(16#75#)) OR
 					(reg_q1955 AND symb_decoder(16#77#)) OR
 					(reg_q1955 AND symb_decoder(16#1b#)) OR
 					(reg_q1955 AND symb_decoder(16#c5#)) OR
 					(reg_q1955 AND symb_decoder(16#ce#)) OR
 					(reg_q1955 AND symb_decoder(16#22#)) OR
 					(reg_q1955 AND symb_decoder(16#80#)) OR
 					(reg_q1955 AND symb_decoder(16#af#)) OR
 					(reg_q1955 AND symb_decoder(16#26#)) OR
 					(reg_q1955 AND symb_decoder(16#bf#)) OR
 					(reg_q1955 AND symb_decoder(16#ad#)) OR
 					(reg_q1955 AND symb_decoder(16#b2#)) OR
 					(reg_q1955 AND symb_decoder(16#07#)) OR
 					(reg_q1955 AND symb_decoder(16#96#)) OR
 					(reg_q1955 AND symb_decoder(16#9c#)) OR
 					(reg_q1955 AND symb_decoder(16#ee#));
reg_q1955_init <= '0' ;
	p_reg_q1955: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1955 <= reg_q1955_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1955 <= reg_q1955_init;
        else
          reg_q1955 <= reg_q1955_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1848_in <= (reg_q1848 AND symb_decoder(16#20#)) OR
 					(reg_q1848 AND symb_decoder(16#0c#)) OR
 					(reg_q1848 AND symb_decoder(16#09#)) OR
 					(reg_q1848 AND symb_decoder(16#0a#)) OR
 					(reg_q1848 AND symb_decoder(16#0d#)) OR
 					(reg_q1846 AND symb_decoder(16#0c#)) OR
 					(reg_q1846 AND symb_decoder(16#0a#)) OR
 					(reg_q1846 AND symb_decoder(16#09#)) OR
 					(reg_q1846 AND symb_decoder(16#20#)) OR
 					(reg_q1846 AND symb_decoder(16#0d#));
reg_q1848_init <= '0' ;
	p_reg_q1848: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1848 <= reg_q1848_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1848 <= reg_q1848_init;
        else
          reg_q1848 <= reg_q1848_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q52_in <= (reg_q50 AND symb_decoder(16#30#));
reg_q52_init <= '0' ;
	p_reg_q52: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q52 <= reg_q52_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q52 <= reg_q52_init;
        else
          reg_q52 <= reg_q52_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q54_in <= (reg_q52 AND symb_decoder(16#4f#)) OR
 					(reg_q52 AND symb_decoder(16#6f#));
reg_q54_init <= '0' ;
	p_reg_q54: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q54 <= reg_q54_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q54 <= reg_q54_init;
        else
          reg_q54 <= reg_q54_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q630_in <= (reg_q628 AND symb_decoder(16#52#)) OR
 					(reg_q628 AND symb_decoder(16#72#));
reg_q630_init <= '0' ;
	p_reg_q630: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q630 <= reg_q630_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q630 <= reg_q630_init;
        else
          reg_q630 <= reg_q630_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q632_in <= (reg_q630 AND symb_decoder(16#0a#)) OR
 					(reg_q630 AND symb_decoder(16#0c#)) OR
 					(reg_q630 AND symb_decoder(16#0d#)) OR
 					(reg_q630 AND symb_decoder(16#09#)) OR
 					(reg_q630 AND symb_decoder(16#20#)) OR
 					(reg_q632 AND symb_decoder(16#0d#)) OR
 					(reg_q632 AND symb_decoder(16#0a#)) OR
 					(reg_q632 AND symb_decoder(16#0c#)) OR
 					(reg_q632 AND symb_decoder(16#20#)) OR
 					(reg_q632 AND symb_decoder(16#09#));
reg_q632_init <= '0' ;
	p_reg_q632: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q632 <= reg_q632_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q632 <= reg_q632_init;
        else
          reg_q632 <= reg_q632_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q703_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q703 AND symb_decoder(16#a5#)) OR
 					(reg_q703 AND symb_decoder(16#40#)) OR
 					(reg_q703 AND symb_decoder(16#1f#)) OR
 					(reg_q703 AND symb_decoder(16#95#)) OR
 					(reg_q703 AND symb_decoder(16#5e#)) OR
 					(reg_q703 AND symb_decoder(16#4b#)) OR
 					(reg_q703 AND symb_decoder(16#8e#)) OR
 					(reg_q703 AND symb_decoder(16#0d#)) OR
 					(reg_q703 AND symb_decoder(16#46#)) OR
 					(reg_q703 AND symb_decoder(16#90#)) OR
 					(reg_q703 AND symb_decoder(16#ad#)) OR
 					(reg_q703 AND symb_decoder(16#e3#)) OR
 					(reg_q703 AND symb_decoder(16#df#)) OR
 					(reg_q703 AND symb_decoder(16#29#)) OR
 					(reg_q703 AND symb_decoder(16#8f#)) OR
 					(reg_q703 AND symb_decoder(16#b8#)) OR
 					(reg_q703 AND symb_decoder(16#a9#)) OR
 					(reg_q703 AND symb_decoder(16#07#)) OR
 					(reg_q703 AND symb_decoder(16#91#)) OR
 					(reg_q703 AND symb_decoder(16#62#)) OR
 					(reg_q703 AND symb_decoder(16#cf#)) OR
 					(reg_q703 AND symb_decoder(16#8c#)) OR
 					(reg_q703 AND symb_decoder(16#7b#)) OR
 					(reg_q703 AND symb_decoder(16#8a#)) OR
 					(reg_q703 AND symb_decoder(16#80#)) OR
 					(reg_q703 AND symb_decoder(16#42#)) OR
 					(reg_q703 AND symb_decoder(16#87#)) OR
 					(reg_q703 AND symb_decoder(16#bc#)) OR
 					(reg_q703 AND symb_decoder(16#36#)) OR
 					(reg_q703 AND symb_decoder(16#9e#)) OR
 					(reg_q703 AND symb_decoder(16#7c#)) OR
 					(reg_q703 AND symb_decoder(16#1b#)) OR
 					(reg_q703 AND symb_decoder(16#70#)) OR
 					(reg_q703 AND symb_decoder(16#71#)) OR
 					(reg_q703 AND symb_decoder(16#a2#)) OR
 					(reg_q703 AND symb_decoder(16#f3#)) OR
 					(reg_q703 AND symb_decoder(16#41#)) OR
 					(reg_q703 AND symb_decoder(16#51#)) OR
 					(reg_q703 AND symb_decoder(16#e9#)) OR
 					(reg_q703 AND symb_decoder(16#f1#)) OR
 					(reg_q703 AND symb_decoder(16#a7#)) OR
 					(reg_q703 AND symb_decoder(16#9c#)) OR
 					(reg_q703 AND symb_decoder(16#1e#)) OR
 					(reg_q703 AND symb_decoder(16#4f#)) OR
 					(reg_q703 AND symb_decoder(16#69#)) OR
 					(reg_q703 AND symb_decoder(16#54#)) OR
 					(reg_q703 AND symb_decoder(16#93#)) OR
 					(reg_q703 AND symb_decoder(16#2b#)) OR
 					(reg_q703 AND symb_decoder(16#eb#)) OR
 					(reg_q703 AND symb_decoder(16#30#)) OR
 					(reg_q703 AND symb_decoder(16#47#)) OR
 					(reg_q703 AND symb_decoder(16#e8#)) OR
 					(reg_q703 AND symb_decoder(16#dc#)) OR
 					(reg_q703 AND symb_decoder(16#73#)) OR
 					(reg_q703 AND symb_decoder(16#63#)) OR
 					(reg_q703 AND symb_decoder(16#a1#)) OR
 					(reg_q703 AND symb_decoder(16#da#)) OR
 					(reg_q703 AND symb_decoder(16#c8#)) OR
 					(reg_q703 AND symb_decoder(16#52#)) OR
 					(reg_q703 AND symb_decoder(16#53#)) OR
 					(reg_q703 AND symb_decoder(16#ef#)) OR
 					(reg_q703 AND symb_decoder(16#75#)) OR
 					(reg_q703 AND symb_decoder(16#56#)) OR
 					(reg_q703 AND symb_decoder(16#c1#)) OR
 					(reg_q703 AND symb_decoder(16#d8#)) OR
 					(reg_q703 AND symb_decoder(16#2a#)) OR
 					(reg_q703 AND symb_decoder(16#68#)) OR
 					(reg_q703 AND symb_decoder(16#0e#)) OR
 					(reg_q703 AND symb_decoder(16#9a#)) OR
 					(reg_q703 AND symb_decoder(16#3a#)) OR
 					(reg_q703 AND symb_decoder(16#43#)) OR
 					(reg_q703 AND symb_decoder(16#0a#)) OR
 					(reg_q703 AND symb_decoder(16#d2#)) OR
 					(reg_q703 AND symb_decoder(16#10#)) OR
 					(reg_q703 AND symb_decoder(16#d4#)) OR
 					(reg_q703 AND symb_decoder(16#92#)) OR
 					(reg_q703 AND symb_decoder(16#8b#)) OR
 					(reg_q703 AND symb_decoder(16#dd#)) OR
 					(reg_q703 AND symb_decoder(16#18#)) OR
 					(reg_q703 AND symb_decoder(16#b7#)) OR
 					(reg_q703 AND symb_decoder(16#5d#)) OR
 					(reg_q703 AND symb_decoder(16#a0#)) OR
 					(reg_q703 AND symb_decoder(16#9d#)) OR
 					(reg_q703 AND symb_decoder(16#4c#)) OR
 					(reg_q703 AND symb_decoder(16#f8#)) OR
 					(reg_q703 AND symb_decoder(16#3e#)) OR
 					(reg_q703 AND symb_decoder(16#17#)) OR
 					(reg_q703 AND symb_decoder(16#1c#)) OR
 					(reg_q703 AND symb_decoder(16#f6#)) OR
 					(reg_q703 AND symb_decoder(16#c5#)) OR
 					(reg_q703 AND symb_decoder(16#4d#)) OR
 					(reg_q703 AND symb_decoder(16#be#)) OR
 					(reg_q703 AND symb_decoder(16#48#)) OR
 					(reg_q703 AND symb_decoder(16#19#)) OR
 					(reg_q703 AND symb_decoder(16#e5#)) OR
 					(reg_q703 AND symb_decoder(16#5f#)) OR
 					(reg_q703 AND symb_decoder(16#c7#)) OR
 					(reg_q703 AND symb_decoder(16#e1#)) OR
 					(reg_q703 AND symb_decoder(16#a4#)) OR
 					(reg_q703 AND symb_decoder(16#c0#)) OR
 					(reg_q703 AND symb_decoder(16#af#)) OR
 					(reg_q703 AND symb_decoder(16#28#)) OR
 					(reg_q703 AND symb_decoder(16#ea#)) OR
 					(reg_q703 AND symb_decoder(16#d5#)) OR
 					(reg_q703 AND symb_decoder(16#3c#)) OR
 					(reg_q703 AND symb_decoder(16#1d#)) OR
 					(reg_q703 AND symb_decoder(16#59#)) OR
 					(reg_q703 AND symb_decoder(16#74#)) OR
 					(reg_q703 AND symb_decoder(16#02#)) OR
 					(reg_q703 AND symb_decoder(16#ce#)) OR
 					(reg_q703 AND symb_decoder(16#16#)) OR
 					(reg_q703 AND symb_decoder(16#64#)) OR
 					(reg_q703 AND symb_decoder(16#50#)) OR
 					(reg_q703 AND symb_decoder(16#b1#)) OR
 					(reg_q703 AND symb_decoder(16#d7#)) OR
 					(reg_q703 AND symb_decoder(16#f7#)) OR
 					(reg_q703 AND symb_decoder(16#6c#)) OR
 					(reg_q703 AND symb_decoder(16#78#)) OR
 					(reg_q703 AND symb_decoder(16#e0#)) OR
 					(reg_q703 AND symb_decoder(16#cd#)) OR
 					(reg_q703 AND symb_decoder(16#cb#)) OR
 					(reg_q703 AND symb_decoder(16#66#)) OR
 					(reg_q703 AND symb_decoder(16#e4#)) OR
 					(reg_q703 AND symb_decoder(16#bd#)) OR
 					(reg_q703 AND symb_decoder(16#04#)) OR
 					(reg_q703 AND symb_decoder(16#81#)) OR
 					(reg_q703 AND symb_decoder(16#2f#)) OR
 					(reg_q703 AND symb_decoder(16#ae#)) OR
 					(reg_q703 AND symb_decoder(16#fc#)) OR
 					(reg_q703 AND symb_decoder(16#6e#)) OR
 					(reg_q703 AND symb_decoder(16#61#)) OR
 					(reg_q703 AND symb_decoder(16#ff#)) OR
 					(reg_q703 AND symb_decoder(16#b5#)) OR
 					(reg_q703 AND symb_decoder(16#38#)) OR
 					(reg_q703 AND symb_decoder(16#8d#)) OR
 					(reg_q703 AND symb_decoder(16#55#)) OR
 					(reg_q703 AND symb_decoder(16#96#)) OR
 					(reg_q703 AND symb_decoder(16#82#)) OR
 					(reg_q703 AND symb_decoder(16#bb#)) OR
 					(reg_q703 AND symb_decoder(16#f9#)) OR
 					(reg_q703 AND symb_decoder(16#a8#)) OR
 					(reg_q703 AND symb_decoder(16#77#)) OR
 					(reg_q703 AND symb_decoder(16#7d#)) OR
 					(reg_q703 AND symb_decoder(16#83#)) OR
 					(reg_q703 AND symb_decoder(16#4a#)) OR
 					(reg_q703 AND symb_decoder(16#f0#)) OR
 					(reg_q703 AND symb_decoder(16#23#)) OR
 					(reg_q703 AND symb_decoder(16#3f#)) OR
 					(reg_q703 AND symb_decoder(16#57#)) OR
 					(reg_q703 AND symb_decoder(16#c4#)) OR
 					(reg_q703 AND symb_decoder(16#97#)) OR
 					(reg_q703 AND symb_decoder(16#d6#)) OR
 					(reg_q703 AND symb_decoder(16#98#)) OR
 					(reg_q703 AND symb_decoder(16#bf#)) OR
 					(reg_q703 AND symb_decoder(16#b0#)) OR
 					(reg_q703 AND symb_decoder(16#ab#)) OR
 					(reg_q703 AND symb_decoder(16#26#)) OR
 					(reg_q703 AND symb_decoder(16#89#)) OR
 					(reg_q703 AND symb_decoder(16#fd#)) OR
 					(reg_q703 AND symb_decoder(16#3d#)) OR
 					(reg_q703 AND symb_decoder(16#21#)) OR
 					(reg_q703 AND symb_decoder(16#67#)) OR
 					(reg_q703 AND symb_decoder(16#20#)) OR
 					(reg_q703 AND symb_decoder(16#5b#)) OR
 					(reg_q703 AND symb_decoder(16#ba#)) OR
 					(reg_q703 AND symb_decoder(16#34#)) OR
 					(reg_q703 AND symb_decoder(16#08#)) OR
 					(reg_q703 AND symb_decoder(16#6f#)) OR
 					(reg_q703 AND symb_decoder(16#15#)) OR
 					(reg_q703 AND symb_decoder(16#ec#)) OR
 					(reg_q703 AND symb_decoder(16#44#)) OR
 					(reg_q703 AND symb_decoder(16#a3#)) OR
 					(reg_q703 AND symb_decoder(16#cc#)) OR
 					(reg_q703 AND symb_decoder(16#d0#)) OR
 					(reg_q703 AND symb_decoder(16#c9#)) OR
 					(reg_q703 AND symb_decoder(16#49#)) OR
 					(reg_q703 AND symb_decoder(16#d9#)) OR
 					(reg_q703 AND symb_decoder(16#fe#)) OR
 					(reg_q703 AND symb_decoder(16#b4#)) OR
 					(reg_q703 AND symb_decoder(16#6a#)) OR
 					(reg_q703 AND symb_decoder(16#f2#)) OR
 					(reg_q703 AND symb_decoder(16#2e#)) OR
 					(reg_q703 AND symb_decoder(16#7f#)) OR
 					(reg_q703 AND symb_decoder(16#aa#)) OR
 					(reg_q703 AND symb_decoder(16#9b#)) OR
 					(reg_q703 AND symb_decoder(16#72#)) OR
 					(reg_q703 AND symb_decoder(16#f4#)) OR
 					(reg_q703 AND symb_decoder(16#b6#)) OR
 					(reg_q703 AND symb_decoder(16#13#)) OR
 					(reg_q703 AND symb_decoder(16#de#)) OR
 					(reg_q703 AND symb_decoder(16#6b#)) OR
 					(reg_q703 AND symb_decoder(16#c3#)) OR
 					(reg_q703 AND symb_decoder(16#39#)) OR
 					(reg_q703 AND symb_decoder(16#e6#)) OR
 					(reg_q703 AND symb_decoder(16#fa#)) OR
 					(reg_q703 AND symb_decoder(16#c6#)) OR
 					(reg_q703 AND symb_decoder(16#a6#)) OR
 					(reg_q703 AND symb_decoder(16#25#)) OR
 					(reg_q703 AND symb_decoder(16#6d#)) OR
 					(reg_q703 AND symb_decoder(16#d1#)) OR
 					(reg_q703 AND symb_decoder(16#94#)) OR
 					(reg_q703 AND symb_decoder(16#0b#)) OR
 					(reg_q703 AND symb_decoder(16#27#)) OR
 					(reg_q703 AND symb_decoder(16#76#)) OR
 					(reg_q703 AND symb_decoder(16#ca#)) OR
 					(reg_q703 AND symb_decoder(16#5a#)) OR
 					(reg_q703 AND symb_decoder(16#e2#)) OR
 					(reg_q703 AND symb_decoder(16#fb#)) OR
 					(reg_q703 AND symb_decoder(16#35#)) OR
 					(reg_q703 AND symb_decoder(16#14#)) OR
 					(reg_q703 AND symb_decoder(16#9f#)) OR
 					(reg_q703 AND symb_decoder(16#37#)) OR
 					(reg_q703 AND symb_decoder(16#0c#)) OR
 					(reg_q703 AND symb_decoder(16#45#)) OR
 					(reg_q703 AND symb_decoder(16#0f#)) OR
 					(reg_q703 AND symb_decoder(16#31#)) OR
 					(reg_q703 AND symb_decoder(16#03#)) OR
 					(reg_q703 AND symb_decoder(16#01#)) OR
 					(reg_q703 AND symb_decoder(16#65#)) OR
 					(reg_q703 AND symb_decoder(16#24#)) OR
 					(reg_q703 AND symb_decoder(16#33#)) OR
 					(reg_q703 AND symb_decoder(16#11#)) OR
 					(reg_q703 AND symb_decoder(16#4e#)) OR
 					(reg_q703 AND symb_decoder(16#22#)) OR
 					(reg_q703 AND symb_decoder(16#b9#)) OR
 					(reg_q703 AND symb_decoder(16#2c#)) OR
 					(reg_q703 AND symb_decoder(16#ee#)) OR
 					(reg_q703 AND symb_decoder(16#e7#)) OR
 					(reg_q703 AND symb_decoder(16#db#)) OR
 					(reg_q703 AND symb_decoder(16#5c#)) OR
 					(reg_q703 AND symb_decoder(16#79#)) OR
 					(reg_q703 AND symb_decoder(16#d3#)) OR
 					(reg_q703 AND symb_decoder(16#05#)) OR
 					(reg_q703 AND symb_decoder(16#86#)) OR
 					(reg_q703 AND symb_decoder(16#b2#)) OR
 					(reg_q703 AND symb_decoder(16#f5#)) OR
 					(reg_q703 AND symb_decoder(16#58#)) OR
 					(reg_q703 AND symb_decoder(16#c2#)) OR
 					(reg_q703 AND symb_decoder(16#06#)) OR
 					(reg_q703 AND symb_decoder(16#99#)) OR
 					(reg_q703 AND symb_decoder(16#85#)) OR
 					(reg_q703 AND symb_decoder(16#3b#)) OR
 					(reg_q703 AND symb_decoder(16#2d#)) OR
 					(reg_q703 AND symb_decoder(16#ac#)) OR
 					(reg_q703 AND symb_decoder(16#00#)) OR
 					(reg_q703 AND symb_decoder(16#84#)) OR
 					(reg_q703 AND symb_decoder(16#12#)) OR
 					(reg_q703 AND symb_decoder(16#ed#)) OR
 					(reg_q703 AND symb_decoder(16#7e#)) OR
 					(reg_q703 AND symb_decoder(16#88#)) OR
 					(reg_q703 AND symb_decoder(16#7a#)) OR
 					(reg_q703 AND symb_decoder(16#60#)) OR
 					(reg_q703 AND symb_decoder(16#32#)) OR
 					(reg_q703 AND symb_decoder(16#09#)) OR
 					(reg_q703 AND symb_decoder(16#1a#)) OR
 					(reg_q703 AND symb_decoder(16#b3#));
reg_q703_init <= '0' ;
	p_reg_q703: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q703 <= reg_q703_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q703 <= reg_q703_init;
        else
          reg_q703 <= reg_q703_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1574_in <= (reg_q1574 AND symb_decoder(16#0c#)) OR
 					(reg_q1574 AND symb_decoder(16#20#)) OR
 					(reg_q1574 AND symb_decoder(16#0d#)) OR
 					(reg_q1574 AND symb_decoder(16#0a#)) OR
 					(reg_q1574 AND symb_decoder(16#09#)) OR
 					(reg_q1572 AND symb_decoder(16#09#)) OR
 					(reg_q1572 AND symb_decoder(16#20#)) OR
 					(reg_q1572 AND symb_decoder(16#0c#)) OR
 					(reg_q1572 AND symb_decoder(16#0a#)) OR
 					(reg_q1572 AND symb_decoder(16#0d#));
reg_q1574_init <= '0' ;
	p_reg_q1574: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1574 <= reg_q1574_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1574 <= reg_q1574_init;
        else
          reg_q1574 <= reg_q1574_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1576_in <= (reg_q1574 AND symb_decoder(16#34#)) OR
 					(reg_q1574 AND symb_decoder(16#32#)) OR
 					(reg_q1574 AND symb_decoder(16#33#)) OR
 					(reg_q1574 AND symb_decoder(16#35#)) OR
 					(reg_q1574 AND symb_decoder(16#31#)) OR
 					(reg_q1574 AND symb_decoder(16#36#)) OR
 					(reg_q1574 AND symb_decoder(16#37#)) OR
 					(reg_q1574 AND symb_decoder(16#38#)) OR
 					(reg_q1574 AND symb_decoder(16#39#)) OR
 					(reg_q1574 AND symb_decoder(16#30#)) OR
 					(reg_q1576 AND symb_decoder(16#30#)) OR
 					(reg_q1576 AND symb_decoder(16#33#)) OR
 					(reg_q1576 AND symb_decoder(16#37#)) OR
 					(reg_q1576 AND symb_decoder(16#35#)) OR
 					(reg_q1576 AND symb_decoder(16#32#)) OR
 					(reg_q1576 AND symb_decoder(16#34#)) OR
 					(reg_q1576 AND symb_decoder(16#39#)) OR
 					(reg_q1576 AND symb_decoder(16#31#)) OR
 					(reg_q1576 AND symb_decoder(16#36#)) OR
 					(reg_q1576 AND symb_decoder(16#38#));
reg_q1576_init <= '0' ;
	p_reg_q1576: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1576 <= reg_q1576_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1576 <= reg_q1576_init;
        else
          reg_q1576 <= reg_q1576_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2172_in <= (reg_q2170 AND symb_decoder(16#4e#)) OR
 					(reg_q2170 AND symb_decoder(16#6e#));
reg_q2172_init <= '0' ;
	p_reg_q2172: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2172 <= reg_q2172_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2172 <= reg_q2172_init;
        else
          reg_q2172 <= reg_q2172_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2208_in <= (reg_q2172 AND symb_decoder(16#41#)) OR
 					(reg_q2172 AND symb_decoder(16#e7#)) OR
 					(reg_q2172 AND symb_decoder(16#7e#)) OR
 					(reg_q2172 AND symb_decoder(16#0e#)) OR
 					(reg_q2172 AND symb_decoder(16#0f#)) OR
 					(reg_q2172 AND symb_decoder(16#d7#)) OR
 					(reg_q2172 AND symb_decoder(16#e2#)) OR
 					(reg_q2172 AND symb_decoder(16#80#)) OR
 					(reg_q2172 AND symb_decoder(16#2f#)) OR
 					(reg_q2172 AND symb_decoder(16#12#)) OR
 					(reg_q2172 AND symb_decoder(16#b8#)) OR
 					(reg_q2172 AND symb_decoder(16#be#)) OR
 					(reg_q2172 AND symb_decoder(16#c9#)) OR
 					(reg_q2172 AND symb_decoder(16#6d#)) OR
 					(reg_q2172 AND symb_decoder(16#af#)) OR
 					(reg_q2172 AND symb_decoder(16#7c#)) OR
 					(reg_q2172 AND symb_decoder(16#e0#)) OR
 					(reg_q2172 AND symb_decoder(16#35#)) OR
 					(reg_q2172 AND symb_decoder(16#a2#)) OR
 					(reg_q2172 AND symb_decoder(16#89#)) OR
 					(reg_q2172 AND symb_decoder(16#27#)) OR
 					(reg_q2172 AND symb_decoder(16#3d#)) OR
 					(reg_q2172 AND symb_decoder(16#56#)) OR
 					(reg_q2172 AND symb_decoder(16#e9#)) OR
 					(reg_q2172 AND symb_decoder(16#97#)) OR
 					(reg_q2172 AND symb_decoder(16#40#)) OR
 					(reg_q2172 AND symb_decoder(16#9d#)) OR
 					(reg_q2172 AND symb_decoder(16#76#)) OR
 					(reg_q2172 AND symb_decoder(16#6b#)) OR
 					(reg_q2172 AND symb_decoder(16#02#)) OR
 					(reg_q2172 AND symb_decoder(16#d5#)) OR
 					(reg_q2172 AND symb_decoder(16#95#)) OR
 					(reg_q2172 AND symb_decoder(16#05#)) OR
 					(reg_q2172 AND symb_decoder(16#ce#)) OR
 					(reg_q2172 AND symb_decoder(16#64#)) OR
 					(reg_q2172 AND symb_decoder(16#98#)) OR
 					(reg_q2172 AND symb_decoder(16#f7#)) OR
 					(reg_q2172 AND symb_decoder(16#83#)) OR
 					(reg_q2172 AND symb_decoder(16#54#)) OR
 					(reg_q2172 AND symb_decoder(16#a3#)) OR
 					(reg_q2172 AND symb_decoder(16#43#)) OR
 					(reg_q2172 AND symb_decoder(16#e1#)) OR
 					(reg_q2172 AND symb_decoder(16#67#)) OR
 					(reg_q2172 AND symb_decoder(16#24#)) OR
 					(reg_q2172 AND symb_decoder(16#e6#)) OR
 					(reg_q2172 AND symb_decoder(16#ac#)) OR
 					(reg_q2172 AND symb_decoder(16#cf#)) OR
 					(reg_q2172 AND symb_decoder(16#fe#)) OR
 					(reg_q2172 AND symb_decoder(16#69#)) OR
 					(reg_q2172 AND symb_decoder(16#dc#)) OR
 					(reg_q2172 AND symb_decoder(16#a0#)) OR
 					(reg_q2172 AND symb_decoder(16#07#)) OR
 					(reg_q2172 AND symb_decoder(16#3e#)) OR
 					(reg_q2172 AND symb_decoder(16#44#)) OR
 					(reg_q2172 AND symb_decoder(16#2b#)) OR
 					(reg_q2172 AND symb_decoder(16#09#)) OR
 					(reg_q2172 AND symb_decoder(16#3a#)) OR
 					(reg_q2172 AND symb_decoder(16#8a#)) OR
 					(reg_q2172 AND symb_decoder(16#66#)) OR
 					(reg_q2172 AND symb_decoder(16#78#)) OR
 					(reg_q2172 AND symb_decoder(16#5f#)) OR
 					(reg_q2172 AND symb_decoder(16#bd#)) OR
 					(reg_q2172 AND symb_decoder(16#aa#)) OR
 					(reg_q2172 AND symb_decoder(16#c1#)) OR
 					(reg_q2172 AND symb_decoder(16#f6#)) OR
 					(reg_q2172 AND symb_decoder(16#4a#)) OR
 					(reg_q2172 AND symb_decoder(16#85#)) OR
 					(reg_q2172 AND symb_decoder(16#a8#)) OR
 					(reg_q2172 AND symb_decoder(16#90#)) OR
 					(reg_q2172 AND symb_decoder(16#03#)) OR
 					(reg_q2172 AND symb_decoder(16#5e#)) OR
 					(reg_q2172 AND symb_decoder(16#1a#)) OR
 					(reg_q2172 AND symb_decoder(16#0d#)) OR
 					(reg_q2172 AND symb_decoder(16#29#)) OR
 					(reg_q2172 AND symb_decoder(16#c0#)) OR
 					(reg_q2172 AND symb_decoder(16#5a#)) OR
 					(reg_q2172 AND symb_decoder(16#5d#)) OR
 					(reg_q2172 AND symb_decoder(16#59#)) OR
 					(reg_q2172 AND symb_decoder(16#b2#)) OR
 					(reg_q2172 AND symb_decoder(16#30#)) OR
 					(reg_q2172 AND symb_decoder(16#8d#)) OR
 					(reg_q2172 AND symb_decoder(16#c4#)) OR
 					(reg_q2172 AND symb_decoder(16#9e#)) OR
 					(reg_q2172 AND symb_decoder(16#46#)) OR
 					(reg_q2172 AND symb_decoder(16#d1#)) OR
 					(reg_q2172 AND symb_decoder(16#b6#)) OR
 					(reg_q2172 AND symb_decoder(16#df#)) OR
 					(reg_q2172 AND symb_decoder(16#c3#)) OR
 					(reg_q2172 AND symb_decoder(16#ea#)) OR
 					(reg_q2172 AND symb_decoder(16#18#)) OR
 					(reg_q2172 AND symb_decoder(16#9b#)) OR
 					(reg_q2172 AND symb_decoder(16#06#)) OR
 					(reg_q2172 AND symb_decoder(16#6c#)) OR
 					(reg_q2172 AND symb_decoder(16#74#)) OR
 					(reg_q2172 AND symb_decoder(16#f3#)) OR
 					(reg_q2172 AND symb_decoder(16#33#)) OR
 					(reg_q2172 AND symb_decoder(16#4b#)) OR
 					(reg_q2172 AND symb_decoder(16#bc#)) OR
 					(reg_q2172 AND symb_decoder(16#ec#)) OR
 					(reg_q2172 AND symb_decoder(16#f0#)) OR
 					(reg_q2172 AND symb_decoder(16#45#)) OR
 					(reg_q2172 AND symb_decoder(16#3f#)) OR
 					(reg_q2172 AND symb_decoder(16#a9#)) OR
 					(reg_q2172 AND symb_decoder(16#73#)) OR
 					(reg_q2172 AND symb_decoder(16#9a#)) OR
 					(reg_q2172 AND symb_decoder(16#38#)) OR
 					(reg_q2172 AND symb_decoder(16#fc#)) OR
 					(reg_q2172 AND symb_decoder(16#cb#)) OR
 					(reg_q2172 AND symb_decoder(16#0b#)) OR
 					(reg_q2172 AND symb_decoder(16#4f#)) OR
 					(reg_q2172 AND symb_decoder(16#d8#)) OR
 					(reg_q2172 AND symb_decoder(16#58#)) OR
 					(reg_q2172 AND symb_decoder(16#16#)) OR
 					(reg_q2172 AND symb_decoder(16#2d#)) OR
 					(reg_q2172 AND symb_decoder(16#75#)) OR
 					(reg_q2172 AND symb_decoder(16#2e#)) OR
 					(reg_q2172 AND symb_decoder(16#7b#)) OR
 					(reg_q2172 AND symb_decoder(16#b9#)) OR
 					(reg_q2172 AND symb_decoder(16#7d#)) OR
 					(reg_q2172 AND symb_decoder(16#01#)) OR
 					(reg_q2172 AND symb_decoder(16#17#)) OR
 					(reg_q2172 AND symb_decoder(16#25#)) OR
 					(reg_q2172 AND symb_decoder(16#d3#)) OR
 					(reg_q2172 AND symb_decoder(16#13#)) OR
 					(reg_q2172 AND symb_decoder(16#47#)) OR
 					(reg_q2172 AND symb_decoder(16#0a#)) OR
 					(reg_q2172 AND symb_decoder(16#31#)) OR
 					(reg_q2172 AND symb_decoder(16#1d#)) OR
 					(reg_q2172 AND symb_decoder(16#57#)) OR
 					(reg_q2172 AND symb_decoder(16#94#)) OR
 					(reg_q2172 AND symb_decoder(16#65#)) OR
 					(reg_q2172 AND symb_decoder(16#84#)) OR
 					(reg_q2172 AND symb_decoder(16#68#)) OR
 					(reg_q2172 AND symb_decoder(16#99#)) OR
 					(reg_q2172 AND symb_decoder(16#21#)) OR
 					(reg_q2172 AND symb_decoder(16#5b#)) OR
 					(reg_q2172 AND symb_decoder(16#60#)) OR
 					(reg_q2172 AND symb_decoder(16#79#)) OR
 					(reg_q2172 AND symb_decoder(16#ab#)) OR
 					(reg_q2172 AND symb_decoder(16#88#)) OR
 					(reg_q2172 AND symb_decoder(16#de#)) OR
 					(reg_q2172 AND symb_decoder(16#dd#)) OR
 					(reg_q2172 AND symb_decoder(16#91#)) OR
 					(reg_q2172 AND symb_decoder(16#87#)) OR
 					(reg_q2172 AND symb_decoder(16#ad#)) OR
 					(reg_q2172 AND symb_decoder(16#bb#)) OR
 					(reg_q2172 AND symb_decoder(16#1e#)) OR
 					(reg_q2172 AND symb_decoder(16#a7#)) OR
 					(reg_q2172 AND symb_decoder(16#a1#)) OR
 					(reg_q2172 AND symb_decoder(16#42#)) OR
 					(reg_q2172 AND symb_decoder(16#8b#)) OR
 					(reg_q2172 AND symb_decoder(16#26#)) OR
 					(reg_q2172 AND symb_decoder(16#8e#)) OR
 					(reg_q2172 AND symb_decoder(16#e5#)) OR
 					(reg_q2172 AND symb_decoder(16#e4#)) OR
 					(reg_q2172 AND symb_decoder(16#b0#)) OR
 					(reg_q2172 AND symb_decoder(16#ba#)) OR
 					(reg_q2172 AND symb_decoder(16#eb#)) OR
 					(reg_q2172 AND symb_decoder(16#3b#)) OR
 					(reg_q2172 AND symb_decoder(16#c7#)) OR
 					(reg_q2172 AND symb_decoder(16#04#)) OR
 					(reg_q2172 AND symb_decoder(16#ed#)) OR
 					(reg_q2172 AND symb_decoder(16#82#)) OR
 					(reg_q2172 AND symb_decoder(16#39#)) OR
 					(reg_q2172 AND symb_decoder(16#28#)) OR
 					(reg_q2172 AND symb_decoder(16#f4#)) OR
 					(reg_q2172 AND symb_decoder(16#f8#)) OR
 					(reg_q2172 AND symb_decoder(16#3c#)) OR
 					(reg_q2172 AND symb_decoder(16#b5#)) OR
 					(reg_q2172 AND symb_decoder(16#14#)) OR
 					(reg_q2172 AND symb_decoder(16#bf#)) OR
 					(reg_q2172 AND symb_decoder(16#1b#)) OR
 					(reg_q2172 AND symb_decoder(16#ae#)) OR
 					(reg_q2172 AND symb_decoder(16#77#)) OR
 					(reg_q2172 AND symb_decoder(16#7a#)) OR
 					(reg_q2172 AND symb_decoder(16#f9#)) OR
 					(reg_q2172 AND symb_decoder(16#da#)) OR
 					(reg_q2172 AND symb_decoder(16#fd#)) OR
 					(reg_q2172 AND symb_decoder(16#2c#)) OR
 					(reg_q2172 AND symb_decoder(16#37#)) OR
 					(reg_q2172 AND symb_decoder(16#51#)) OR
 					(reg_q2172 AND symb_decoder(16#2a#)) OR
 					(reg_q2172 AND symb_decoder(16#f5#)) OR
 					(reg_q2172 AND symb_decoder(16#81#)) OR
 					(reg_q2172 AND symb_decoder(16#cd#)) OR
 					(reg_q2172 AND symb_decoder(16#08#)) OR
 					(reg_q2172 AND symb_decoder(16#15#)) OR
 					(reg_q2172 AND symb_decoder(16#d6#)) OR
 					(reg_q2172 AND symb_decoder(16#a5#)) OR
 					(reg_q2172 AND symb_decoder(16#a4#)) OR
 					(reg_q2172 AND symb_decoder(16#72#)) OR
 					(reg_q2172 AND symb_decoder(16#4d#)) OR
 					(reg_q2172 AND symb_decoder(16#50#)) OR
 					(reg_q2172 AND symb_decoder(16#d0#)) OR
 					(reg_q2172 AND symb_decoder(16#c2#)) OR
 					(reg_q2172 AND symb_decoder(16#48#)) OR
 					(reg_q2172 AND symb_decoder(16#0c#)) OR
 					(reg_q2172 AND symb_decoder(16#6a#)) OR
 					(reg_q2172 AND symb_decoder(16#23#)) OR
 					(reg_q2172 AND symb_decoder(16#49#)) OR
 					(reg_q2172 AND symb_decoder(16#fb#)) OR
 					(reg_q2172 AND symb_decoder(16#34#)) OR
 					(reg_q2172 AND symb_decoder(16#4e#)) OR
 					(reg_q2172 AND symb_decoder(16#55#)) OR
 					(reg_q2172 AND symb_decoder(16#d4#)) OR
 					(reg_q2172 AND symb_decoder(16#11#)) OR
 					(reg_q2172 AND symb_decoder(16#32#)) OR
 					(reg_q2172 AND symb_decoder(16#1f#)) OR
 					(reg_q2172 AND symb_decoder(16#61#)) OR
 					(reg_q2172 AND symb_decoder(16#e8#)) OR
 					(reg_q2172 AND symb_decoder(16#cc#)) OR
 					(reg_q2172 AND symb_decoder(16#71#)) OR
 					(reg_q2172 AND symb_decoder(16#8c#)) OR
 					(reg_q2172 AND symb_decoder(16#d2#)) OR
 					(reg_q2172 AND symb_decoder(16#19#)) OR
 					(reg_q2172 AND symb_decoder(16#53#)) OR
 					(reg_q2172 AND symb_decoder(16#62#)) OR
 					(reg_q2172 AND symb_decoder(16#e3#)) OR
 					(reg_q2172 AND symb_decoder(16#a6#)) OR
 					(reg_q2172 AND symb_decoder(16#f1#)) OR
 					(reg_q2172 AND symb_decoder(16#fa#)) OR
 					(reg_q2172 AND symb_decoder(16#10#)) OR
 					(reg_q2172 AND symb_decoder(16#4c#)) OR
 					(reg_q2172 AND symb_decoder(16#96#)) OR
 					(reg_q2172 AND symb_decoder(16#c6#)) OR
 					(reg_q2172 AND symb_decoder(16#1c#)) OR
 					(reg_q2172 AND symb_decoder(16#8f#)) OR
 					(reg_q2172 AND symb_decoder(16#f2#)) OR
 					(reg_q2172 AND symb_decoder(16#b3#)) OR
 					(reg_q2172 AND symb_decoder(16#6e#)) OR
 					(reg_q2172 AND symb_decoder(16#c5#)) OR
 					(reg_q2172 AND symb_decoder(16#52#)) OR
 					(reg_q2172 AND symb_decoder(16#ca#)) OR
 					(reg_q2172 AND symb_decoder(16#9c#)) OR
 					(reg_q2172 AND symb_decoder(16#b7#)) OR
 					(reg_q2172 AND symb_decoder(16#63#)) OR
 					(reg_q2172 AND symb_decoder(16#ef#)) OR
 					(reg_q2172 AND symb_decoder(16#b1#)) OR
 					(reg_q2172 AND symb_decoder(16#5c#)) OR
 					(reg_q2172 AND symb_decoder(16#c8#)) OR
 					(reg_q2172 AND symb_decoder(16#36#)) OR
 					(reg_q2172 AND symb_decoder(16#9f#)) OR
 					(reg_q2172 AND symb_decoder(16#d9#)) OR
 					(reg_q2172 AND symb_decoder(16#db#)) OR
 					(reg_q2172 AND symb_decoder(16#20#)) OR
 					(reg_q2172 AND symb_decoder(16#22#)) OR
 					(reg_q2172 AND symb_decoder(16#93#)) OR
 					(reg_q2172 AND symb_decoder(16#00#)) OR
 					(reg_q2172 AND symb_decoder(16#70#)) OR
 					(reg_q2172 AND symb_decoder(16#7f#)) OR
 					(reg_q2172 AND symb_decoder(16#92#)) OR
 					(reg_q2172 AND symb_decoder(16#ff#)) OR
 					(reg_q2172 AND symb_decoder(16#86#)) OR
 					(reg_q2172 AND symb_decoder(16#b4#)) OR
 					(reg_q2172 AND symb_decoder(16#ee#)) OR
 					(reg_q2172 AND symb_decoder(16#6f#)) OR
 					(reg_q2208 AND symb_decoder(16#c0#)) OR
 					(reg_q2208 AND symb_decoder(16#72#)) OR
 					(reg_q2208 AND symb_decoder(16#c7#)) OR
 					(reg_q2208 AND symb_decoder(16#b0#)) OR
 					(reg_q2208 AND symb_decoder(16#d1#)) OR
 					(reg_q2208 AND symb_decoder(16#0e#)) OR
 					(reg_q2208 AND symb_decoder(16#0d#)) OR
 					(reg_q2208 AND symb_decoder(16#5b#)) OR
 					(reg_q2208 AND symb_decoder(16#bf#)) OR
 					(reg_q2208 AND symb_decoder(16#37#)) OR
 					(reg_q2208 AND symb_decoder(16#dd#)) OR
 					(reg_q2208 AND symb_decoder(16#bd#)) OR
 					(reg_q2208 AND symb_decoder(16#08#)) OR
 					(reg_q2208 AND symb_decoder(16#fe#)) OR
 					(reg_q2208 AND symb_decoder(16#54#)) OR
 					(reg_q2208 AND symb_decoder(16#86#)) OR
 					(reg_q2208 AND symb_decoder(16#13#)) OR
 					(reg_q2208 AND symb_decoder(16#0a#)) OR
 					(reg_q2208 AND symb_decoder(16#8a#)) OR
 					(reg_q2208 AND symb_decoder(16#8b#)) OR
 					(reg_q2208 AND symb_decoder(16#22#)) OR
 					(reg_q2208 AND symb_decoder(16#89#)) OR
 					(reg_q2208 AND symb_decoder(16#1f#)) OR
 					(reg_q2208 AND symb_decoder(16#87#)) OR
 					(reg_q2208 AND symb_decoder(16#6f#)) OR
 					(reg_q2208 AND symb_decoder(16#28#)) OR
 					(reg_q2208 AND symb_decoder(16#70#)) OR
 					(reg_q2208 AND symb_decoder(16#4f#)) OR
 					(reg_q2208 AND symb_decoder(16#12#)) OR
 					(reg_q2208 AND symb_decoder(16#af#)) OR
 					(reg_q2208 AND symb_decoder(16#eb#)) OR
 					(reg_q2208 AND symb_decoder(16#f8#)) OR
 					(reg_q2208 AND symb_decoder(16#00#)) OR
 					(reg_q2208 AND symb_decoder(16#7e#)) OR
 					(reg_q2208 AND symb_decoder(16#be#)) OR
 					(reg_q2208 AND symb_decoder(16#f9#)) OR
 					(reg_q2208 AND symb_decoder(16#29#)) OR
 					(reg_q2208 AND symb_decoder(16#25#)) OR
 					(reg_q2208 AND symb_decoder(16#3d#)) OR
 					(reg_q2208 AND symb_decoder(16#c5#)) OR
 					(reg_q2208 AND symb_decoder(16#ef#)) OR
 					(reg_q2208 AND symb_decoder(16#90#)) OR
 					(reg_q2208 AND symb_decoder(16#61#)) OR
 					(reg_q2208 AND symb_decoder(16#9e#)) OR
 					(reg_q2208 AND symb_decoder(16#b9#)) OR
 					(reg_q2208 AND symb_decoder(16#6e#)) OR
 					(reg_q2208 AND symb_decoder(16#ff#)) OR
 					(reg_q2208 AND symb_decoder(16#f2#)) OR
 					(reg_q2208 AND symb_decoder(16#15#)) OR
 					(reg_q2208 AND symb_decoder(16#14#)) OR
 					(reg_q2208 AND symb_decoder(16#ac#)) OR
 					(reg_q2208 AND symb_decoder(16#05#)) OR
 					(reg_q2208 AND symb_decoder(16#75#)) OR
 					(reg_q2208 AND symb_decoder(16#da#)) OR
 					(reg_q2208 AND symb_decoder(16#a0#)) OR
 					(reg_q2208 AND symb_decoder(16#5f#)) OR
 					(reg_q2208 AND symb_decoder(16#51#)) OR
 					(reg_q2208 AND symb_decoder(16#bc#)) OR
 					(reg_q2208 AND symb_decoder(16#2e#)) OR
 					(reg_q2208 AND symb_decoder(16#df#)) OR
 					(reg_q2208 AND symb_decoder(16#91#)) OR
 					(reg_q2208 AND symb_decoder(16#4b#)) OR
 					(reg_q2208 AND symb_decoder(16#41#)) OR
 					(reg_q2208 AND symb_decoder(16#73#)) OR
 					(reg_q2208 AND symb_decoder(16#ea#)) OR
 					(reg_q2208 AND symb_decoder(16#56#)) OR
 					(reg_q2208 AND symb_decoder(16#57#)) OR
 					(reg_q2208 AND symb_decoder(16#a8#)) OR
 					(reg_q2208 AND symb_decoder(16#ee#)) OR
 					(reg_q2208 AND symb_decoder(16#44#)) OR
 					(reg_q2208 AND symb_decoder(16#c6#)) OR
 					(reg_q2208 AND symb_decoder(16#1c#)) OR
 					(reg_q2208 AND symb_decoder(16#66#)) OR
 					(reg_q2208 AND symb_decoder(16#98#)) OR
 					(reg_q2208 AND symb_decoder(16#33#)) OR
 					(reg_q2208 AND symb_decoder(16#db#)) OR
 					(reg_q2208 AND symb_decoder(16#1d#)) OR
 					(reg_q2208 AND symb_decoder(16#5e#)) OR
 					(reg_q2208 AND symb_decoder(16#d3#)) OR
 					(reg_q2208 AND symb_decoder(16#99#)) OR
 					(reg_q2208 AND symb_decoder(16#c8#)) OR
 					(reg_q2208 AND symb_decoder(16#46#)) OR
 					(reg_q2208 AND symb_decoder(16#d5#)) OR
 					(reg_q2208 AND symb_decoder(16#de#)) OR
 					(reg_q2208 AND symb_decoder(16#16#)) OR
 					(reg_q2208 AND symb_decoder(16#d0#)) OR
 					(reg_q2208 AND symb_decoder(16#a9#)) OR
 					(reg_q2208 AND symb_decoder(16#5d#)) OR
 					(reg_q2208 AND symb_decoder(16#62#)) OR
 					(reg_q2208 AND symb_decoder(16#3a#)) OR
 					(reg_q2208 AND symb_decoder(16#65#)) OR
 					(reg_q2208 AND symb_decoder(16#36#)) OR
 					(reg_q2208 AND symb_decoder(16#d7#)) OR
 					(reg_q2208 AND symb_decoder(16#e2#)) OR
 					(reg_q2208 AND symb_decoder(16#9d#)) OR
 					(reg_q2208 AND symb_decoder(16#ec#)) OR
 					(reg_q2208 AND symb_decoder(16#f0#)) OR
 					(reg_q2208 AND symb_decoder(16#21#)) OR
 					(reg_q2208 AND symb_decoder(16#0b#)) OR
 					(reg_q2208 AND symb_decoder(16#9a#)) OR
 					(reg_q2208 AND symb_decoder(16#fc#)) OR
 					(reg_q2208 AND symb_decoder(16#5c#)) OR
 					(reg_q2208 AND symb_decoder(16#ca#)) OR
 					(reg_q2208 AND symb_decoder(16#b4#)) OR
 					(reg_q2208 AND symb_decoder(16#f6#)) OR
 					(reg_q2208 AND symb_decoder(16#7b#)) OR
 					(reg_q2208 AND symb_decoder(16#6b#)) OR
 					(reg_q2208 AND symb_decoder(16#4a#)) OR
 					(reg_q2208 AND symb_decoder(16#e6#)) OR
 					(reg_q2208 AND symb_decoder(16#64#)) OR
 					(reg_q2208 AND symb_decoder(16#93#)) OR
 					(reg_q2208 AND symb_decoder(16#fb#)) OR
 					(reg_q2208 AND symb_decoder(16#e0#)) OR
 					(reg_q2208 AND symb_decoder(16#a5#)) OR
 					(reg_q2208 AND symb_decoder(16#4e#)) OR
 					(reg_q2208 AND symb_decoder(16#3e#)) OR
 					(reg_q2208 AND symb_decoder(16#18#)) OR
 					(reg_q2208 AND symb_decoder(16#d8#)) OR
 					(reg_q2208 AND symb_decoder(16#2a#)) OR
 					(reg_q2208 AND symb_decoder(16#35#)) OR
 					(reg_q2208 AND symb_decoder(16#e3#)) OR
 					(reg_q2208 AND symb_decoder(16#cd#)) OR
 					(reg_q2208 AND symb_decoder(16#e4#)) OR
 					(reg_q2208 AND symb_decoder(16#81#)) OR
 					(reg_q2208 AND symb_decoder(16#85#)) OR
 					(reg_q2208 AND symb_decoder(16#8f#)) OR
 					(reg_q2208 AND symb_decoder(16#80#)) OR
 					(reg_q2208 AND symb_decoder(16#84#)) OR
 					(reg_q2208 AND symb_decoder(16#aa#)) OR
 					(reg_q2208 AND symb_decoder(16#d4#)) OR
 					(reg_q2208 AND symb_decoder(16#3b#)) OR
 					(reg_q2208 AND symb_decoder(16#ed#)) OR
 					(reg_q2208 AND symb_decoder(16#2f#)) OR
 					(reg_q2208 AND symb_decoder(16#88#)) OR
 					(reg_q2208 AND symb_decoder(16#01#)) OR
 					(reg_q2208 AND symb_decoder(16#2d#)) OR
 					(reg_q2208 AND symb_decoder(16#24#)) OR
 					(reg_q2208 AND symb_decoder(16#d6#)) OR
 					(reg_q2208 AND symb_decoder(16#1a#)) OR
 					(reg_q2208 AND symb_decoder(16#ba#)) OR
 					(reg_q2208 AND symb_decoder(16#b6#)) OR
 					(reg_q2208 AND symb_decoder(16#97#)) OR
 					(reg_q2208 AND symb_decoder(16#45#)) OR
 					(reg_q2208 AND symb_decoder(16#49#)) OR
 					(reg_q2208 AND symb_decoder(16#7d#)) OR
 					(reg_q2208 AND symb_decoder(16#b1#)) OR
 					(reg_q2208 AND symb_decoder(16#04#)) OR
 					(reg_q2208 AND symb_decoder(16#68#)) OR
 					(reg_q2208 AND symb_decoder(16#8c#)) OR
 					(reg_q2208 AND symb_decoder(16#c4#)) OR
 					(reg_q2208 AND symb_decoder(16#e7#)) OR
 					(reg_q2208 AND symb_decoder(16#f7#)) OR
 					(reg_q2208 AND symb_decoder(16#cf#)) OR
 					(reg_q2208 AND symb_decoder(16#67#)) OR
 					(reg_q2208 AND symb_decoder(16#e1#)) OR
 					(reg_q2208 AND symb_decoder(16#e9#)) OR
 					(reg_q2208 AND symb_decoder(16#a3#)) OR
 					(reg_q2208 AND symb_decoder(16#cc#)) OR
 					(reg_q2208 AND symb_decoder(16#c1#)) OR
 					(reg_q2208 AND symb_decoder(16#7f#)) OR
 					(reg_q2208 AND symb_decoder(16#17#)) OR
 					(reg_q2208 AND symb_decoder(16#38#)) OR
 					(reg_q2208 AND symb_decoder(16#11#)) OR
 					(reg_q2208 AND symb_decoder(16#02#)) OR
 					(reg_q2208 AND symb_decoder(16#82#)) OR
 					(reg_q2208 AND symb_decoder(16#23#)) OR
 					(reg_q2208 AND symb_decoder(16#43#)) OR
 					(reg_q2208 AND symb_decoder(16#6a#)) OR
 					(reg_q2208 AND symb_decoder(16#26#)) OR
 					(reg_q2208 AND symb_decoder(16#92#)) OR
 					(reg_q2208 AND symb_decoder(16#03#)) OR
 					(reg_q2208 AND symb_decoder(16#47#)) OR
 					(reg_q2208 AND symb_decoder(16#a2#)) OR
 					(reg_q2208 AND symb_decoder(16#d2#)) OR
 					(reg_q2208 AND symb_decoder(16#40#)) OR
 					(reg_q2208 AND symb_decoder(16#79#)) OR
 					(reg_q2208 AND symb_decoder(16#2c#)) OR
 					(reg_q2208 AND symb_decoder(16#95#)) OR
 					(reg_q2208 AND symb_decoder(16#39#)) OR
 					(reg_q2208 AND symb_decoder(16#55#)) OR
 					(reg_q2208 AND symb_decoder(16#83#)) OR
 					(reg_q2208 AND symb_decoder(16#9c#)) OR
 					(reg_q2208 AND symb_decoder(16#a4#)) OR
 					(reg_q2208 AND symb_decoder(16#4c#)) OR
 					(reg_q2208 AND symb_decoder(16#6d#)) OR
 					(reg_q2208 AND symb_decoder(16#94#)) OR
 					(reg_q2208 AND symb_decoder(16#c2#)) OR
 					(reg_q2208 AND symb_decoder(16#8e#)) OR
 					(reg_q2208 AND symb_decoder(16#e5#)) OR
 					(reg_q2208 AND symb_decoder(16#6c#)) OR
 					(reg_q2208 AND symb_decoder(16#a1#)) OR
 					(reg_q2208 AND symb_decoder(16#bb#)) OR
 					(reg_q2208 AND symb_decoder(16#07#)) OR
 					(reg_q2208 AND symb_decoder(16#69#)) OR
 					(reg_q2208 AND symb_decoder(16#fa#)) OR
 					(reg_q2208 AND symb_decoder(16#76#)) OR
 					(reg_q2208 AND symb_decoder(16#7a#)) OR
 					(reg_q2208 AND symb_decoder(16#f3#)) OR
 					(reg_q2208 AND symb_decoder(16#42#)) OR
 					(reg_q2208 AND symb_decoder(16#ad#)) OR
 					(reg_q2208 AND symb_decoder(16#77#)) OR
 					(reg_q2208 AND symb_decoder(16#1e#)) OR
 					(reg_q2208 AND symb_decoder(16#b5#)) OR
 					(reg_q2208 AND symb_decoder(16#59#)) OR
 					(reg_q2208 AND symb_decoder(16#2b#)) OR
 					(reg_q2208 AND symb_decoder(16#20#)) OR
 					(reg_q2208 AND symb_decoder(16#d9#)) OR
 					(reg_q2208 AND symb_decoder(16#58#)) OR
 					(reg_q2208 AND symb_decoder(16#96#)) OR
 					(reg_q2208 AND symb_decoder(16#50#)) OR
 					(reg_q2208 AND symb_decoder(16#9f#)) OR
 					(reg_q2208 AND symb_decoder(16#60#)) OR
 					(reg_q2208 AND symb_decoder(16#53#)) OR
 					(reg_q2208 AND symb_decoder(16#b8#)) OR
 					(reg_q2208 AND symb_decoder(16#a6#)) OR
 					(reg_q2208 AND symb_decoder(16#0f#)) OR
 					(reg_q2208 AND symb_decoder(16#cb#)) OR
 					(reg_q2208 AND symb_decoder(16#a7#)) OR
 					(reg_q2208 AND symb_decoder(16#f1#)) OR
 					(reg_q2208 AND symb_decoder(16#5a#)) OR
 					(reg_q2208 AND symb_decoder(16#06#)) OR
 					(reg_q2208 AND symb_decoder(16#09#)) OR
 					(reg_q2208 AND symb_decoder(16#dc#)) OR
 					(reg_q2208 AND symb_decoder(16#9b#)) OR
 					(reg_q2208 AND symb_decoder(16#74#)) OR
 					(reg_q2208 AND symb_decoder(16#ce#)) OR
 					(reg_q2208 AND symb_decoder(16#63#)) OR
 					(reg_q2208 AND symb_decoder(16#31#)) OR
 					(reg_q2208 AND symb_decoder(16#27#)) OR
 					(reg_q2208 AND symb_decoder(16#7c#)) OR
 					(reg_q2208 AND symb_decoder(16#8d#)) OR
 					(reg_q2208 AND symb_decoder(16#b3#)) OR
 					(reg_q2208 AND symb_decoder(16#b7#)) OR
 					(reg_q2208 AND symb_decoder(16#10#)) OR
 					(reg_q2208 AND symb_decoder(16#4d#)) OR
 					(reg_q2208 AND symb_decoder(16#f5#)) OR
 					(reg_q2208 AND symb_decoder(16#ae#)) OR
 					(reg_q2208 AND symb_decoder(16#78#)) OR
 					(reg_q2208 AND symb_decoder(16#0c#)) OR
 					(reg_q2208 AND symb_decoder(16#71#)) OR
 					(reg_q2208 AND symb_decoder(16#3f#)) OR
 					(reg_q2208 AND symb_decoder(16#e8#)) OR
 					(reg_q2208 AND symb_decoder(16#34#)) OR
 					(reg_q2208 AND symb_decoder(16#19#)) OR
 					(reg_q2208 AND symb_decoder(16#fd#)) OR
 					(reg_q2208 AND symb_decoder(16#1b#)) OR
 					(reg_q2208 AND symb_decoder(16#f4#)) OR
 					(reg_q2208 AND symb_decoder(16#32#)) OR
 					(reg_q2208 AND symb_decoder(16#b2#)) OR
 					(reg_q2208 AND symb_decoder(16#52#)) OR
 					(reg_q2208 AND symb_decoder(16#c3#)) OR
 					(reg_q2208 AND symb_decoder(16#48#)) OR
 					(reg_q2208 AND symb_decoder(16#3c#)) OR
 					(reg_q2208 AND symb_decoder(16#c9#)) OR
 					(reg_q2208 AND symb_decoder(16#ab#)) OR
 					(reg_q2208 AND symb_decoder(16#30#));
reg_q2208_init <= '0' ;
	p_reg_q2208: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2208 <= reg_q2208_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2208 <= reg_q2208_init;
        else
          reg_q2208 <= reg_q2208_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1997_in <= (reg_q1997 AND symb_decoder(16#a3#)) OR
 					(reg_q1997 AND symb_decoder(16#d5#)) OR
 					(reg_q1997 AND symb_decoder(16#a7#)) OR
 					(reg_q1997 AND symb_decoder(16#b8#)) OR
 					(reg_q1997 AND symb_decoder(16#a4#)) OR
 					(reg_q1997 AND symb_decoder(16#45#)) OR
 					(reg_q1997 AND symb_decoder(16#92#)) OR
 					(reg_q1997 AND symb_decoder(16#db#)) OR
 					(reg_q1997 AND symb_decoder(16#22#)) OR
 					(reg_q1997 AND symb_decoder(16#44#)) OR
 					(reg_q1997 AND symb_decoder(16#16#)) OR
 					(reg_q1997 AND symb_decoder(16#d8#)) OR
 					(reg_q1997 AND symb_decoder(16#05#)) OR
 					(reg_q1997 AND symb_decoder(16#26#)) OR
 					(reg_q1997 AND symb_decoder(16#14#)) OR
 					(reg_q1997 AND symb_decoder(16#0b#)) OR
 					(reg_q1997 AND symb_decoder(16#df#)) OR
 					(reg_q1997 AND symb_decoder(16#53#)) OR
 					(reg_q1997 AND symb_decoder(16#b0#)) OR
 					(reg_q1997 AND symb_decoder(16#54#)) OR
 					(reg_q1997 AND symb_decoder(16#40#)) OR
 					(reg_q1997 AND symb_decoder(16#d9#)) OR
 					(reg_q1997 AND symb_decoder(16#50#)) OR
 					(reg_q1997 AND symb_decoder(16#4d#)) OR
 					(reg_q1997 AND symb_decoder(16#73#)) OR
 					(reg_q1997 AND symb_decoder(16#2a#)) OR
 					(reg_q1997 AND symb_decoder(16#76#)) OR
 					(reg_q1997 AND symb_decoder(16#7e#)) OR
 					(reg_q1997 AND symb_decoder(16#8f#)) OR
 					(reg_q1997 AND symb_decoder(16#b9#)) OR
 					(reg_q1997 AND symb_decoder(16#88#)) OR
 					(reg_q1997 AND symb_decoder(16#0e#)) OR
 					(reg_q1997 AND symb_decoder(16#b3#)) OR
 					(reg_q1997 AND symb_decoder(16#83#)) OR
 					(reg_q1997 AND symb_decoder(16#5c#)) OR
 					(reg_q1997 AND symb_decoder(16#08#)) OR
 					(reg_q1997 AND symb_decoder(16#4a#)) OR
 					(reg_q1997 AND symb_decoder(16#91#)) OR
 					(reg_q1997 AND symb_decoder(16#27#)) OR
 					(reg_q1997 AND symb_decoder(16#18#)) OR
 					(reg_q1997 AND symb_decoder(16#9e#)) OR
 					(reg_q1997 AND symb_decoder(16#79#)) OR
 					(reg_q1997 AND symb_decoder(16#ef#)) OR
 					(reg_q1997 AND symb_decoder(16#95#)) OR
 					(reg_q1997 AND symb_decoder(16#b7#)) OR
 					(reg_q1997 AND symb_decoder(16#67#)) OR
 					(reg_q1997 AND symb_decoder(16#31#)) OR
 					(reg_q1997 AND symb_decoder(16#1a#)) OR
 					(reg_q1997 AND symb_decoder(16#37#)) OR
 					(reg_q1997 AND symb_decoder(16#b5#)) OR
 					(reg_q1997 AND symb_decoder(16#5f#)) OR
 					(reg_q1997 AND symb_decoder(16#47#)) OR
 					(reg_q1997 AND symb_decoder(16#15#)) OR
 					(reg_q1997 AND symb_decoder(16#bd#)) OR
 					(reg_q1997 AND symb_decoder(16#25#)) OR
 					(reg_q1997 AND symb_decoder(16#ce#)) OR
 					(reg_q1997 AND symb_decoder(16#d3#)) OR
 					(reg_q1997 AND symb_decoder(16#01#)) OR
 					(reg_q1997 AND symb_decoder(16#d0#)) OR
 					(reg_q1997 AND symb_decoder(16#f3#)) OR
 					(reg_q1997 AND symb_decoder(16#6a#)) OR
 					(reg_q1997 AND symb_decoder(16#fd#)) OR
 					(reg_q1997 AND symb_decoder(16#cc#)) OR
 					(reg_q1997 AND symb_decoder(16#90#)) OR
 					(reg_q1997 AND symb_decoder(16#ba#)) OR
 					(reg_q1997 AND symb_decoder(16#d4#)) OR
 					(reg_q1997 AND symb_decoder(16#a6#)) OR
 					(reg_q1997 AND symb_decoder(16#24#)) OR
 					(reg_q1997 AND symb_decoder(16#bc#)) OR
 					(reg_q1997 AND symb_decoder(16#93#)) OR
 					(reg_q1997 AND symb_decoder(16#11#)) OR
 					(reg_q1997 AND symb_decoder(16#f6#)) OR
 					(reg_q1997 AND symb_decoder(16#f7#)) OR
 					(reg_q1997 AND symb_decoder(16#d2#)) OR
 					(reg_q1997 AND symb_decoder(16#5d#)) OR
 					(reg_q1997 AND symb_decoder(16#63#)) OR
 					(reg_q1997 AND symb_decoder(16#02#)) OR
 					(reg_q1997 AND symb_decoder(16#8b#)) OR
 					(reg_q1997 AND symb_decoder(16#60#)) OR
 					(reg_q1997 AND symb_decoder(16#9f#)) OR
 					(reg_q1997 AND symb_decoder(16#86#)) OR
 					(reg_q1997 AND symb_decoder(16#48#)) OR
 					(reg_q1997 AND symb_decoder(16#cb#)) OR
 					(reg_q1997 AND symb_decoder(16#6f#)) OR
 					(reg_q1997 AND symb_decoder(16#c1#)) OR
 					(reg_q1997 AND symb_decoder(16#9c#)) OR
 					(reg_q1997 AND symb_decoder(16#28#)) OR
 					(reg_q1997 AND symb_decoder(16#0c#)) OR
 					(reg_q1997 AND symb_decoder(16#f9#)) OR
 					(reg_q1997 AND symb_decoder(16#a0#)) OR
 					(reg_q1997 AND symb_decoder(16#a5#)) OR
 					(reg_q1997 AND symb_decoder(16#4e#)) OR
 					(reg_q1997 AND symb_decoder(16#87#)) OR
 					(reg_q1997 AND symb_decoder(16#e2#)) OR
 					(reg_q1997 AND symb_decoder(16#e3#)) OR
 					(reg_q1997 AND symb_decoder(16#2e#)) OR
 					(reg_q1997 AND symb_decoder(16#3a#)) OR
 					(reg_q1997 AND symb_decoder(16#8c#)) OR
 					(reg_q1997 AND symb_decoder(16#10#)) OR
 					(reg_q1997 AND symb_decoder(16#2c#)) OR
 					(reg_q1997 AND symb_decoder(16#3f#)) OR
 					(reg_q1997 AND symb_decoder(16#ae#)) OR
 					(reg_q1997 AND symb_decoder(16#97#)) OR
 					(reg_q1997 AND symb_decoder(16#21#)) OR
 					(reg_q1997 AND symb_decoder(16#29#)) OR
 					(reg_q1997 AND symb_decoder(16#17#)) OR
 					(reg_q1997 AND symb_decoder(16#c8#)) OR
 					(reg_q1997 AND symb_decoder(16#39#)) OR
 					(reg_q1997 AND symb_decoder(16#35#)) OR
 					(reg_q1997 AND symb_decoder(16#6e#)) OR
 					(reg_q1997 AND symb_decoder(16#ff#)) OR
 					(reg_q1997 AND symb_decoder(16#4b#)) OR
 					(reg_q1997 AND symb_decoder(16#13#)) OR
 					(reg_q1997 AND symb_decoder(16#ec#)) OR
 					(reg_q1997 AND symb_decoder(16#3c#)) OR
 					(reg_q1997 AND symb_decoder(16#59#)) OR
 					(reg_q1997 AND symb_decoder(16#ca#)) OR
 					(reg_q1997 AND symb_decoder(16#72#)) OR
 					(reg_q1997 AND symb_decoder(16#64#)) OR
 					(reg_q1997 AND symb_decoder(16#b2#)) OR
 					(reg_q1997 AND symb_decoder(16#84#)) OR
 					(reg_q1997 AND symb_decoder(16#04#)) OR
 					(reg_q1997 AND symb_decoder(16#c4#)) OR
 					(reg_q1997 AND symb_decoder(16#20#)) OR
 					(reg_q1997 AND symb_decoder(16#fc#)) OR
 					(reg_q1997 AND symb_decoder(16#2f#)) OR
 					(reg_q1997 AND symb_decoder(16#e7#)) OR
 					(reg_q1997 AND symb_decoder(16#71#)) OR
 					(reg_q1997 AND symb_decoder(16#cf#)) OR
 					(reg_q1997 AND symb_decoder(16#9b#)) OR
 					(reg_q1997 AND symb_decoder(16#c2#)) OR
 					(reg_q1997 AND symb_decoder(16#e5#)) OR
 					(reg_q1997 AND symb_decoder(16#36#)) OR
 					(reg_q1997 AND symb_decoder(16#65#)) OR
 					(reg_q1997 AND symb_decoder(16#32#)) OR
 					(reg_q1997 AND symb_decoder(16#fa#)) OR
 					(reg_q1997 AND symb_decoder(16#68#)) OR
 					(reg_q1997 AND symb_decoder(16#89#)) OR
 					(reg_q1997 AND symb_decoder(16#19#)) OR
 					(reg_q1997 AND symb_decoder(16#fe#)) OR
 					(reg_q1997 AND symb_decoder(16#dc#)) OR
 					(reg_q1997 AND symb_decoder(16#23#)) OR
 					(reg_q1997 AND symb_decoder(16#1f#)) OR
 					(reg_q1997 AND symb_decoder(16#80#)) OR
 					(reg_q1997 AND symb_decoder(16#be#)) OR
 					(reg_q1997 AND symb_decoder(16#ee#)) OR
 					(reg_q1997 AND symb_decoder(16#03#)) OR
 					(reg_q1997 AND symb_decoder(16#d6#)) OR
 					(reg_q1997 AND symb_decoder(16#82#)) OR
 					(reg_q1997 AND symb_decoder(16#c3#)) OR
 					(reg_q1997 AND symb_decoder(16#f2#)) OR
 					(reg_q1997 AND symb_decoder(16#f1#)) OR
 					(reg_q1997 AND symb_decoder(16#1c#)) OR
 					(reg_q1997 AND symb_decoder(16#5b#)) OR
 					(reg_q1997 AND symb_decoder(16#2d#)) OR
 					(reg_q1997 AND symb_decoder(16#ad#)) OR
 					(reg_q1997 AND symb_decoder(16#b6#)) OR
 					(reg_q1997 AND symb_decoder(16#55#)) OR
 					(reg_q1997 AND symb_decoder(16#30#)) OR
 					(reg_q1997 AND symb_decoder(16#ac#)) OR
 					(reg_q1997 AND symb_decoder(16#58#)) OR
 					(reg_q1997 AND symb_decoder(16#00#)) OR
 					(reg_q1997 AND symb_decoder(16#e0#)) OR
 					(reg_q1997 AND symb_decoder(16#52#)) OR
 					(reg_q1997 AND symb_decoder(16#77#)) OR
 					(reg_q1997 AND symb_decoder(16#66#)) OR
 					(reg_q1997 AND symb_decoder(16#7d#)) OR
 					(reg_q1997 AND symb_decoder(16#f4#)) OR
 					(reg_q1997 AND symb_decoder(16#8e#)) OR
 					(reg_q1997 AND symb_decoder(16#33#)) OR
 					(reg_q1997 AND symb_decoder(16#56#)) OR
 					(reg_q1997 AND symb_decoder(16#bf#)) OR
 					(reg_q1997 AND symb_decoder(16#3b#)) OR
 					(reg_q1997 AND symb_decoder(16#4c#)) OR
 					(reg_q1997 AND symb_decoder(16#85#)) OR
 					(reg_q1997 AND symb_decoder(16#ab#)) OR
 					(reg_q1997 AND symb_decoder(16#b1#)) OR
 					(reg_q1997 AND symb_decoder(16#de#)) OR
 					(reg_q1997 AND symb_decoder(16#8a#)) OR
 					(reg_q1997 AND symb_decoder(16#69#)) OR
 					(reg_q1997 AND symb_decoder(16#f5#)) OR
 					(reg_q1997 AND symb_decoder(16#aa#)) OR
 					(reg_q1997 AND symb_decoder(16#4f#)) OR
 					(reg_q1997 AND symb_decoder(16#41#)) OR
 					(reg_q1997 AND symb_decoder(16#c6#)) OR
 					(reg_q1997 AND symb_decoder(16#a2#)) OR
 					(reg_q1997 AND symb_decoder(16#bb#)) OR
 					(reg_q1997 AND symb_decoder(16#ed#)) OR
 					(reg_q1997 AND symb_decoder(16#7b#)) OR
 					(reg_q1997 AND symb_decoder(16#f0#)) OR
 					(reg_q1997 AND symb_decoder(16#ea#)) OR
 					(reg_q1997 AND symb_decoder(16#94#)) OR
 					(reg_q1997 AND symb_decoder(16#74#)) OR
 					(reg_q1997 AND symb_decoder(16#3d#)) OR
 					(reg_q1997 AND symb_decoder(16#78#)) OR
 					(reg_q1997 AND symb_decoder(16#a8#)) OR
 					(reg_q1997 AND symb_decoder(16#e6#)) OR
 					(reg_q1997 AND symb_decoder(16#57#)) OR
 					(reg_q1997 AND symb_decoder(16#d7#)) OR
 					(reg_q1997 AND symb_decoder(16#8d#)) OR
 					(reg_q1997 AND symb_decoder(16#70#)) OR
 					(reg_q1997 AND symb_decoder(16#e8#)) OR
 					(reg_q1997 AND symb_decoder(16#d1#)) OR
 					(reg_q1997 AND symb_decoder(16#b4#)) OR
 					(reg_q1997 AND symb_decoder(16#09#)) OR
 					(reg_q1997 AND symb_decoder(16#1b#)) OR
 					(reg_q1997 AND symb_decoder(16#cd#)) OR
 					(reg_q1997 AND symb_decoder(16#07#)) OR
 					(reg_q1997 AND symb_decoder(16#fb#)) OR
 					(reg_q1997 AND symb_decoder(16#7a#)) OR
 					(reg_q1997 AND symb_decoder(16#62#)) OR
 					(reg_q1997 AND symb_decoder(16#1e#)) OR
 					(reg_q1997 AND symb_decoder(16#3e#)) OR
 					(reg_q1997 AND symb_decoder(16#2b#)) OR
 					(reg_q1997 AND symb_decoder(16#c0#)) OR
 					(reg_q1997 AND symb_decoder(16#49#)) OR
 					(reg_q1997 AND symb_decoder(16#51#)) OR
 					(reg_q1997 AND symb_decoder(16#12#)) OR
 					(reg_q1997 AND symb_decoder(16#af#)) OR
 					(reg_q1997 AND symb_decoder(16#c7#)) OR
 					(reg_q1997 AND symb_decoder(16#a9#)) OR
 					(reg_q1997 AND symb_decoder(16#42#)) OR
 					(reg_q1997 AND symb_decoder(16#75#)) OR
 					(reg_q1997 AND symb_decoder(16#6b#)) OR
 					(reg_q1997 AND symb_decoder(16#38#)) OR
 					(reg_q1997 AND symb_decoder(16#98#)) OR
 					(reg_q1997 AND symb_decoder(16#96#)) OR
 					(reg_q1997 AND symb_decoder(16#a1#)) OR
 					(reg_q1997 AND symb_decoder(16#dd#)) OR
 					(reg_q1997 AND symb_decoder(16#1d#)) OR
 					(reg_q1997 AND symb_decoder(16#7f#)) OR
 					(reg_q1997 AND symb_decoder(16#f8#)) OR
 					(reg_q1997 AND symb_decoder(16#0f#)) OR
 					(reg_q1997 AND symb_decoder(16#c5#)) OR
 					(reg_q1997 AND symb_decoder(16#da#)) OR
 					(reg_q1997 AND symb_decoder(16#81#)) OR
 					(reg_q1997 AND symb_decoder(16#e4#)) OR
 					(reg_q1997 AND symb_decoder(16#34#)) OR
 					(reg_q1997 AND symb_decoder(16#6c#)) OR
 					(reg_q1997 AND symb_decoder(16#9d#)) OR
 					(reg_q1997 AND symb_decoder(16#5a#)) OR
 					(reg_q1997 AND symb_decoder(16#5e#)) OR
 					(reg_q1997 AND symb_decoder(16#7c#)) OR
 					(reg_q1997 AND symb_decoder(16#43#)) OR
 					(reg_q1997 AND symb_decoder(16#9a#)) OR
 					(reg_q1997 AND symb_decoder(16#46#)) OR
 					(reg_q1997 AND symb_decoder(16#06#)) OR
 					(reg_q1997 AND symb_decoder(16#6d#)) OR
 					(reg_q1997 AND symb_decoder(16#eb#)) OR
 					(reg_q1997 AND symb_decoder(16#e9#)) OR
 					(reg_q1997 AND symb_decoder(16#e1#)) OR
 					(reg_q1997 AND symb_decoder(16#61#)) OR
 					(reg_q1997 AND symb_decoder(16#c9#)) OR
 					(reg_q1997 AND symb_decoder(16#99#)) OR
 					(reg_q1975 AND symb_decoder(16#a3#)) OR
 					(reg_q1975 AND symb_decoder(16#ce#)) OR
 					(reg_q1975 AND symb_decoder(16#36#)) OR
 					(reg_q1975 AND symb_decoder(16#48#)) OR
 					(reg_q1975 AND symb_decoder(16#6a#)) OR
 					(reg_q1975 AND symb_decoder(16#53#)) OR
 					(reg_q1975 AND symb_decoder(16#0b#)) OR
 					(reg_q1975 AND symb_decoder(16#46#)) OR
 					(reg_q1975 AND symb_decoder(16#66#)) OR
 					(reg_q1975 AND symb_decoder(16#52#)) OR
 					(reg_q1975 AND symb_decoder(16#d7#)) OR
 					(reg_q1975 AND symb_decoder(16#cc#)) OR
 					(reg_q1975 AND symb_decoder(16#29#)) OR
 					(reg_q1975 AND symb_decoder(16#a0#)) OR
 					(reg_q1975 AND symb_decoder(16#12#)) OR
 					(reg_q1975 AND symb_decoder(16#b9#)) OR
 					(reg_q1975 AND symb_decoder(16#e3#)) OR
 					(reg_q1975 AND symb_decoder(16#ed#)) OR
 					(reg_q1975 AND symb_decoder(16#91#)) OR
 					(reg_q1975 AND symb_decoder(16#eb#)) OR
 					(reg_q1975 AND symb_decoder(16#f1#)) OR
 					(reg_q1975 AND symb_decoder(16#86#)) OR
 					(reg_q1975 AND symb_decoder(16#60#)) OR
 					(reg_q1975 AND symb_decoder(16#99#)) OR
 					(reg_q1975 AND symb_decoder(16#b5#)) OR
 					(reg_q1975 AND symb_decoder(16#f4#)) OR
 					(reg_q1975 AND symb_decoder(16#77#)) OR
 					(reg_q1975 AND symb_decoder(16#95#)) OR
 					(reg_q1975 AND symb_decoder(16#0e#)) OR
 					(reg_q1975 AND symb_decoder(16#96#)) OR
 					(reg_q1975 AND symb_decoder(16#ec#)) OR
 					(reg_q1975 AND symb_decoder(16#63#)) OR
 					(reg_q1975 AND symb_decoder(16#b1#)) OR
 					(reg_q1975 AND symb_decoder(16#a2#)) OR
 					(reg_q1975 AND symb_decoder(16#4e#)) OR
 					(reg_q1975 AND symb_decoder(16#20#)) OR
 					(reg_q1975 AND symb_decoder(16#f2#)) OR
 					(reg_q1975 AND symb_decoder(16#7c#)) OR
 					(reg_q1975 AND symb_decoder(16#a1#)) OR
 					(reg_q1975 AND symb_decoder(16#ca#)) OR
 					(reg_q1975 AND symb_decoder(16#fa#)) OR
 					(reg_q1975 AND symb_decoder(16#c4#)) OR
 					(reg_q1975 AND symb_decoder(16#d3#)) OR
 					(reg_q1975 AND symb_decoder(16#dd#)) OR
 					(reg_q1975 AND symb_decoder(16#10#)) OR
 					(reg_q1975 AND symb_decoder(16#fe#)) OR
 					(reg_q1975 AND symb_decoder(16#5e#)) OR
 					(reg_q1975 AND symb_decoder(16#1e#)) OR
 					(reg_q1975 AND symb_decoder(16#3d#)) OR
 					(reg_q1975 AND symb_decoder(16#28#)) OR
 					(reg_q1975 AND symb_decoder(16#15#)) OR
 					(reg_q1975 AND symb_decoder(16#38#)) OR
 					(reg_q1975 AND symb_decoder(16#82#)) OR
 					(reg_q1975 AND symb_decoder(16#75#)) OR
 					(reg_q1975 AND symb_decoder(16#d5#)) OR
 					(reg_q1975 AND symb_decoder(16#56#)) OR
 					(reg_q1975 AND symb_decoder(16#98#)) OR
 					(reg_q1975 AND symb_decoder(16#8c#)) OR
 					(reg_q1975 AND symb_decoder(16#ae#)) OR
 					(reg_q1975 AND symb_decoder(16#b7#)) OR
 					(reg_q1975 AND symb_decoder(16#ac#)) OR
 					(reg_q1975 AND symb_decoder(16#21#)) OR
 					(reg_q1975 AND symb_decoder(16#7a#)) OR
 					(reg_q1975 AND symb_decoder(16#49#)) OR
 					(reg_q1975 AND symb_decoder(16#89#)) OR
 					(reg_q1975 AND symb_decoder(16#5d#)) OR
 					(reg_q1975 AND symb_decoder(16#51#)) OR
 					(reg_q1975 AND symb_decoder(16#24#)) OR
 					(reg_q1975 AND symb_decoder(16#ad#)) OR
 					(reg_q1975 AND symb_decoder(16#67#)) OR
 					(reg_q1975 AND symb_decoder(16#81#)) OR
 					(reg_q1975 AND symb_decoder(16#64#)) OR
 					(reg_q1975 AND symb_decoder(16#79#)) OR
 					(reg_q1975 AND symb_decoder(16#90#)) OR
 					(reg_q1975 AND symb_decoder(16#cf#)) OR
 					(reg_q1975 AND symb_decoder(16#00#)) OR
 					(reg_q1975 AND symb_decoder(16#3b#)) OR
 					(reg_q1975 AND symb_decoder(16#06#)) OR
 					(reg_q1975 AND symb_decoder(16#da#)) OR
 					(reg_q1975 AND symb_decoder(16#e6#)) OR
 					(reg_q1975 AND symb_decoder(16#6d#)) OR
 					(reg_q1975 AND symb_decoder(16#25#)) OR
 					(reg_q1975 AND symb_decoder(16#3a#)) OR
 					(reg_q1975 AND symb_decoder(16#cd#)) OR
 					(reg_q1975 AND symb_decoder(16#8f#)) OR
 					(reg_q1975 AND symb_decoder(16#bb#)) OR
 					(reg_q1975 AND symb_decoder(16#6b#)) OR
 					(reg_q1975 AND symb_decoder(16#2e#)) OR
 					(reg_q1975 AND symb_decoder(16#80#)) OR
 					(reg_q1975 AND symb_decoder(16#e4#)) OR
 					(reg_q1975 AND symb_decoder(16#42#)) OR
 					(reg_q1975 AND symb_decoder(16#4f#)) OR
 					(reg_q1975 AND symb_decoder(16#ee#)) OR
 					(reg_q1975 AND symb_decoder(16#2d#)) OR
 					(reg_q1975 AND symb_decoder(16#69#)) OR
 					(reg_q1975 AND symb_decoder(16#8a#)) OR
 					(reg_q1975 AND symb_decoder(16#37#)) OR
 					(reg_q1975 AND symb_decoder(16#9d#)) OR
 					(reg_q1975 AND symb_decoder(16#9e#)) OR
 					(reg_q1975 AND symb_decoder(16#9f#)) OR
 					(reg_q1975 AND symb_decoder(16#df#)) OR
 					(reg_q1975 AND symb_decoder(16#27#)) OR
 					(reg_q1975 AND symb_decoder(16#70#)) OR
 					(reg_q1975 AND symb_decoder(16#07#)) OR
 					(reg_q1975 AND symb_decoder(16#6f#)) OR
 					(reg_q1975 AND symb_decoder(16#d0#)) OR
 					(reg_q1975 AND symb_decoder(16#e7#)) OR
 					(reg_q1975 AND symb_decoder(16#4b#)) OR
 					(reg_q1975 AND symb_decoder(16#68#)) OR
 					(reg_q1975 AND symb_decoder(16#db#)) OR
 					(reg_q1975 AND symb_decoder(16#9b#)) OR
 					(reg_q1975 AND symb_decoder(16#af#)) OR
 					(reg_q1975 AND symb_decoder(16#97#)) OR
 					(reg_q1975 AND symb_decoder(16#c7#)) OR
 					(reg_q1975 AND symb_decoder(16#8b#)) OR
 					(reg_q1975 AND symb_decoder(16#a7#)) OR
 					(reg_q1975 AND symb_decoder(16#34#)) OR
 					(reg_q1975 AND symb_decoder(16#f6#)) OR
 					(reg_q1975 AND symb_decoder(16#57#)) OR
 					(reg_q1975 AND symb_decoder(16#2f#)) OR
 					(reg_q1975 AND symb_decoder(16#fd#)) OR
 					(reg_q1975 AND symb_decoder(16#de#)) OR
 					(reg_q1975 AND symb_decoder(16#4c#)) OR
 					(reg_q1975 AND symb_decoder(16#fb#)) OR
 					(reg_q1975 AND symb_decoder(16#30#)) OR
 					(reg_q1975 AND symb_decoder(16#f8#)) OR
 					(reg_q1975 AND symb_decoder(16#19#)) OR
 					(reg_q1975 AND symb_decoder(16#7d#)) OR
 					(reg_q1975 AND symb_decoder(16#c9#)) OR
 					(reg_q1975 AND symb_decoder(16#c6#)) OR
 					(reg_q1975 AND symb_decoder(16#4d#)) OR
 					(reg_q1975 AND symb_decoder(16#b3#)) OR
 					(reg_q1975 AND symb_decoder(16#1a#)) OR
 					(reg_q1975 AND symb_decoder(16#1c#)) OR
 					(reg_q1975 AND symb_decoder(16#55#)) OR
 					(reg_q1975 AND symb_decoder(16#f5#)) OR
 					(reg_q1975 AND symb_decoder(16#bc#)) OR
 					(reg_q1975 AND symb_decoder(16#85#)) OR
 					(reg_q1975 AND symb_decoder(16#5f#)) OR
 					(reg_q1975 AND symb_decoder(16#d2#)) OR
 					(reg_q1975 AND symb_decoder(16#f0#)) OR
 					(reg_q1975 AND symb_decoder(16#c0#)) OR
 					(reg_q1975 AND symb_decoder(16#11#)) OR
 					(reg_q1975 AND symb_decoder(16#7f#)) OR
 					(reg_q1975 AND symb_decoder(16#18#)) OR
 					(reg_q1975 AND symb_decoder(16#2a#)) OR
 					(reg_q1975 AND symb_decoder(16#e2#)) OR
 					(reg_q1975 AND symb_decoder(16#1f#)) OR
 					(reg_q1975 AND symb_decoder(16#9a#)) OR
 					(reg_q1975 AND symb_decoder(16#a4#)) OR
 					(reg_q1975 AND symb_decoder(16#e0#)) OR
 					(reg_q1975 AND symb_decoder(16#5b#)) OR
 					(reg_q1975 AND symb_decoder(16#45#)) OR
 					(reg_q1975 AND symb_decoder(16#44#)) OR
 					(reg_q1975 AND symb_decoder(16#6c#)) OR
 					(reg_q1975 AND symb_decoder(16#c5#)) OR
 					(reg_q1975 AND symb_decoder(16#c1#)) OR
 					(reg_q1975 AND symb_decoder(16#8e#)) OR
 					(reg_q1975 AND symb_decoder(16#39#)) OR
 					(reg_q1975 AND symb_decoder(16#05#)) OR
 					(reg_q1975 AND symb_decoder(16#d9#)) OR
 					(reg_q1975 AND symb_decoder(16#1b#)) OR
 					(reg_q1975 AND symb_decoder(16#ea#)) OR
 					(reg_q1975 AND symb_decoder(16#bf#)) OR
 					(reg_q1975 AND symb_decoder(16#a5#)) OR
 					(reg_q1975 AND symb_decoder(16#93#)) OR
 					(reg_q1975 AND symb_decoder(16#73#)) OR
 					(reg_q1975 AND symb_decoder(16#04#)) OR
 					(reg_q1975 AND symb_decoder(16#92#)) OR
 					(reg_q1975 AND symb_decoder(16#01#)) OR
 					(reg_q1975 AND symb_decoder(16#47#)) OR
 					(reg_q1975 AND symb_decoder(16#33#)) OR
 					(reg_q1975 AND symb_decoder(16#1d#)) OR
 					(reg_q1975 AND symb_decoder(16#40#)) OR
 					(reg_q1975 AND symb_decoder(16#17#)) OR
 					(reg_q1975 AND symb_decoder(16#c8#)) OR
 					(reg_q1975 AND symb_decoder(16#4a#)) OR
 					(reg_q1975 AND symb_decoder(16#59#)) OR
 					(reg_q1975 AND symb_decoder(16#88#)) OR
 					(reg_q1975 AND symb_decoder(16#2c#)) OR
 					(reg_q1975 AND symb_decoder(16#a8#)) OR
 					(reg_q1975 AND symb_decoder(16#0c#)) OR
 					(reg_q1975 AND symb_decoder(16#08#)) OR
 					(reg_q1975 AND symb_decoder(16#b6#)) OR
 					(reg_q1975 AND symb_decoder(16#09#)) OR
 					(reg_q1975 AND symb_decoder(16#03#)) OR
 					(reg_q1975 AND symb_decoder(16#f3#)) OR
 					(reg_q1975 AND symb_decoder(16#e9#)) OR
 					(reg_q1975 AND symb_decoder(16#02#)) OR
 					(reg_q1975 AND symb_decoder(16#dc#)) OR
 					(reg_q1975 AND symb_decoder(16#c2#)) OR
 					(reg_q1975 AND symb_decoder(16#d8#)) OR
 					(reg_q1975 AND symb_decoder(16#3e#)) OR
 					(reg_q1975 AND symb_decoder(16#c3#)) OR
 					(reg_q1975 AND symb_decoder(16#23#)) OR
 					(reg_q1975 AND symb_decoder(16#35#)) OR
 					(reg_q1975 AND symb_decoder(16#83#)) OR
 					(reg_q1975 AND symb_decoder(16#41#)) OR
 					(reg_q1975 AND symb_decoder(16#58#)) OR
 					(reg_q1975 AND symb_decoder(16#3f#)) OR
 					(reg_q1975 AND symb_decoder(16#9c#)) OR
 					(reg_q1975 AND symb_decoder(16#87#)) OR
 					(reg_q1975 AND symb_decoder(16#5a#)) OR
 					(reg_q1975 AND symb_decoder(16#d1#)) OR
 					(reg_q1975 AND symb_decoder(16#32#)) OR
 					(reg_q1975 AND symb_decoder(16#62#)) OR
 					(reg_q1975 AND symb_decoder(16#61#)) OR
 					(reg_q1975 AND symb_decoder(16#6e#)) OR
 					(reg_q1975 AND symb_decoder(16#0f#)) OR
 					(reg_q1975 AND symb_decoder(16#13#)) OR
 					(reg_q1975 AND symb_decoder(16#e8#)) OR
 					(reg_q1975 AND symb_decoder(16#ab#)) OR
 					(reg_q1975 AND symb_decoder(16#43#)) OR
 					(reg_q1975 AND symb_decoder(16#72#)) OR
 					(reg_q1975 AND symb_decoder(16#a6#)) OR
 					(reg_q1975 AND symb_decoder(16#16#)) OR
 					(reg_q1975 AND symb_decoder(16#22#)) OR
 					(reg_q1975 AND symb_decoder(16#ba#)) OR
 					(reg_q1975 AND symb_decoder(16#e1#)) OR
 					(reg_q1975 AND symb_decoder(16#b2#)) OR
 					(reg_q1975 AND symb_decoder(16#aa#)) OR
 					(reg_q1975 AND symb_decoder(16#78#)) OR
 					(reg_q1975 AND symb_decoder(16#5c#)) OR
 					(reg_q1975 AND symb_decoder(16#8d#)) OR
 					(reg_q1975 AND symb_decoder(16#f7#)) OR
 					(reg_q1975 AND symb_decoder(16#76#)) OR
 					(reg_q1975 AND symb_decoder(16#cb#)) OR
 					(reg_q1975 AND symb_decoder(16#e5#)) OR
 					(reg_q1975 AND symb_decoder(16#3c#)) OR
 					(reg_q1975 AND symb_decoder(16#31#)) OR
 					(reg_q1975 AND symb_decoder(16#2b#)) OR
 					(reg_q1975 AND symb_decoder(16#b4#)) OR
 					(reg_q1975 AND symb_decoder(16#84#)) OR
 					(reg_q1975 AND symb_decoder(16#94#)) OR
 					(reg_q1975 AND symb_decoder(16#74#)) OR
 					(reg_q1975 AND symb_decoder(16#ef#)) OR
 					(reg_q1975 AND symb_decoder(16#d4#)) OR
 					(reg_q1975 AND symb_decoder(16#7b#)) OR
 					(reg_q1975 AND symb_decoder(16#d6#)) OR
 					(reg_q1975 AND symb_decoder(16#71#)) OR
 					(reg_q1975 AND symb_decoder(16#bd#)) OR
 					(reg_q1975 AND symb_decoder(16#50#)) OR
 					(reg_q1975 AND symb_decoder(16#54#)) OR
 					(reg_q1975 AND symb_decoder(16#b8#)) OR
 					(reg_q1975 AND symb_decoder(16#65#)) OR
 					(reg_q1975 AND symb_decoder(16#fc#)) OR
 					(reg_q1975 AND symb_decoder(16#26#)) OR
 					(reg_q1975 AND symb_decoder(16#b0#)) OR
 					(reg_q1975 AND symb_decoder(16#ff#)) OR
 					(reg_q1975 AND symb_decoder(16#be#)) OR
 					(reg_q1975 AND symb_decoder(16#a9#)) OR
 					(reg_q1975 AND symb_decoder(16#7e#)) OR
 					(reg_q1975 AND symb_decoder(16#14#)) OR
 					(reg_q1975 AND symb_decoder(16#f9#));
reg_q1997_init <= '0' ;
	p_reg_q1997: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1997 <= reg_q1997_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1997 <= reg_q1997_init;
        else
          reg_q1997 <= reg_q1997_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q933_in <= (reg_q931 AND symb_decoder(16#00#));
reg_q933_init <= '0' ;
	p_reg_q933: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q933 <= reg_q933_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q933 <= reg_q933_init;
        else
          reg_q933 <= reg_q933_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q955_in <= (reg_q933 AND symb_decoder(16#37#)) OR
 					(reg_q933 AND symb_decoder(16#c6#)) OR
 					(reg_q933 AND symb_decoder(16#66#)) OR
 					(reg_q933 AND symb_decoder(16#73#)) OR
 					(reg_q933 AND symb_decoder(16#7e#)) OR
 					(reg_q933 AND symb_decoder(16#b6#)) OR
 					(reg_q933 AND symb_decoder(16#d8#)) OR
 					(reg_q933 AND symb_decoder(16#7f#)) OR
 					(reg_q933 AND symb_decoder(16#e6#)) OR
 					(reg_q933 AND symb_decoder(16#7d#)) OR
 					(reg_q933 AND symb_decoder(16#63#)) OR
 					(reg_q933 AND symb_decoder(16#22#)) OR
 					(reg_q933 AND symb_decoder(16#e4#)) OR
 					(reg_q933 AND symb_decoder(16#c0#)) OR
 					(reg_q933 AND symb_decoder(16#8b#)) OR
 					(reg_q933 AND symb_decoder(16#cb#)) OR
 					(reg_q933 AND symb_decoder(16#06#)) OR
 					(reg_q933 AND symb_decoder(16#ed#)) OR
 					(reg_q933 AND symb_decoder(16#4a#)) OR
 					(reg_q933 AND symb_decoder(16#e8#)) OR
 					(reg_q933 AND symb_decoder(16#9d#)) OR
 					(reg_q933 AND symb_decoder(16#33#)) OR
 					(reg_q933 AND symb_decoder(16#a2#)) OR
 					(reg_q933 AND symb_decoder(16#db#)) OR
 					(reg_q933 AND symb_decoder(16#69#)) OR
 					(reg_q933 AND symb_decoder(16#ac#)) OR
 					(reg_q933 AND symb_decoder(16#1c#)) OR
 					(reg_q933 AND symb_decoder(16#c7#)) OR
 					(reg_q933 AND symb_decoder(16#cd#)) OR
 					(reg_q933 AND symb_decoder(16#8f#)) OR
 					(reg_q933 AND symb_decoder(16#40#)) OR
 					(reg_q933 AND symb_decoder(16#03#)) OR
 					(reg_q933 AND symb_decoder(16#f1#)) OR
 					(reg_q933 AND symb_decoder(16#68#)) OR
 					(reg_q933 AND symb_decoder(16#54#)) OR
 					(reg_q933 AND symb_decoder(16#bb#)) OR
 					(reg_q933 AND symb_decoder(16#71#)) OR
 					(reg_q933 AND symb_decoder(16#0f#)) OR
 					(reg_q933 AND symb_decoder(16#c4#)) OR
 					(reg_q933 AND symb_decoder(16#87#)) OR
 					(reg_q933 AND symb_decoder(16#8c#)) OR
 					(reg_q933 AND symb_decoder(16#9a#)) OR
 					(reg_q933 AND symb_decoder(16#f2#)) OR
 					(reg_q933 AND symb_decoder(16#b9#)) OR
 					(reg_q933 AND symb_decoder(16#90#)) OR
 					(reg_q933 AND symb_decoder(16#d9#)) OR
 					(reg_q933 AND symb_decoder(16#e3#)) OR
 					(reg_q933 AND symb_decoder(16#30#)) OR
 					(reg_q933 AND symb_decoder(16#ee#)) OR
 					(reg_q933 AND symb_decoder(16#c9#)) OR
 					(reg_q933 AND symb_decoder(16#f6#)) OR
 					(reg_q933 AND symb_decoder(16#e7#)) OR
 					(reg_q933 AND symb_decoder(16#18#)) OR
 					(reg_q933 AND symb_decoder(16#00#)) OR
 					(reg_q933 AND symb_decoder(16#a6#)) OR
 					(reg_q933 AND symb_decoder(16#39#)) OR
 					(reg_q933 AND symb_decoder(16#4f#)) OR
 					(reg_q933 AND symb_decoder(16#42#)) OR
 					(reg_q933 AND symb_decoder(16#36#)) OR
 					(reg_q933 AND symb_decoder(16#20#)) OR
 					(reg_q933 AND symb_decoder(16#4c#)) OR
 					(reg_q933 AND symb_decoder(16#a4#)) OR
 					(reg_q933 AND symb_decoder(16#15#)) OR
 					(reg_q933 AND symb_decoder(16#1a#)) OR
 					(reg_q933 AND symb_decoder(16#fc#)) OR
 					(reg_q933 AND symb_decoder(16#4e#)) OR
 					(reg_q933 AND symb_decoder(16#83#)) OR
 					(reg_q933 AND symb_decoder(16#79#)) OR
 					(reg_q933 AND symb_decoder(16#be#)) OR
 					(reg_q933 AND symb_decoder(16#d0#)) OR
 					(reg_q933 AND symb_decoder(16#c8#)) OR
 					(reg_q933 AND symb_decoder(16#24#)) OR
 					(reg_q933 AND symb_decoder(16#6d#)) OR
 					(reg_q933 AND symb_decoder(16#89#)) OR
 					(reg_q933 AND symb_decoder(16#94#)) OR
 					(reg_q933 AND symb_decoder(16#88#)) OR
 					(reg_q933 AND symb_decoder(16#5a#)) OR
 					(reg_q933 AND symb_decoder(16#bd#)) OR
 					(reg_q933 AND symb_decoder(16#ba#)) OR
 					(reg_q933 AND symb_decoder(16#ef#)) OR
 					(reg_q933 AND symb_decoder(16#51#)) OR
 					(reg_q933 AND symb_decoder(16#c2#)) OR
 					(reg_q933 AND symb_decoder(16#8e#)) OR
 					(reg_q933 AND symb_decoder(16#27#)) OR
 					(reg_q933 AND symb_decoder(16#4b#)) OR
 					(reg_q933 AND symb_decoder(16#5c#)) OR
 					(reg_q933 AND symb_decoder(16#3d#)) OR
 					(reg_q933 AND symb_decoder(16#07#)) OR
 					(reg_q933 AND symb_decoder(16#b5#)) OR
 					(reg_q933 AND symb_decoder(16#e1#)) OR
 					(reg_q933 AND symb_decoder(16#2a#)) OR
 					(reg_q933 AND symb_decoder(16#cc#)) OR
 					(reg_q933 AND symb_decoder(16#43#)) OR
 					(reg_q933 AND symb_decoder(16#19#)) OR
 					(reg_q933 AND symb_decoder(16#65#)) OR
 					(reg_q933 AND symb_decoder(16#f9#)) OR
 					(reg_q933 AND symb_decoder(16#b2#)) OR
 					(reg_q933 AND symb_decoder(16#96#)) OR
 					(reg_q933 AND symb_decoder(16#d1#)) OR
 					(reg_q933 AND symb_decoder(16#2c#)) OR
 					(reg_q933 AND symb_decoder(16#dd#)) OR
 					(reg_q933 AND symb_decoder(16#7b#)) OR
 					(reg_q933 AND symb_decoder(16#76#)) OR
 					(reg_q933 AND symb_decoder(16#9e#)) OR
 					(reg_q933 AND symb_decoder(16#84#)) OR
 					(reg_q933 AND symb_decoder(16#df#)) OR
 					(reg_q933 AND symb_decoder(16#78#)) OR
 					(reg_q933 AND symb_decoder(16#a8#)) OR
 					(reg_q933 AND symb_decoder(16#55#)) OR
 					(reg_q933 AND symb_decoder(16#45#)) OR
 					(reg_q933 AND symb_decoder(16#e9#)) OR
 					(reg_q933 AND symb_decoder(16#f5#)) OR
 					(reg_q933 AND symb_decoder(16#12#)) OR
 					(reg_q933 AND symb_decoder(16#bc#)) OR
 					(reg_q933 AND symb_decoder(16#48#)) OR
 					(reg_q933 AND symb_decoder(16#8a#)) OR
 					(reg_q933 AND symb_decoder(16#f8#)) OR
 					(reg_q933 AND symb_decoder(16#98#)) OR
 					(reg_q933 AND symb_decoder(16#0b#)) OR
 					(reg_q933 AND symb_decoder(16#91#)) OR
 					(reg_q933 AND symb_decoder(16#60#)) OR
 					(reg_q933 AND symb_decoder(16#80#)) OR
 					(reg_q933 AND symb_decoder(16#fb#)) OR
 					(reg_q933 AND symb_decoder(16#92#)) OR
 					(reg_q933 AND symb_decoder(16#ff#)) OR
 					(reg_q933 AND symb_decoder(16#3c#)) OR
 					(reg_q933 AND symb_decoder(16#67#)) OR
 					(reg_q933 AND symb_decoder(16#ca#)) OR
 					(reg_q933 AND symb_decoder(16#af#)) OR
 					(reg_q933 AND symb_decoder(16#52#)) OR
 					(reg_q933 AND symb_decoder(16#d7#)) OR
 					(reg_q933 AND symb_decoder(16#ad#)) OR
 					(reg_q933 AND symb_decoder(16#17#)) OR
 					(reg_q933 AND symb_decoder(16#9f#)) OR
 					(reg_q933 AND symb_decoder(16#97#)) OR
 					(reg_q933 AND symb_decoder(16#f3#)) OR
 					(reg_q933 AND symb_decoder(16#ec#)) OR
 					(reg_q933 AND symb_decoder(16#02#)) OR
 					(reg_q933 AND symb_decoder(16#2e#)) OR
 					(reg_q933 AND symb_decoder(16#11#)) OR
 					(reg_q933 AND symb_decoder(16#a3#)) OR
 					(reg_q933 AND symb_decoder(16#6e#)) OR
 					(reg_q933 AND symb_decoder(16#de#)) OR
 					(reg_q933 AND symb_decoder(16#b7#)) OR
 					(reg_q933 AND symb_decoder(16#d6#)) OR
 					(reg_q933 AND symb_decoder(16#7a#)) OR
 					(reg_q933 AND symb_decoder(16#46#)) OR
 					(reg_q933 AND symb_decoder(16#e2#)) OR
 					(reg_q933 AND symb_decoder(16#f7#)) OR
 					(reg_q933 AND symb_decoder(16#95#)) OR
 					(reg_q933 AND symb_decoder(16#fd#)) OR
 					(reg_q933 AND symb_decoder(16#56#)) OR
 					(reg_q933 AND symb_decoder(16#fa#)) OR
 					(reg_q933 AND symb_decoder(16#28#)) OR
 					(reg_q933 AND symb_decoder(16#3f#)) OR
 					(reg_q933 AND symb_decoder(16#2f#)) OR
 					(reg_q933 AND symb_decoder(16#29#)) OR
 					(reg_q933 AND symb_decoder(16#72#)) OR
 					(reg_q933 AND symb_decoder(16#bf#)) OR
 					(reg_q933 AND symb_decoder(16#85#)) OR
 					(reg_q933 AND symb_decoder(16#26#)) OR
 					(reg_q933 AND symb_decoder(16#59#)) OR
 					(reg_q933 AND symb_decoder(16#53#)) OR
 					(reg_q933 AND symb_decoder(16#75#)) OR
 					(reg_q933 AND symb_decoder(16#58#)) OR
 					(reg_q933 AND symb_decoder(16#34#)) OR
 					(reg_q933 AND symb_decoder(16#04#)) OR
 					(reg_q933 AND symb_decoder(16#05#)) OR
 					(reg_q933 AND symb_decoder(16#7c#)) OR
 					(reg_q933 AND symb_decoder(16#44#)) OR
 					(reg_q933 AND symb_decoder(16#1f#)) OR
 					(reg_q933 AND symb_decoder(16#6c#)) OR
 					(reg_q933 AND symb_decoder(16#2b#)) OR
 					(reg_q933 AND symb_decoder(16#2d#)) OR
 					(reg_q933 AND symb_decoder(16#6f#)) OR
 					(reg_q933 AND symb_decoder(16#1e#)) OR
 					(reg_q933 AND symb_decoder(16#d4#)) OR
 					(reg_q933 AND symb_decoder(16#f4#)) OR
 					(reg_q933 AND symb_decoder(16#01#)) OR
 					(reg_q933 AND symb_decoder(16#9c#)) OR
 					(reg_q933 AND symb_decoder(16#d3#)) OR
 					(reg_q933 AND symb_decoder(16#62#)) OR
 					(reg_q933 AND symb_decoder(16#eb#)) OR
 					(reg_q933 AND symb_decoder(16#82#)) OR
 					(reg_q933 AND symb_decoder(16#86#)) OR
 					(reg_q933 AND symb_decoder(16#74#)) OR
 					(reg_q933 AND symb_decoder(16#08#)) OR
 					(reg_q933 AND symb_decoder(16#b8#)) OR
 					(reg_q933 AND symb_decoder(16#dc#)) OR
 					(reg_q933 AND symb_decoder(16#c1#)) OR
 					(reg_q933 AND symb_decoder(16#35#)) OR
 					(reg_q933 AND symb_decoder(16#47#)) OR
 					(reg_q933 AND symb_decoder(16#14#)) OR
 					(reg_q933 AND symb_decoder(16#ab#)) OR
 					(reg_q933 AND symb_decoder(16#6a#)) OR
 					(reg_q933 AND symb_decoder(16#c3#)) OR
 					(reg_q933 AND symb_decoder(16#99#)) OR
 					(reg_q933 AND symb_decoder(16#5b#)) OR
 					(reg_q933 AND symb_decoder(16#3e#)) OR
 					(reg_q933 AND symb_decoder(16#0c#)) OR
 					(reg_q933 AND symb_decoder(16#b4#)) OR
 					(reg_q933 AND symb_decoder(16#09#)) OR
 					(reg_q933 AND symb_decoder(16#32#)) OR
 					(reg_q933 AND symb_decoder(16#4d#)) OR
 					(reg_q933 AND symb_decoder(16#cf#)) OR
 					(reg_q933 AND symb_decoder(16#a7#)) OR
 					(reg_q933 AND symb_decoder(16#0e#)) OR
 					(reg_q933 AND symb_decoder(16#31#)) OR
 					(reg_q933 AND symb_decoder(16#64#)) OR
 					(reg_q933 AND symb_decoder(16#13#)) OR
 					(reg_q933 AND symb_decoder(16#61#)) OR
 					(reg_q933 AND symb_decoder(16#70#)) OR
 					(reg_q933 AND symb_decoder(16#16#)) OR
 					(reg_q933 AND symb_decoder(16#21#)) OR
 					(reg_q933 AND symb_decoder(16#5e#)) OR
 					(reg_q933 AND symb_decoder(16#49#)) OR
 					(reg_q933 AND symb_decoder(16#b3#)) OR
 					(reg_q933 AND symb_decoder(16#23#)) OR
 					(reg_q933 AND symb_decoder(16#a9#)) OR
 					(reg_q933 AND symb_decoder(16#e5#)) OR
 					(reg_q933 AND symb_decoder(16#1d#)) OR
 					(reg_q933 AND symb_decoder(16#da#)) OR
 					(reg_q933 AND symb_decoder(16#a5#)) OR
 					(reg_q933 AND symb_decoder(16#9b#)) OR
 					(reg_q933 AND symb_decoder(16#a0#)) OR
 					(reg_q933 AND symb_decoder(16#5d#)) OR
 					(reg_q933 AND symb_decoder(16#77#)) OR
 					(reg_q933 AND symb_decoder(16#d2#)) OR
 					(reg_q933 AND symb_decoder(16#10#)) OR
 					(reg_q933 AND symb_decoder(16#f0#)) OR
 					(reg_q933 AND symb_decoder(16#ea#)) OR
 					(reg_q933 AND symb_decoder(16#d5#)) OR
 					(reg_q933 AND symb_decoder(16#50#)) OR
 					(reg_q933 AND symb_decoder(16#3a#)) OR
 					(reg_q933 AND symb_decoder(16#38#)) OR
 					(reg_q933 AND symb_decoder(16#b0#)) OR
 					(reg_q933 AND symb_decoder(16#fe#)) OR
 					(reg_q933 AND symb_decoder(16#3b#)) OR
 					(reg_q933 AND symb_decoder(16#c5#)) OR
 					(reg_q933 AND symb_decoder(16#a1#)) OR
 					(reg_q933 AND symb_decoder(16#aa#)) OR
 					(reg_q933 AND symb_decoder(16#e0#)) OR
 					(reg_q933 AND symb_decoder(16#93#)) OR
 					(reg_q933 AND symb_decoder(16#ce#)) OR
 					(reg_q933 AND symb_decoder(16#1b#)) OR
 					(reg_q933 AND symb_decoder(16#6b#)) OR
 					(reg_q933 AND symb_decoder(16#41#)) OR
 					(reg_q933 AND symb_decoder(16#57#)) OR
 					(reg_q933 AND symb_decoder(16#81#)) OR
 					(reg_q933 AND symb_decoder(16#8d#)) OR
 					(reg_q933 AND symb_decoder(16#ae#)) OR
 					(reg_q933 AND symb_decoder(16#25#)) OR
 					(reg_q933 AND symb_decoder(16#5f#)) OR
 					(reg_q933 AND symb_decoder(16#b1#)) OR
 					(reg_q955 AND symb_decoder(16#08#)) OR
 					(reg_q955 AND symb_decoder(16#52#)) OR
 					(reg_q955 AND symb_decoder(16#67#)) OR
 					(reg_q955 AND symb_decoder(16#4c#)) OR
 					(reg_q955 AND symb_decoder(16#40#)) OR
 					(reg_q955 AND symb_decoder(16#ee#)) OR
 					(reg_q955 AND symb_decoder(16#2f#)) OR
 					(reg_q955 AND symb_decoder(16#7b#)) OR
 					(reg_q955 AND symb_decoder(16#cf#)) OR
 					(reg_q955 AND symb_decoder(16#de#)) OR
 					(reg_q955 AND symb_decoder(16#8b#)) OR
 					(reg_q955 AND symb_decoder(16#c3#)) OR
 					(reg_q955 AND symb_decoder(16#e5#)) OR
 					(reg_q955 AND symb_decoder(16#b6#)) OR
 					(reg_q955 AND symb_decoder(16#05#)) OR
 					(reg_q955 AND symb_decoder(16#18#)) OR
 					(reg_q955 AND symb_decoder(16#15#)) OR
 					(reg_q955 AND symb_decoder(16#17#)) OR
 					(reg_q955 AND symb_decoder(16#1a#)) OR
 					(reg_q955 AND symb_decoder(16#01#)) OR
 					(reg_q955 AND symb_decoder(16#1f#)) OR
 					(reg_q955 AND symb_decoder(16#00#)) OR
 					(reg_q955 AND symb_decoder(16#ba#)) OR
 					(reg_q955 AND symb_decoder(16#df#)) OR
 					(reg_q955 AND symb_decoder(16#36#)) OR
 					(reg_q955 AND symb_decoder(16#84#)) OR
 					(reg_q955 AND symb_decoder(16#f3#)) OR
 					(reg_q955 AND symb_decoder(16#a5#)) OR
 					(reg_q955 AND symb_decoder(16#1d#)) OR
 					(reg_q955 AND symb_decoder(16#f1#)) OR
 					(reg_q955 AND symb_decoder(16#3b#)) OR
 					(reg_q955 AND symb_decoder(16#b3#)) OR
 					(reg_q955 AND symb_decoder(16#f2#)) OR
 					(reg_q955 AND symb_decoder(16#20#)) OR
 					(reg_q955 AND symb_decoder(16#be#)) OR
 					(reg_q955 AND symb_decoder(16#d4#)) OR
 					(reg_q955 AND symb_decoder(16#3c#)) OR
 					(reg_q955 AND symb_decoder(16#dc#)) OR
 					(reg_q955 AND symb_decoder(16#9d#)) OR
 					(reg_q955 AND symb_decoder(16#44#)) OR
 					(reg_q955 AND symb_decoder(16#e8#)) OR
 					(reg_q955 AND symb_decoder(16#46#)) OR
 					(reg_q955 AND symb_decoder(16#80#)) OR
 					(reg_q955 AND symb_decoder(16#9c#)) OR
 					(reg_q955 AND symb_decoder(16#9e#)) OR
 					(reg_q955 AND symb_decoder(16#c6#)) OR
 					(reg_q955 AND symb_decoder(16#64#)) OR
 					(reg_q955 AND symb_decoder(16#b1#)) OR
 					(reg_q955 AND symb_decoder(16#9a#)) OR
 					(reg_q955 AND symb_decoder(16#11#)) OR
 					(reg_q955 AND symb_decoder(16#7a#)) OR
 					(reg_q955 AND symb_decoder(16#57#)) OR
 					(reg_q955 AND symb_decoder(16#ed#)) OR
 					(reg_q955 AND symb_decoder(16#1e#)) OR
 					(reg_q955 AND symb_decoder(16#fa#)) OR
 					(reg_q955 AND symb_decoder(16#dd#)) OR
 					(reg_q955 AND symb_decoder(16#94#)) OR
 					(reg_q955 AND symb_decoder(16#a4#)) OR
 					(reg_q955 AND symb_decoder(16#af#)) OR
 					(reg_q955 AND symb_decoder(16#6d#)) OR
 					(reg_q955 AND symb_decoder(16#63#)) OR
 					(reg_q955 AND symb_decoder(16#47#)) OR
 					(reg_q955 AND symb_decoder(16#76#)) OR
 					(reg_q955 AND symb_decoder(16#6b#)) OR
 					(reg_q955 AND symb_decoder(16#70#)) OR
 					(reg_q955 AND symb_decoder(16#ad#)) OR
 					(reg_q955 AND symb_decoder(16#b8#)) OR
 					(reg_q955 AND symb_decoder(16#4f#)) OR
 					(reg_q955 AND symb_decoder(16#e2#)) OR
 					(reg_q955 AND symb_decoder(16#a7#)) OR
 					(reg_q955 AND symb_decoder(16#06#)) OR
 					(reg_q955 AND symb_decoder(16#81#)) OR
 					(reg_q955 AND symb_decoder(16#cd#)) OR
 					(reg_q955 AND symb_decoder(16#ae#)) OR
 					(reg_q955 AND symb_decoder(16#8e#)) OR
 					(reg_q955 AND symb_decoder(16#31#)) OR
 					(reg_q955 AND symb_decoder(16#bd#)) OR
 					(reg_q955 AND symb_decoder(16#69#)) OR
 					(reg_q955 AND symb_decoder(16#32#)) OR
 					(reg_q955 AND symb_decoder(16#9b#)) OR
 					(reg_q955 AND symb_decoder(16#16#)) OR
 					(reg_q955 AND symb_decoder(16#30#)) OR
 					(reg_q955 AND symb_decoder(16#49#)) OR
 					(reg_q955 AND symb_decoder(16#eb#)) OR
 					(reg_q955 AND symb_decoder(16#82#)) OR
 					(reg_q955 AND symb_decoder(16#97#)) OR
 					(reg_q955 AND symb_decoder(16#98#)) OR
 					(reg_q955 AND symb_decoder(16#f5#)) OR
 					(reg_q955 AND symb_decoder(16#72#)) OR
 					(reg_q955 AND symb_decoder(16#19#)) OR
 					(reg_q955 AND symb_decoder(16#58#)) OR
 					(reg_q955 AND symb_decoder(16#99#)) OR
 					(reg_q955 AND symb_decoder(16#1b#)) OR
 					(reg_q955 AND symb_decoder(16#41#)) OR
 					(reg_q955 AND symb_decoder(16#53#)) OR
 					(reg_q955 AND symb_decoder(16#34#)) OR
 					(reg_q955 AND symb_decoder(16#ea#)) OR
 					(reg_q955 AND symb_decoder(16#3e#)) OR
 					(reg_q955 AND symb_decoder(16#f0#)) OR
 					(reg_q955 AND symb_decoder(16#6f#)) OR
 					(reg_q955 AND symb_decoder(16#e1#)) OR
 					(reg_q955 AND symb_decoder(16#d6#)) OR
 					(reg_q955 AND symb_decoder(16#78#)) OR
 					(reg_q955 AND symb_decoder(16#56#)) OR
 					(reg_q955 AND symb_decoder(16#03#)) OR
 					(reg_q955 AND symb_decoder(16#2a#)) OR
 					(reg_q955 AND symb_decoder(16#4b#)) OR
 					(reg_q955 AND symb_decoder(16#3d#)) OR
 					(reg_q955 AND symb_decoder(16#61#)) OR
 					(reg_q955 AND symb_decoder(16#cb#)) OR
 					(reg_q955 AND symb_decoder(16#b4#)) OR
 					(reg_q955 AND symb_decoder(16#48#)) OR
 					(reg_q955 AND symb_decoder(16#86#)) OR
 					(reg_q955 AND symb_decoder(16#c8#)) OR
 					(reg_q955 AND symb_decoder(16#74#)) OR
 					(reg_q955 AND symb_decoder(16#a8#)) OR
 					(reg_q955 AND symb_decoder(16#7d#)) OR
 					(reg_q955 AND symb_decoder(16#79#)) OR
 					(reg_q955 AND symb_decoder(16#e6#)) OR
 					(reg_q955 AND symb_decoder(16#0f#)) OR
 					(reg_q955 AND symb_decoder(16#e9#)) OR
 					(reg_q955 AND symb_decoder(16#59#)) OR
 					(reg_q955 AND symb_decoder(16#25#)) OR
 					(reg_q955 AND symb_decoder(16#5d#)) OR
 					(reg_q955 AND symb_decoder(16#35#)) OR
 					(reg_q955 AND symb_decoder(16#50#)) OR
 					(reg_q955 AND symb_decoder(16#22#)) OR
 					(reg_q955 AND symb_decoder(16#87#)) OR
 					(reg_q955 AND symb_decoder(16#d7#)) OR
 					(reg_q955 AND symb_decoder(16#3a#)) OR
 					(reg_q955 AND symb_decoder(16#42#)) OR
 					(reg_q955 AND symb_decoder(16#c9#)) OR
 					(reg_q955 AND symb_decoder(16#b5#)) OR
 					(reg_q955 AND symb_decoder(16#10#)) OR
 					(reg_q955 AND symb_decoder(16#d9#)) OR
 					(reg_q955 AND symb_decoder(16#13#)) OR
 					(reg_q955 AND symb_decoder(16#71#)) OR
 					(reg_q955 AND symb_decoder(16#33#)) OR
 					(reg_q955 AND symb_decoder(16#4d#)) OR
 					(reg_q955 AND symb_decoder(16#e7#)) OR
 					(reg_q955 AND symb_decoder(16#ce#)) OR
 					(reg_q955 AND symb_decoder(16#c1#)) OR
 					(reg_q955 AND symb_decoder(16#93#)) OR
 					(reg_q955 AND symb_decoder(16#91#)) OR
 					(reg_q955 AND symb_decoder(16#29#)) OR
 					(reg_q955 AND symb_decoder(16#bb#)) OR
 					(reg_q955 AND symb_decoder(16#0e#)) OR
 					(reg_q955 AND symb_decoder(16#fe#)) OR
 					(reg_q955 AND symb_decoder(16#a6#)) OR
 					(reg_q955 AND symb_decoder(16#c0#)) OR
 					(reg_q955 AND symb_decoder(16#75#)) OR
 					(reg_q955 AND symb_decoder(16#37#)) OR
 					(reg_q955 AND symb_decoder(16#5c#)) OR
 					(reg_q955 AND symb_decoder(16#6c#)) OR
 					(reg_q955 AND symb_decoder(16#39#)) OR
 					(reg_q955 AND symb_decoder(16#66#)) OR
 					(reg_q955 AND symb_decoder(16#09#)) OR
 					(reg_q955 AND symb_decoder(16#c2#)) OR
 					(reg_q955 AND symb_decoder(16#8d#)) OR
 					(reg_q955 AND symb_decoder(16#4a#)) OR
 					(reg_q955 AND symb_decoder(16#b9#)) OR
 					(reg_q955 AND symb_decoder(16#24#)) OR
 					(reg_q955 AND symb_decoder(16#3f#)) OR
 					(reg_q955 AND symb_decoder(16#85#)) OR
 					(reg_q955 AND symb_decoder(16#0c#)) OR
 					(reg_q955 AND symb_decoder(16#1c#)) OR
 					(reg_q955 AND symb_decoder(16#65#)) OR
 					(reg_q955 AND symb_decoder(16#60#)) OR
 					(reg_q955 AND symb_decoder(16#6e#)) OR
 					(reg_q955 AND symb_decoder(16#8a#)) OR
 					(reg_q955 AND symb_decoder(16#6a#)) OR
 					(reg_q955 AND symb_decoder(16#90#)) OR
 					(reg_q955 AND symb_decoder(16#68#)) OR
 					(reg_q955 AND symb_decoder(16#7e#)) OR
 					(reg_q955 AND symb_decoder(16#2c#)) OR
 					(reg_q955 AND symb_decoder(16#4e#)) OR
 					(reg_q955 AND symb_decoder(16#5a#)) OR
 					(reg_q955 AND symb_decoder(16#f6#)) OR
 					(reg_q955 AND symb_decoder(16#ac#)) OR
 					(reg_q955 AND symb_decoder(16#02#)) OR
 					(reg_q955 AND symb_decoder(16#5f#)) OR
 					(reg_q955 AND symb_decoder(16#92#)) OR
 					(reg_q955 AND symb_decoder(16#89#)) OR
 					(reg_q955 AND symb_decoder(16#2b#)) OR
 					(reg_q955 AND symb_decoder(16#ef#)) OR
 					(reg_q955 AND symb_decoder(16#5b#)) OR
 					(reg_q955 AND symb_decoder(16#f4#)) OR
 					(reg_q955 AND symb_decoder(16#f7#)) OR
 					(reg_q955 AND symb_decoder(16#bf#)) OR
 					(reg_q955 AND symb_decoder(16#c4#)) OR
 					(reg_q955 AND symb_decoder(16#a0#)) OR
 					(reg_q955 AND symb_decoder(16#a9#)) OR
 					(reg_q955 AND symb_decoder(16#45#)) OR
 					(reg_q955 AND symb_decoder(16#c7#)) OR
 					(reg_q955 AND symb_decoder(16#95#)) OR
 					(reg_q955 AND symb_decoder(16#96#)) OR
 					(reg_q955 AND symb_decoder(16#12#)) OR
 					(reg_q955 AND symb_decoder(16#55#)) OR
 					(reg_q955 AND symb_decoder(16#d2#)) OR
 					(reg_q955 AND symb_decoder(16#8c#)) OR
 					(reg_q955 AND symb_decoder(16#fb#)) OR
 					(reg_q955 AND symb_decoder(16#7f#)) OR
 					(reg_q955 AND symb_decoder(16#28#)) OR
 					(reg_q955 AND symb_decoder(16#a1#)) OR
 					(reg_q955 AND symb_decoder(16#f9#)) OR
 					(reg_q955 AND symb_decoder(16#e3#)) OR
 					(reg_q955 AND symb_decoder(16#b2#)) OR
 					(reg_q955 AND symb_decoder(16#d1#)) OR
 					(reg_q955 AND symb_decoder(16#26#)) OR
 					(reg_q955 AND symb_decoder(16#51#)) OR
 					(reg_q955 AND symb_decoder(16#23#)) OR
 					(reg_q955 AND symb_decoder(16#c5#)) OR
 					(reg_q955 AND symb_decoder(16#ab#)) OR
 					(reg_q955 AND symb_decoder(16#a2#)) OR
 					(reg_q955 AND symb_decoder(16#ff#)) OR
 					(reg_q955 AND symb_decoder(16#0b#)) OR
 					(reg_q955 AND symb_decoder(16#73#)) OR
 					(reg_q955 AND symb_decoder(16#d5#)) OR
 					(reg_q955 AND symb_decoder(16#62#)) OR
 					(reg_q955 AND symb_decoder(16#aa#)) OR
 					(reg_q955 AND symb_decoder(16#9f#)) OR
 					(reg_q955 AND symb_decoder(16#f8#)) OR
 					(reg_q955 AND symb_decoder(16#db#)) OR
 					(reg_q955 AND symb_decoder(16#da#)) OR
 					(reg_q955 AND symb_decoder(16#2d#)) OR
 					(reg_q955 AND symb_decoder(16#07#)) OR
 					(reg_q955 AND symb_decoder(16#fd#)) OR
 					(reg_q955 AND symb_decoder(16#43#)) OR
 					(reg_q955 AND symb_decoder(16#bc#)) OR
 					(reg_q955 AND symb_decoder(16#e4#)) OR
 					(reg_q955 AND symb_decoder(16#04#)) OR
 					(reg_q955 AND symb_decoder(16#d3#)) OR
 					(reg_q955 AND symb_decoder(16#fc#)) OR
 					(reg_q955 AND symb_decoder(16#83#)) OR
 					(reg_q955 AND symb_decoder(16#38#)) OR
 					(reg_q955 AND symb_decoder(16#e0#)) OR
 					(reg_q955 AND symb_decoder(16#54#)) OR
 					(reg_q955 AND symb_decoder(16#ec#)) OR
 					(reg_q955 AND symb_decoder(16#7c#)) OR
 					(reg_q955 AND symb_decoder(16#14#)) OR
 					(reg_q955 AND symb_decoder(16#21#)) OR
 					(reg_q955 AND symb_decoder(16#27#)) OR
 					(reg_q955 AND symb_decoder(16#77#)) OR
 					(reg_q955 AND symb_decoder(16#5e#)) OR
 					(reg_q955 AND symb_decoder(16#b0#)) OR
 					(reg_q955 AND symb_decoder(16#b7#)) OR
 					(reg_q955 AND symb_decoder(16#2e#)) OR
 					(reg_q955 AND symb_decoder(16#88#)) OR
 					(reg_q955 AND symb_decoder(16#d8#)) OR
 					(reg_q955 AND symb_decoder(16#8f#)) OR
 					(reg_q955 AND symb_decoder(16#d0#)) OR
 					(reg_q955 AND symb_decoder(16#a3#)) OR
 					(reg_q955 AND symb_decoder(16#cc#)) OR
 					(reg_q955 AND symb_decoder(16#ca#));
reg_q955_init <= '0' ;
	p_reg_q955: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q955 <= reg_q955_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q955 <= reg_q955_init;
        else
          reg_q955 <= reg_q955_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2091_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2091 AND symb_decoder(16#33#)) OR
 					(reg_q2091 AND symb_decoder(16#3a#)) OR
 					(reg_q2091 AND symb_decoder(16#7a#)) OR
 					(reg_q2091 AND symb_decoder(16#be#)) OR
 					(reg_q2091 AND symb_decoder(16#62#)) OR
 					(reg_q2091 AND symb_decoder(16#43#)) OR
 					(reg_q2091 AND symb_decoder(16#cd#)) OR
 					(reg_q2091 AND symb_decoder(16#10#)) OR
 					(reg_q2091 AND symb_decoder(16#29#)) OR
 					(reg_q2091 AND symb_decoder(16#85#)) OR
 					(reg_q2091 AND symb_decoder(16#db#)) OR
 					(reg_q2091 AND symb_decoder(16#0e#)) OR
 					(reg_q2091 AND symb_decoder(16#46#)) OR
 					(reg_q2091 AND symb_decoder(16#ac#)) OR
 					(reg_q2091 AND symb_decoder(16#56#)) OR
 					(reg_q2091 AND symb_decoder(16#ef#)) OR
 					(reg_q2091 AND symb_decoder(16#9b#)) OR
 					(reg_q2091 AND symb_decoder(16#50#)) OR
 					(reg_q2091 AND symb_decoder(16#91#)) OR
 					(reg_q2091 AND symb_decoder(16#2e#)) OR
 					(reg_q2091 AND symb_decoder(16#13#)) OR
 					(reg_q2091 AND symb_decoder(16#da#)) OR
 					(reg_q2091 AND symb_decoder(16#d5#)) OR
 					(reg_q2091 AND symb_decoder(16#4c#)) OR
 					(reg_q2091 AND symb_decoder(16#ab#)) OR
 					(reg_q2091 AND symb_decoder(16#0a#)) OR
 					(reg_q2091 AND symb_decoder(16#5c#)) OR
 					(reg_q2091 AND symb_decoder(16#1d#)) OR
 					(reg_q2091 AND symb_decoder(16#dc#)) OR
 					(reg_q2091 AND symb_decoder(16#5e#)) OR
 					(reg_q2091 AND symb_decoder(16#84#)) OR
 					(reg_q2091 AND symb_decoder(16#fe#)) OR
 					(reg_q2091 AND symb_decoder(16#4d#)) OR
 					(reg_q2091 AND symb_decoder(16#24#)) OR
 					(reg_q2091 AND symb_decoder(16#73#)) OR
 					(reg_q2091 AND symb_decoder(16#8c#)) OR
 					(reg_q2091 AND symb_decoder(16#60#)) OR
 					(reg_q2091 AND symb_decoder(16#c8#)) OR
 					(reg_q2091 AND symb_decoder(16#3f#)) OR
 					(reg_q2091 AND symb_decoder(16#19#)) OR
 					(reg_q2091 AND symb_decoder(16#44#)) OR
 					(reg_q2091 AND symb_decoder(16#12#)) OR
 					(reg_q2091 AND symb_decoder(16#bd#)) OR
 					(reg_q2091 AND symb_decoder(16#c4#)) OR
 					(reg_q2091 AND symb_decoder(16#31#)) OR
 					(reg_q2091 AND symb_decoder(16#0b#)) OR
 					(reg_q2091 AND symb_decoder(16#d0#)) OR
 					(reg_q2091 AND symb_decoder(16#ca#)) OR
 					(reg_q2091 AND symb_decoder(16#58#)) OR
 					(reg_q2091 AND symb_decoder(16#9d#)) OR
 					(reg_q2091 AND symb_decoder(16#d6#)) OR
 					(reg_q2091 AND symb_decoder(16#86#)) OR
 					(reg_q2091 AND symb_decoder(16#d8#)) OR
 					(reg_q2091 AND symb_decoder(16#8b#)) OR
 					(reg_q2091 AND symb_decoder(16#cc#)) OR
 					(reg_q2091 AND symb_decoder(16#38#)) OR
 					(reg_q2091 AND symb_decoder(16#68#)) OR
 					(reg_q2091 AND symb_decoder(16#bf#)) OR
 					(reg_q2091 AND symb_decoder(16#2f#)) OR
 					(reg_q2091 AND symb_decoder(16#d2#)) OR
 					(reg_q2091 AND symb_decoder(16#98#)) OR
 					(reg_q2091 AND symb_decoder(16#3e#)) OR
 					(reg_q2091 AND symb_decoder(16#e2#)) OR
 					(reg_q2091 AND symb_decoder(16#40#)) OR
 					(reg_q2091 AND symb_decoder(16#ec#)) OR
 					(reg_q2091 AND symb_decoder(16#b0#)) OR
 					(reg_q2091 AND symb_decoder(16#d4#)) OR
 					(reg_q2091 AND symb_decoder(16#b8#)) OR
 					(reg_q2091 AND symb_decoder(16#5a#)) OR
 					(reg_q2091 AND symb_decoder(16#c5#)) OR
 					(reg_q2091 AND symb_decoder(16#b6#)) OR
 					(reg_q2091 AND symb_decoder(16#f2#)) OR
 					(reg_q2091 AND symb_decoder(16#55#)) OR
 					(reg_q2091 AND symb_decoder(16#54#)) OR
 					(reg_q2091 AND symb_decoder(16#08#)) OR
 					(reg_q2091 AND symb_decoder(16#c7#)) OR
 					(reg_q2091 AND symb_decoder(16#a9#)) OR
 					(reg_q2091 AND symb_decoder(16#ba#)) OR
 					(reg_q2091 AND symb_decoder(16#48#)) OR
 					(reg_q2091 AND symb_decoder(16#01#)) OR
 					(reg_q2091 AND symb_decoder(16#3c#)) OR
 					(reg_q2091 AND symb_decoder(16#1f#)) OR
 					(reg_q2091 AND symb_decoder(16#1c#)) OR
 					(reg_q2091 AND symb_decoder(16#97#)) OR
 					(reg_q2091 AND symb_decoder(16#ff#)) OR
 					(reg_q2091 AND symb_decoder(16#15#)) OR
 					(reg_q2091 AND symb_decoder(16#93#)) OR
 					(reg_q2091 AND symb_decoder(16#d9#)) OR
 					(reg_q2091 AND symb_decoder(16#74#)) OR
 					(reg_q2091 AND symb_decoder(16#b2#)) OR
 					(reg_q2091 AND symb_decoder(16#f7#)) OR
 					(reg_q2091 AND symb_decoder(16#76#)) OR
 					(reg_q2091 AND symb_decoder(16#fc#)) OR
 					(reg_q2091 AND symb_decoder(16#e6#)) OR
 					(reg_q2091 AND symb_decoder(16#99#)) OR
 					(reg_q2091 AND symb_decoder(16#b9#)) OR
 					(reg_q2091 AND symb_decoder(16#9a#)) OR
 					(reg_q2091 AND symb_decoder(16#e1#)) OR
 					(reg_q2091 AND symb_decoder(16#36#)) OR
 					(reg_q2091 AND symb_decoder(16#1a#)) OR
 					(reg_q2091 AND symb_decoder(16#6c#)) OR
 					(reg_q2091 AND symb_decoder(16#e4#)) OR
 					(reg_q2091 AND symb_decoder(16#3b#)) OR
 					(reg_q2091 AND symb_decoder(16#b3#)) OR
 					(reg_q2091 AND symb_decoder(16#d3#)) OR
 					(reg_q2091 AND symb_decoder(16#7f#)) OR
 					(reg_q2091 AND symb_decoder(16#32#)) OR
 					(reg_q2091 AND symb_decoder(16#b5#)) OR
 					(reg_q2091 AND symb_decoder(16#94#)) OR
 					(reg_q2091 AND symb_decoder(16#4a#)) OR
 					(reg_q2091 AND symb_decoder(16#4e#)) OR
 					(reg_q2091 AND symb_decoder(16#82#)) OR
 					(reg_q2091 AND symb_decoder(16#72#)) OR
 					(reg_q2091 AND symb_decoder(16#30#)) OR
 					(reg_q2091 AND symb_decoder(16#6e#)) OR
 					(reg_q2091 AND symb_decoder(16#39#)) OR
 					(reg_q2091 AND symb_decoder(16#a4#)) OR
 					(reg_q2091 AND symb_decoder(16#b1#)) OR
 					(reg_q2091 AND symb_decoder(16#cb#)) OR
 					(reg_q2091 AND symb_decoder(16#14#)) OR
 					(reg_q2091 AND symb_decoder(16#96#)) OR
 					(reg_q2091 AND symb_decoder(16#e3#)) OR
 					(reg_q2091 AND symb_decoder(16#f0#)) OR
 					(reg_q2091 AND symb_decoder(16#51#)) OR
 					(reg_q2091 AND symb_decoder(16#92#)) OR
 					(reg_q2091 AND symb_decoder(16#0d#)) OR
 					(reg_q2091 AND symb_decoder(16#52#)) OR
 					(reg_q2091 AND symb_decoder(16#4f#)) OR
 					(reg_q2091 AND symb_decoder(16#fd#)) OR
 					(reg_q2091 AND symb_decoder(16#e7#)) OR
 					(reg_q2091 AND symb_decoder(16#90#)) OR
 					(reg_q2091 AND symb_decoder(16#6f#)) OR
 					(reg_q2091 AND symb_decoder(16#59#)) OR
 					(reg_q2091 AND symb_decoder(16#8d#)) OR
 					(reg_q2091 AND symb_decoder(16#71#)) OR
 					(reg_q2091 AND symb_decoder(16#25#)) OR
 					(reg_q2091 AND symb_decoder(16#34#)) OR
 					(reg_q2091 AND symb_decoder(16#53#)) OR
 					(reg_q2091 AND symb_decoder(16#f5#)) OR
 					(reg_q2091 AND symb_decoder(16#a2#)) OR
 					(reg_q2091 AND symb_decoder(16#37#)) OR
 					(reg_q2091 AND symb_decoder(16#c9#)) OR
 					(reg_q2091 AND symb_decoder(16#05#)) OR
 					(reg_q2091 AND symb_decoder(16#9f#)) OR
 					(reg_q2091 AND symb_decoder(16#2b#)) OR
 					(reg_q2091 AND symb_decoder(16#ea#)) OR
 					(reg_q2091 AND symb_decoder(16#f6#)) OR
 					(reg_q2091 AND symb_decoder(16#22#)) OR
 					(reg_q2091 AND symb_decoder(16#78#)) OR
 					(reg_q2091 AND symb_decoder(16#f8#)) OR
 					(reg_q2091 AND symb_decoder(16#47#)) OR
 					(reg_q2091 AND symb_decoder(16#07#)) OR
 					(reg_q2091 AND symb_decoder(16#a3#)) OR
 					(reg_q2091 AND symb_decoder(16#f1#)) OR
 					(reg_q2091 AND symb_decoder(16#57#)) OR
 					(reg_q2091 AND symb_decoder(16#8f#)) OR
 					(reg_q2091 AND symb_decoder(16#0c#)) OR
 					(reg_q2091 AND symb_decoder(16#16#)) OR
 					(reg_q2091 AND symb_decoder(16#dd#)) OR
 					(reg_q2091 AND symb_decoder(16#fa#)) OR
 					(reg_q2091 AND symb_decoder(16#7c#)) OR
 					(reg_q2091 AND symb_decoder(16#e8#)) OR
 					(reg_q2091 AND symb_decoder(16#4b#)) OR
 					(reg_q2091 AND symb_decoder(16#5d#)) OR
 					(reg_q2091 AND symb_decoder(16#20#)) OR
 					(reg_q2091 AND symb_decoder(16#af#)) OR
 					(reg_q2091 AND symb_decoder(16#c6#)) OR
 					(reg_q2091 AND symb_decoder(16#89#)) OR
 					(reg_q2091 AND symb_decoder(16#a6#)) OR
 					(reg_q2091 AND symb_decoder(16#e0#)) OR
 					(reg_q2091 AND symb_decoder(16#2c#)) OR
 					(reg_q2091 AND symb_decoder(16#61#)) OR
 					(reg_q2091 AND symb_decoder(16#21#)) OR
 					(reg_q2091 AND symb_decoder(16#83#)) OR
 					(reg_q2091 AND symb_decoder(16#69#)) OR
 					(reg_q2091 AND symb_decoder(16#27#)) OR
 					(reg_q2091 AND symb_decoder(16#c1#)) OR
 					(reg_q2091 AND symb_decoder(16#2a#)) OR
 					(reg_q2091 AND symb_decoder(16#5b#)) OR
 					(reg_q2091 AND symb_decoder(16#cf#)) OR
 					(reg_q2091 AND symb_decoder(16#ee#)) OR
 					(reg_q2091 AND symb_decoder(16#06#)) OR
 					(reg_q2091 AND symb_decoder(16#17#)) OR
 					(reg_q2091 AND symb_decoder(16#b4#)) OR
 					(reg_q2091 AND symb_decoder(16#02#)) OR
 					(reg_q2091 AND symb_decoder(16#87#)) OR
 					(reg_q2091 AND symb_decoder(16#0f#)) OR
 					(reg_q2091 AND symb_decoder(16#b7#)) OR
 					(reg_q2091 AND symb_decoder(16#18#)) OR
 					(reg_q2091 AND symb_decoder(16#1e#)) OR
 					(reg_q2091 AND symb_decoder(16#04#)) OR
 					(reg_q2091 AND symb_decoder(16#d1#)) OR
 					(reg_q2091 AND symb_decoder(16#f9#)) OR
 					(reg_q2091 AND symb_decoder(16#66#)) OR
 					(reg_q2091 AND symb_decoder(16#26#)) OR
 					(reg_q2091 AND symb_decoder(16#a7#)) OR
 					(reg_q2091 AND symb_decoder(16#41#)) OR
 					(reg_q2091 AND symb_decoder(16#6d#)) OR
 					(reg_q2091 AND symb_decoder(16#49#)) OR
 					(reg_q2091 AND symb_decoder(16#65#)) OR
 					(reg_q2091 AND symb_decoder(16#63#)) OR
 					(reg_q2091 AND symb_decoder(16#6b#)) OR
 					(reg_q2091 AND symb_decoder(16#77#)) OR
 					(reg_q2091 AND symb_decoder(16#80#)) OR
 					(reg_q2091 AND symb_decoder(16#fb#)) OR
 					(reg_q2091 AND symb_decoder(16#7d#)) OR
 					(reg_q2091 AND symb_decoder(16#09#)) OR
 					(reg_q2091 AND symb_decoder(16#3d#)) OR
 					(reg_q2091 AND symb_decoder(16#75#)) OR
 					(reg_q2091 AND symb_decoder(16#03#)) OR
 					(reg_q2091 AND symb_decoder(16#7e#)) OR
 					(reg_q2091 AND symb_decoder(16#8e#)) OR
 					(reg_q2091 AND symb_decoder(16#45#)) OR
 					(reg_q2091 AND symb_decoder(16#ae#)) OR
 					(reg_q2091 AND symb_decoder(16#ed#)) OR
 					(reg_q2091 AND symb_decoder(16#d7#)) OR
 					(reg_q2091 AND symb_decoder(16#64#)) OR
 					(reg_q2091 AND symb_decoder(16#aa#)) OR
 					(reg_q2091 AND symb_decoder(16#9c#)) OR
 					(reg_q2091 AND symb_decoder(16#8a#)) OR
 					(reg_q2091 AND symb_decoder(16#c2#)) OR
 					(reg_q2091 AND symb_decoder(16#f3#)) OR
 					(reg_q2091 AND symb_decoder(16#5f#)) OR
 					(reg_q2091 AND symb_decoder(16#ce#)) OR
 					(reg_q2091 AND symb_decoder(16#c3#)) OR
 					(reg_q2091 AND symb_decoder(16#2d#)) OR
 					(reg_q2091 AND symb_decoder(16#e5#)) OR
 					(reg_q2091 AND symb_decoder(16#7b#)) OR
 					(reg_q2091 AND symb_decoder(16#11#)) OR
 					(reg_q2091 AND symb_decoder(16#f4#)) OR
 					(reg_q2091 AND symb_decoder(16#67#)) OR
 					(reg_q2091 AND symb_decoder(16#bc#)) OR
 					(reg_q2091 AND symb_decoder(16#81#)) OR
 					(reg_q2091 AND symb_decoder(16#95#)) OR
 					(reg_q2091 AND symb_decoder(16#a0#)) OR
 					(reg_q2091 AND symb_decoder(16#c0#)) OR
 					(reg_q2091 AND symb_decoder(16#28#)) OR
 					(reg_q2091 AND symb_decoder(16#70#)) OR
 					(reg_q2091 AND symb_decoder(16#df#)) OR
 					(reg_q2091 AND symb_decoder(16#42#)) OR
 					(reg_q2091 AND symb_decoder(16#eb#)) OR
 					(reg_q2091 AND symb_decoder(16#00#)) OR
 					(reg_q2091 AND symb_decoder(16#a1#)) OR
 					(reg_q2091 AND symb_decoder(16#88#)) OR
 					(reg_q2091 AND symb_decoder(16#e9#)) OR
 					(reg_q2091 AND symb_decoder(16#35#)) OR
 					(reg_q2091 AND symb_decoder(16#6a#)) OR
 					(reg_q2091 AND symb_decoder(16#23#)) OR
 					(reg_q2091 AND symb_decoder(16#bb#)) OR
 					(reg_q2091 AND symb_decoder(16#79#)) OR
 					(reg_q2091 AND symb_decoder(16#a5#)) OR
 					(reg_q2091 AND symb_decoder(16#1b#)) OR
 					(reg_q2091 AND symb_decoder(16#a8#)) OR
 					(reg_q2091 AND symb_decoder(16#ad#)) OR
 					(reg_q2091 AND symb_decoder(16#de#)) OR
 					(reg_q2091 AND symb_decoder(16#9e#));
reg_q2091_init <= '0' ;
	p_reg_q2091: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2091 <= reg_q2091_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2091 <= reg_q2091_init;
        else
          reg_q2091 <= reg_q2091_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2636_in <= (reg_q2634 AND symb_decoder(16#73#)) OR
 					(reg_q2634 AND symb_decoder(16#53#));
reg_q2636_init <= '0' ;
	p_reg_q2636: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2636 <= reg_q2636_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2636 <= reg_q2636_init;
        else
          reg_q2636 <= reg_q2636_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2638_in <= (reg_q2636 AND symb_decoder(16#65#)) OR
 					(reg_q2636 AND symb_decoder(16#45#));
reg_q2638_init <= '0' ;
	p_reg_q2638: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2638 <= reg_q2638_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2638 <= reg_q2638_init;
        else
          reg_q2638 <= reg_q2638_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q606_in <= (reg_q604 AND symb_decoder(16#56#)) OR
 					(reg_q604 AND symb_decoder(16#76#));
reg_q606_init <= '0' ;
	p_reg_q606: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q606 <= reg_q606_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q606 <= reg_q606_init;
        else
          reg_q606 <= reg_q606_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q608_in <= (reg_q606 AND symb_decoder(16#36#)) OR
 					(reg_q606 AND symb_decoder(16#34#)) OR
 					(reg_q606 AND symb_decoder(16#37#)) OR
 					(reg_q606 AND symb_decoder(16#39#)) OR
 					(reg_q606 AND symb_decoder(16#30#)) OR
 					(reg_q606 AND symb_decoder(16#38#)) OR
 					(reg_q606 AND symb_decoder(16#31#)) OR
 					(reg_q606 AND symb_decoder(16#35#)) OR
 					(reg_q606 AND symb_decoder(16#32#)) OR
 					(reg_q606 AND symb_decoder(16#33#)) OR
 					(reg_q608 AND symb_decoder(16#32#)) OR
 					(reg_q608 AND symb_decoder(16#37#)) OR
 					(reg_q608 AND symb_decoder(16#33#)) OR
 					(reg_q608 AND symb_decoder(16#39#)) OR
 					(reg_q608 AND symb_decoder(16#38#)) OR
 					(reg_q608 AND symb_decoder(16#36#)) OR
 					(reg_q608 AND symb_decoder(16#30#)) OR
 					(reg_q608 AND symb_decoder(16#31#)) OR
 					(reg_q608 AND symb_decoder(16#35#)) OR
 					(reg_q608 AND symb_decoder(16#34#));
reg_q608_init <= '0' ;
	p_reg_q608: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q608 <= reg_q608_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q608 <= reg_q608_init;
        else
          reg_q608 <= reg_q608_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1355_in <= (reg_q1355 AND symb_decoder(16#0a#)) OR
 					(reg_q1355 AND symb_decoder(16#0d#)) OR
 					(reg_q1355 AND symb_decoder(16#09#)) OR
 					(reg_q1355 AND symb_decoder(16#20#)) OR
 					(reg_q1355 AND symb_decoder(16#0c#)) OR
 					(reg_q1353 AND symb_decoder(16#09#)) OR
 					(reg_q1353 AND symb_decoder(16#0d#)) OR
 					(reg_q1353 AND symb_decoder(16#0c#)) OR
 					(reg_q1353 AND symb_decoder(16#20#)) OR
 					(reg_q1353 AND symb_decoder(16#0a#));
reg_q1355_init <= '0' ;
	p_reg_q1355: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1355 <= reg_q1355_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1355 <= reg_q1355_init;
        else
          reg_q1355 <= reg_q1355_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q618_in <= (reg_q618 AND symb_decoder(16#63#)) OR
 					(reg_q618 AND symb_decoder(16#df#)) OR
 					(reg_q618 AND symb_decoder(16#c9#)) OR
 					(reg_q618 AND symb_decoder(16#dc#)) OR
 					(reg_q618 AND symb_decoder(16#2e#)) OR
 					(reg_q618 AND symb_decoder(16#79#)) OR
 					(reg_q618 AND symb_decoder(16#bc#)) OR
 					(reg_q618 AND symb_decoder(16#f3#)) OR
 					(reg_q618 AND symb_decoder(16#53#)) OR
 					(reg_q618 AND symb_decoder(16#41#)) OR
 					(reg_q618 AND symb_decoder(16#71#)) OR
 					(reg_q618 AND symb_decoder(16#24#)) OR
 					(reg_q618 AND symb_decoder(16#b7#)) OR
 					(reg_q618 AND symb_decoder(16#0b#)) OR
 					(reg_q618 AND symb_decoder(16#60#)) OR
 					(reg_q618 AND symb_decoder(16#07#)) OR
 					(reg_q618 AND symb_decoder(16#9d#)) OR
 					(reg_q618 AND symb_decoder(16#c8#)) OR
 					(reg_q618 AND symb_decoder(16#44#)) OR
 					(reg_q618 AND symb_decoder(16#ba#)) OR
 					(reg_q618 AND symb_decoder(16#54#)) OR
 					(reg_q618 AND symb_decoder(16#69#)) OR
 					(reg_q618 AND symb_decoder(16#96#)) OR
 					(reg_q618 AND symb_decoder(16#e6#)) OR
 					(reg_q618 AND symb_decoder(16#33#)) OR
 					(reg_q618 AND symb_decoder(16#31#)) OR
 					(reg_q618 AND symb_decoder(16#d9#)) OR
 					(reg_q618 AND symb_decoder(16#d6#)) OR
 					(reg_q618 AND symb_decoder(16#aa#)) OR
 					(reg_q618 AND symb_decoder(16#88#)) OR
 					(reg_q618 AND symb_decoder(16#5f#)) OR
 					(reg_q618 AND symb_decoder(16#73#)) OR
 					(reg_q618 AND symb_decoder(16#c3#)) OR
 					(reg_q618 AND symb_decoder(16#45#)) OR
 					(reg_q618 AND symb_decoder(16#9f#)) OR
 					(reg_q618 AND symb_decoder(16#1b#)) OR
 					(reg_q618 AND symb_decoder(16#9c#)) OR
 					(reg_q618 AND symb_decoder(16#80#)) OR
 					(reg_q618 AND symb_decoder(16#c0#)) OR
 					(reg_q618 AND symb_decoder(16#50#)) OR
 					(reg_q618 AND symb_decoder(16#65#)) OR
 					(reg_q618 AND symb_decoder(16#ec#)) OR
 					(reg_q618 AND symb_decoder(16#35#)) OR
 					(reg_q618 AND symb_decoder(16#ac#)) OR
 					(reg_q618 AND symb_decoder(16#6e#)) OR
 					(reg_q618 AND symb_decoder(16#02#)) OR
 					(reg_q618 AND symb_decoder(16#ca#)) OR
 					(reg_q618 AND symb_decoder(16#4d#)) OR
 					(reg_q618 AND symb_decoder(16#48#)) OR
 					(reg_q618 AND symb_decoder(16#b9#)) OR
 					(reg_q618 AND symb_decoder(16#e8#)) OR
 					(reg_q618 AND symb_decoder(16#90#)) OR
 					(reg_q618 AND symb_decoder(16#af#)) OR
 					(reg_q618 AND symb_decoder(16#f0#)) OR
 					(reg_q618 AND symb_decoder(16#32#)) OR
 					(reg_q618 AND symb_decoder(16#0f#)) OR
 					(reg_q618 AND symb_decoder(16#36#)) OR
 					(reg_q618 AND symb_decoder(16#10#)) OR
 					(reg_q618 AND symb_decoder(16#9a#)) OR
 					(reg_q618 AND symb_decoder(16#5b#)) OR
 					(reg_q618 AND symb_decoder(16#7c#)) OR
 					(reg_q618 AND symb_decoder(16#15#)) OR
 					(reg_q618 AND symb_decoder(16#f6#)) OR
 					(reg_q618 AND symb_decoder(16#6d#)) OR
 					(reg_q618 AND symb_decoder(16#2c#)) OR
 					(reg_q618 AND symb_decoder(16#5d#)) OR
 					(reg_q618 AND symb_decoder(16#b0#)) OR
 					(reg_q618 AND symb_decoder(16#be#)) OR
 					(reg_q618 AND symb_decoder(16#d0#)) OR
 					(reg_q618 AND symb_decoder(16#d1#)) OR
 					(reg_q618 AND symb_decoder(16#8f#)) OR
 					(reg_q618 AND symb_decoder(16#1d#)) OR
 					(reg_q618 AND symb_decoder(16#8e#)) OR
 					(reg_q618 AND symb_decoder(16#fc#)) OR
 					(reg_q618 AND symb_decoder(16#2d#)) OR
 					(reg_q618 AND symb_decoder(16#9e#)) OR
 					(reg_q618 AND symb_decoder(16#a7#)) OR
 					(reg_q618 AND symb_decoder(16#3e#)) OR
 					(reg_q618 AND symb_decoder(16#cb#)) OR
 					(reg_q618 AND symb_decoder(16#b6#)) OR
 					(reg_q618 AND symb_decoder(16#16#)) OR
 					(reg_q618 AND symb_decoder(16#ab#)) OR
 					(reg_q618 AND symb_decoder(16#03#)) OR
 					(reg_q618 AND symb_decoder(16#81#)) OR
 					(reg_q618 AND symb_decoder(16#cf#)) OR
 					(reg_q618 AND symb_decoder(16#f4#)) OR
 					(reg_q618 AND symb_decoder(16#bf#)) OR
 					(reg_q618 AND symb_decoder(16#8b#)) OR
 					(reg_q618 AND symb_decoder(16#87#)) OR
 					(reg_q618 AND symb_decoder(16#5a#)) OR
 					(reg_q618 AND symb_decoder(16#72#)) OR
 					(reg_q618 AND symb_decoder(16#fb#)) OR
 					(reg_q618 AND symb_decoder(16#ad#)) OR
 					(reg_q618 AND symb_decoder(16#6a#)) OR
 					(reg_q618 AND symb_decoder(16#5e#)) OR
 					(reg_q618 AND symb_decoder(16#b1#)) OR
 					(reg_q618 AND symb_decoder(16#4b#)) OR
 					(reg_q618 AND symb_decoder(16#86#)) OR
 					(reg_q618 AND symb_decoder(16#ed#)) OR
 					(reg_q618 AND symb_decoder(16#34#)) OR
 					(reg_q618 AND symb_decoder(16#89#)) OR
 					(reg_q618 AND symb_decoder(16#77#)) OR
 					(reg_q618 AND symb_decoder(16#3b#)) OR
 					(reg_q618 AND symb_decoder(16#8a#)) OR
 					(reg_q618 AND symb_decoder(16#f8#)) OR
 					(reg_q618 AND symb_decoder(16#d2#)) OR
 					(reg_q618 AND symb_decoder(16#e0#)) OR
 					(reg_q618 AND symb_decoder(16#bd#)) OR
 					(reg_q618 AND symb_decoder(16#62#)) OR
 					(reg_q618 AND symb_decoder(16#99#)) OR
 					(reg_q618 AND symb_decoder(16#2f#)) OR
 					(reg_q618 AND symb_decoder(16#fa#)) OR
 					(reg_q618 AND symb_decoder(16#1f#)) OR
 					(reg_q618 AND symb_decoder(16#bb#)) OR
 					(reg_q618 AND symb_decoder(16#12#)) OR
 					(reg_q618 AND symb_decoder(16#95#)) OR
 					(reg_q618 AND symb_decoder(16#7f#)) OR
 					(reg_q618 AND symb_decoder(16#fe#)) OR
 					(reg_q618 AND symb_decoder(16#3d#)) OR
 					(reg_q618 AND symb_decoder(16#4c#)) OR
 					(reg_q618 AND symb_decoder(16#01#)) OR
 					(reg_q618 AND symb_decoder(16#7e#)) OR
 					(reg_q618 AND symb_decoder(16#8d#)) OR
 					(reg_q618 AND symb_decoder(16#f5#)) OR
 					(reg_q618 AND symb_decoder(16#11#)) OR
 					(reg_q618 AND symb_decoder(16#1a#)) OR
 					(reg_q618 AND symb_decoder(16#47#)) OR
 					(reg_q618 AND symb_decoder(16#98#)) OR
 					(reg_q618 AND symb_decoder(16#94#)) OR
 					(reg_q618 AND symb_decoder(16#2b#)) OR
 					(reg_q618 AND symb_decoder(16#a4#)) OR
 					(reg_q618 AND symb_decoder(16#3f#)) OR
 					(reg_q618 AND symb_decoder(16#a5#)) OR
 					(reg_q618 AND symb_decoder(16#28#)) OR
 					(reg_q618 AND symb_decoder(16#75#)) OR
 					(reg_q618 AND symb_decoder(16#26#)) OR
 					(reg_q618 AND symb_decoder(16#e9#)) OR
 					(reg_q618 AND symb_decoder(16#e2#)) OR
 					(reg_q618 AND symb_decoder(16#d7#)) OR
 					(reg_q618 AND symb_decoder(16#6f#)) OR
 					(reg_q618 AND symb_decoder(16#30#)) OR
 					(reg_q618 AND symb_decoder(16#83#)) OR
 					(reg_q618 AND symb_decoder(16#08#)) OR
 					(reg_q618 AND symb_decoder(16#a9#)) OR
 					(reg_q618 AND symb_decoder(16#f1#)) OR
 					(reg_q618 AND symb_decoder(16#f2#)) OR
 					(reg_q618 AND symb_decoder(16#25#)) OR
 					(reg_q618 AND symb_decoder(16#23#)) OR
 					(reg_q618 AND symb_decoder(16#c2#)) OR
 					(reg_q618 AND symb_decoder(16#6b#)) OR
 					(reg_q618 AND symb_decoder(16#14#)) OR
 					(reg_q618 AND symb_decoder(16#db#)) OR
 					(reg_q618 AND symb_decoder(16#58#)) OR
 					(reg_q618 AND symb_decoder(16#d3#)) OR
 					(reg_q618 AND symb_decoder(16#b4#)) OR
 					(reg_q618 AND symb_decoder(16#e3#)) OR
 					(reg_q618 AND symb_decoder(16#da#)) OR
 					(reg_q618 AND symb_decoder(16#22#)) OR
 					(reg_q618 AND symb_decoder(16#27#)) OR
 					(reg_q618 AND symb_decoder(16#fd#)) OR
 					(reg_q618 AND symb_decoder(16#46#)) OR
 					(reg_q618 AND symb_decoder(16#13#)) OR
 					(reg_q618 AND symb_decoder(16#67#)) OR
 					(reg_q618 AND symb_decoder(16#e4#)) OR
 					(reg_q618 AND symb_decoder(16#40#)) OR
 					(reg_q618 AND symb_decoder(16#38#)) OR
 					(reg_q618 AND symb_decoder(16#e1#)) OR
 					(reg_q618 AND symb_decoder(16#d5#)) OR
 					(reg_q618 AND symb_decoder(16#06#)) OR
 					(reg_q618 AND symb_decoder(16#dd#)) OR
 					(reg_q618 AND symb_decoder(16#43#)) OR
 					(reg_q618 AND symb_decoder(16#4e#)) OR
 					(reg_q618 AND symb_decoder(16#d4#)) OR
 					(reg_q618 AND symb_decoder(16#7d#)) OR
 					(reg_q618 AND symb_decoder(16#7a#)) OR
 					(reg_q618 AND symb_decoder(16#55#)) OR
 					(reg_q618 AND symb_decoder(16#04#)) OR
 					(reg_q618 AND symb_decoder(16#c6#)) OR
 					(reg_q618 AND symb_decoder(16#c4#)) OR
 					(reg_q618 AND symb_decoder(16#cc#)) OR
 					(reg_q618 AND symb_decoder(16#97#)) OR
 					(reg_q618 AND symb_decoder(16#1e#)) OR
 					(reg_q618 AND symb_decoder(16#a6#)) OR
 					(reg_q618 AND symb_decoder(16#a8#)) OR
 					(reg_q618 AND symb_decoder(16#b2#)) OR
 					(reg_q618 AND symb_decoder(16#a3#)) OR
 					(reg_q618 AND symb_decoder(16#d8#)) OR
 					(reg_q618 AND symb_decoder(16#18#)) OR
 					(reg_q618 AND symb_decoder(16#51#)) OR
 					(reg_q618 AND symb_decoder(16#c1#)) OR
 					(reg_q618 AND symb_decoder(16#ae#)) OR
 					(reg_q618 AND symb_decoder(16#b8#)) OR
 					(reg_q618 AND symb_decoder(16#2a#)) OR
 					(reg_q618 AND symb_decoder(16#e5#)) OR
 					(reg_q618 AND symb_decoder(16#3a#)) OR
 					(reg_q618 AND symb_decoder(16#a1#)) OR
 					(reg_q618 AND symb_decoder(16#b5#)) OR
 					(reg_q618 AND symb_decoder(16#3c#)) OR
 					(reg_q618 AND symb_decoder(16#f9#)) OR
 					(reg_q618 AND symb_decoder(16#19#)) OR
 					(reg_q618 AND symb_decoder(16#74#)) OR
 					(reg_q618 AND symb_decoder(16#c7#)) OR
 					(reg_q618 AND symb_decoder(16#85#)) OR
 					(reg_q618 AND symb_decoder(16#ea#)) OR
 					(reg_q618 AND symb_decoder(16#68#)) OR
 					(reg_q618 AND symb_decoder(16#7b#)) OR
 					(reg_q618 AND symb_decoder(16#cd#)) OR
 					(reg_q618 AND symb_decoder(16#4f#)) OR
 					(reg_q618 AND symb_decoder(16#61#)) OR
 					(reg_q618 AND symb_decoder(16#70#)) OR
 					(reg_q618 AND symb_decoder(16#eb#)) OR
 					(reg_q618 AND symb_decoder(16#05#)) OR
 					(reg_q618 AND symb_decoder(16#b3#)) OR
 					(reg_q618 AND symb_decoder(16#1c#)) OR
 					(reg_q618 AND symb_decoder(16#0e#)) OR
 					(reg_q618 AND symb_decoder(16#00#)) OR
 					(reg_q618 AND symb_decoder(16#17#)) OR
 					(reg_q618 AND symb_decoder(16#76#)) OR
 					(reg_q618 AND symb_decoder(16#5c#)) OR
 					(reg_q618 AND symb_decoder(16#e7#)) OR
 					(reg_q618 AND symb_decoder(16#29#)) OR
 					(reg_q618 AND symb_decoder(16#9b#)) OR
 					(reg_q618 AND symb_decoder(16#39#)) OR
 					(reg_q618 AND symb_decoder(16#91#)) OR
 					(reg_q618 AND symb_decoder(16#37#)) OR
 					(reg_q618 AND symb_decoder(16#82#)) OR
 					(reg_q618 AND symb_decoder(16#66#)) OR
 					(reg_q618 AND symb_decoder(16#ee#)) OR
 					(reg_q618 AND symb_decoder(16#84#)) OR
 					(reg_q618 AND symb_decoder(16#a0#)) OR
 					(reg_q618 AND symb_decoder(16#ce#)) OR
 					(reg_q618 AND symb_decoder(16#59#)) OR
 					(reg_q618 AND symb_decoder(16#f7#)) OR
 					(reg_q618 AND symb_decoder(16#42#)) OR
 					(reg_q618 AND symb_decoder(16#56#)) OR
 					(reg_q618 AND symb_decoder(16#c5#)) OR
 					(reg_q618 AND symb_decoder(16#52#)) OR
 					(reg_q618 AND symb_decoder(16#78#)) OR
 					(reg_q618 AND symb_decoder(16#ef#)) OR
 					(reg_q618 AND symb_decoder(16#a2#)) OR
 					(reg_q618 AND symb_decoder(16#93#)) OR
 					(reg_q618 AND symb_decoder(16#de#)) OR
 					(reg_q618 AND symb_decoder(16#21#)) OR
 					(reg_q618 AND symb_decoder(16#ff#)) OR
 					(reg_q618 AND symb_decoder(16#8c#)) OR
 					(reg_q618 AND symb_decoder(16#6c#)) OR
 					(reg_q618 AND symb_decoder(16#49#)) OR
 					(reg_q618 AND symb_decoder(16#57#)) OR
 					(reg_q618 AND symb_decoder(16#4a#)) OR
 					(reg_q618 AND symb_decoder(16#64#)) OR
 					(reg_q618 AND symb_decoder(16#92#)) OR
 					(reg_q616 AND symb_decoder(16#5b#)) OR
 					(reg_q616 AND symb_decoder(16#82#)) OR
 					(reg_q616 AND symb_decoder(16#98#)) OR
 					(reg_q616 AND symb_decoder(16#74#)) OR
 					(reg_q616 AND symb_decoder(16#1b#)) OR
 					(reg_q616 AND symb_decoder(16#bf#)) OR
 					(reg_q616 AND symb_decoder(16#f9#)) OR
 					(reg_q616 AND symb_decoder(16#19#)) OR
 					(reg_q616 AND symb_decoder(16#dd#)) OR
 					(reg_q616 AND symb_decoder(16#ff#)) OR
 					(reg_q616 AND symb_decoder(16#d7#)) OR
 					(reg_q616 AND symb_decoder(16#b6#)) OR
 					(reg_q616 AND symb_decoder(16#41#)) OR
 					(reg_q616 AND symb_decoder(16#53#)) OR
 					(reg_q616 AND symb_decoder(16#ae#)) OR
 					(reg_q616 AND symb_decoder(16#2e#)) OR
 					(reg_q616 AND symb_decoder(16#38#)) OR
 					(reg_q616 AND symb_decoder(16#c4#)) OR
 					(reg_q616 AND symb_decoder(16#d3#)) OR
 					(reg_q616 AND symb_decoder(16#c0#)) OR
 					(reg_q616 AND symb_decoder(16#b1#)) OR
 					(reg_q616 AND symb_decoder(16#ed#)) OR
 					(reg_q616 AND symb_decoder(16#be#)) OR
 					(reg_q616 AND symb_decoder(16#0b#)) OR
 					(reg_q616 AND symb_decoder(16#72#)) OR
 					(reg_q616 AND symb_decoder(16#a0#)) OR
 					(reg_q616 AND symb_decoder(16#17#)) OR
 					(reg_q616 AND symb_decoder(16#25#)) OR
 					(reg_q616 AND symb_decoder(16#ea#)) OR
 					(reg_q616 AND symb_decoder(16#32#)) OR
 					(reg_q616 AND symb_decoder(16#ee#)) OR
 					(reg_q616 AND symb_decoder(16#60#)) OR
 					(reg_q616 AND symb_decoder(16#56#)) OR
 					(reg_q616 AND symb_decoder(16#bb#)) OR
 					(reg_q616 AND symb_decoder(16#b4#)) OR
 					(reg_q616 AND symb_decoder(16#45#)) OR
 					(reg_q616 AND symb_decoder(16#69#)) OR
 					(reg_q616 AND symb_decoder(16#86#)) OR
 					(reg_q616 AND symb_decoder(16#33#)) OR
 					(reg_q616 AND symb_decoder(16#3a#)) OR
 					(reg_q616 AND symb_decoder(16#44#)) OR
 					(reg_q616 AND symb_decoder(16#93#)) OR
 					(reg_q616 AND symb_decoder(16#f2#)) OR
 					(reg_q616 AND symb_decoder(16#9c#)) OR
 					(reg_q616 AND symb_decoder(16#fc#)) OR
 					(reg_q616 AND symb_decoder(16#ca#)) OR
 					(reg_q616 AND symb_decoder(16#1e#)) OR
 					(reg_q616 AND symb_decoder(16#a1#)) OR
 					(reg_q616 AND symb_decoder(16#90#)) OR
 					(reg_q616 AND symb_decoder(16#5d#)) OR
 					(reg_q616 AND symb_decoder(16#bc#)) OR
 					(reg_q616 AND symb_decoder(16#5a#)) OR
 					(reg_q616 AND symb_decoder(16#2d#)) OR
 					(reg_q616 AND symb_decoder(16#f5#)) OR
 					(reg_q616 AND symb_decoder(16#35#)) OR
 					(reg_q616 AND symb_decoder(16#a9#)) OR
 					(reg_q616 AND symb_decoder(16#97#)) OR
 					(reg_q616 AND symb_decoder(16#80#)) OR
 					(reg_q616 AND symb_decoder(16#9f#)) OR
 					(reg_q616 AND symb_decoder(16#df#)) OR
 					(reg_q616 AND symb_decoder(16#c2#)) OR
 					(reg_q616 AND symb_decoder(16#eb#)) OR
 					(reg_q616 AND symb_decoder(16#30#)) OR
 					(reg_q616 AND symb_decoder(16#12#)) OR
 					(reg_q616 AND symb_decoder(16#f7#)) OR
 					(reg_q616 AND symb_decoder(16#2b#)) OR
 					(reg_q616 AND symb_decoder(16#a7#)) OR
 					(reg_q616 AND symb_decoder(16#15#)) OR
 					(reg_q616 AND symb_decoder(16#78#)) OR
 					(reg_q616 AND symb_decoder(16#e5#)) OR
 					(reg_q616 AND symb_decoder(16#06#)) OR
 					(reg_q616 AND symb_decoder(16#4b#)) OR
 					(reg_q616 AND symb_decoder(16#24#)) OR
 					(reg_q616 AND symb_decoder(16#55#)) OR
 					(reg_q616 AND symb_decoder(16#ef#)) OR
 					(reg_q616 AND symb_decoder(16#3d#)) OR
 					(reg_q616 AND symb_decoder(16#26#)) OR
 					(reg_q616 AND symb_decoder(16#da#)) OR
 					(reg_q616 AND symb_decoder(16#e7#)) OR
 					(reg_q616 AND symb_decoder(16#36#)) OR
 					(reg_q616 AND symb_decoder(16#43#)) OR
 					(reg_q616 AND symb_decoder(16#e8#)) OR
 					(reg_q616 AND symb_decoder(16#c1#)) OR
 					(reg_q616 AND symb_decoder(16#95#)) OR
 					(reg_q616 AND symb_decoder(16#91#)) OR
 					(reg_q616 AND symb_decoder(16#1c#)) OR
 					(reg_q616 AND symb_decoder(16#75#)) OR
 					(reg_q616 AND symb_decoder(16#9b#)) OR
 					(reg_q616 AND symb_decoder(16#16#)) OR
 					(reg_q616 AND symb_decoder(16#46#)) OR
 					(reg_q616 AND symb_decoder(16#84#)) OR
 					(reg_q616 AND symb_decoder(16#48#)) OR
 					(reg_q616 AND symb_decoder(16#cc#)) OR
 					(reg_q616 AND symb_decoder(16#f3#)) OR
 					(reg_q616 AND symb_decoder(16#8e#)) OR
 					(reg_q616 AND symb_decoder(16#d5#)) OR
 					(reg_q616 AND symb_decoder(16#e9#)) OR
 					(reg_q616 AND symb_decoder(16#3b#)) OR
 					(reg_q616 AND symb_decoder(16#3e#)) OR
 					(reg_q616 AND symb_decoder(16#88#)) OR
 					(reg_q616 AND symb_decoder(16#f4#)) OR
 					(reg_q616 AND symb_decoder(16#ac#)) OR
 					(reg_q616 AND symb_decoder(16#e1#)) OR
 					(reg_q616 AND symb_decoder(16#c3#)) OR
 					(reg_q616 AND symb_decoder(16#c7#)) OR
 					(reg_q616 AND symb_decoder(16#63#)) OR
 					(reg_q616 AND symb_decoder(16#08#)) OR
 					(reg_q616 AND symb_decoder(16#d9#)) OR
 					(reg_q616 AND symb_decoder(16#79#)) OR
 					(reg_q616 AND symb_decoder(16#d2#)) OR
 					(reg_q616 AND symb_decoder(16#47#)) OR
 					(reg_q616 AND symb_decoder(16#76#)) OR
 					(reg_q616 AND symb_decoder(16#29#)) OR
 					(reg_q616 AND symb_decoder(16#65#)) OR
 					(reg_q616 AND symb_decoder(16#39#)) OR
 					(reg_q616 AND symb_decoder(16#a8#)) OR
 					(reg_q616 AND symb_decoder(16#7a#)) OR
 					(reg_q616 AND symb_decoder(16#31#)) OR
 					(reg_q616 AND symb_decoder(16#4c#)) OR
 					(reg_q616 AND symb_decoder(16#27#)) OR
 					(reg_q616 AND symb_decoder(16#07#)) OR
 					(reg_q616 AND symb_decoder(16#8c#)) OR
 					(reg_q616 AND symb_decoder(16#89#)) OR
 					(reg_q616 AND symb_decoder(16#5c#)) OR
 					(reg_q616 AND symb_decoder(16#b3#)) OR
 					(reg_q616 AND symb_decoder(16#22#)) OR
 					(reg_q616 AND symb_decoder(16#01#)) OR
 					(reg_q616 AND symb_decoder(16#de#)) OR
 					(reg_q616 AND symb_decoder(16#ab#)) OR
 					(reg_q616 AND symb_decoder(16#87#)) OR
 					(reg_q616 AND symb_decoder(16#14#)) OR
 					(reg_q616 AND symb_decoder(16#1a#)) OR
 					(reg_q616 AND symb_decoder(16#58#)) OR
 					(reg_q616 AND symb_decoder(16#11#)) OR
 					(reg_q616 AND symb_decoder(16#6f#)) OR
 					(reg_q616 AND symb_decoder(16#37#)) OR
 					(reg_q616 AND symb_decoder(16#02#)) OR
 					(reg_q616 AND symb_decoder(16#ce#)) OR
 					(reg_q616 AND symb_decoder(16#9a#)) OR
 					(reg_q616 AND symb_decoder(16#b5#)) OR
 					(reg_q616 AND symb_decoder(16#94#)) OR
 					(reg_q616 AND symb_decoder(16#6d#)) OR
 					(reg_q616 AND symb_decoder(16#04#)) OR
 					(reg_q616 AND symb_decoder(16#8f#)) OR
 					(reg_q616 AND symb_decoder(16#71#)) OR
 					(reg_q616 AND symb_decoder(16#b2#)) OR
 					(reg_q616 AND symb_decoder(16#73#)) OR
 					(reg_q616 AND symb_decoder(16#7e#)) OR
 					(reg_q616 AND symb_decoder(16#81#)) OR
 					(reg_q616 AND symb_decoder(16#4e#)) OR
 					(reg_q616 AND symb_decoder(16#52#)) OR
 					(reg_q616 AND symb_decoder(16#bd#)) OR
 					(reg_q616 AND symb_decoder(16#f6#)) OR
 					(reg_q616 AND symb_decoder(16#50#)) OR
 					(reg_q616 AND symb_decoder(16#6e#)) OR
 					(reg_q616 AND symb_decoder(16#96#)) OR
 					(reg_q616 AND symb_decoder(16#d8#)) OR
 					(reg_q616 AND symb_decoder(16#e4#)) OR
 					(reg_q616 AND symb_decoder(16#92#)) OR
 					(reg_q616 AND symb_decoder(16#4d#)) OR
 					(reg_q616 AND symb_decoder(16#a2#)) OR
 					(reg_q616 AND symb_decoder(16#ec#)) OR
 					(reg_q616 AND symb_decoder(16#b9#)) OR
 					(reg_q616 AND symb_decoder(16#d6#)) OR
 					(reg_q616 AND symb_decoder(16#64#)) OR
 					(reg_q616 AND symb_decoder(16#8b#)) OR
 					(reg_q616 AND symb_decoder(16#1d#)) OR
 					(reg_q616 AND symb_decoder(16#8a#)) OR
 					(reg_q616 AND symb_decoder(16#c8#)) OR
 					(reg_q616 AND symb_decoder(16#4a#)) OR
 					(reg_q616 AND symb_decoder(16#fe#)) OR
 					(reg_q616 AND symb_decoder(16#4f#)) OR
 					(reg_q616 AND symb_decoder(16#9e#)) OR
 					(reg_q616 AND symb_decoder(16#40#)) OR
 					(reg_q616 AND symb_decoder(16#7b#)) OR
 					(reg_q616 AND symb_decoder(16#e2#)) OR
 					(reg_q616 AND symb_decoder(16#f8#)) OR
 					(reg_q616 AND symb_decoder(16#a3#)) OR
 					(reg_q616 AND symb_decoder(16#7d#)) OR
 					(reg_q616 AND symb_decoder(16#34#)) OR
 					(reg_q616 AND symb_decoder(16#b0#)) OR
 					(reg_q616 AND symb_decoder(16#2a#)) OR
 					(reg_q616 AND symb_decoder(16#c9#)) OR
 					(reg_q616 AND symb_decoder(16#18#)) OR
 					(reg_q616 AND symb_decoder(16#59#)) OR
 					(reg_q616 AND symb_decoder(16#6b#)) OR
 					(reg_q616 AND symb_decoder(16#70#)) OR
 					(reg_q616 AND symb_decoder(16#cd#)) OR
 					(reg_q616 AND symb_decoder(16#aa#)) OR
 					(reg_q616 AND symb_decoder(16#00#)) OR
 					(reg_q616 AND symb_decoder(16#dc#)) OR
 					(reg_q616 AND symb_decoder(16#85#)) OR
 					(reg_q616 AND symb_decoder(16#05#)) OR
 					(reg_q616 AND symb_decoder(16#62#)) OR
 					(reg_q616 AND symb_decoder(16#57#)) OR
 					(reg_q616 AND symb_decoder(16#ad#)) OR
 					(reg_q616 AND symb_decoder(16#28#)) OR
 					(reg_q616 AND symb_decoder(16#13#)) OR
 					(reg_q616 AND symb_decoder(16#c5#)) OR
 					(reg_q616 AND symb_decoder(16#67#)) OR
 					(reg_q616 AND symb_decoder(16#db#)) OR
 					(reg_q616 AND symb_decoder(16#2f#)) OR
 					(reg_q616 AND symb_decoder(16#5f#)) OR
 					(reg_q616 AND symb_decoder(16#03#)) OR
 					(reg_q616 AND symb_decoder(16#f0#)) OR
 					(reg_q616 AND symb_decoder(16#2c#)) OR
 					(reg_q616 AND symb_decoder(16#a5#)) OR
 					(reg_q616 AND symb_decoder(16#6c#)) OR
 					(reg_q616 AND symb_decoder(16#6a#)) OR
 					(reg_q616 AND symb_decoder(16#10#)) OR
 					(reg_q616 AND symb_decoder(16#66#)) OR
 					(reg_q616 AND symb_decoder(16#cb#)) OR
 					(reg_q616 AND symb_decoder(16#b8#)) OR
 					(reg_q616 AND symb_decoder(16#fa#)) OR
 					(reg_q616 AND symb_decoder(16#7f#)) OR
 					(reg_q616 AND symb_decoder(16#3f#)) OR
 					(reg_q616 AND symb_decoder(16#fd#)) OR
 					(reg_q616 AND symb_decoder(16#7c#)) OR
 					(reg_q616 AND symb_decoder(16#3c#)) OR
 					(reg_q616 AND symb_decoder(16#61#)) OR
 					(reg_q616 AND symb_decoder(16#8d#)) OR
 					(reg_q616 AND symb_decoder(16#68#)) OR
 					(reg_q616 AND symb_decoder(16#d4#)) OR
 					(reg_q616 AND symb_decoder(16#5e#)) OR
 					(reg_q616 AND symb_decoder(16#0f#)) OR
 					(reg_q616 AND symb_decoder(16#f1#)) OR
 					(reg_q616 AND symb_decoder(16#af#)) OR
 					(reg_q616 AND symb_decoder(16#54#)) OR
 					(reg_q616 AND symb_decoder(16#a6#)) OR
 					(reg_q616 AND symb_decoder(16#99#)) OR
 					(reg_q616 AND symb_decoder(16#77#)) OR
 					(reg_q616 AND symb_decoder(16#c6#)) OR
 					(reg_q616 AND symb_decoder(16#83#)) OR
 					(reg_q616 AND symb_decoder(16#cf#)) OR
 					(reg_q616 AND symb_decoder(16#21#)) OR
 					(reg_q616 AND symb_decoder(16#51#)) OR
 					(reg_q616 AND symb_decoder(16#a4#)) OR
 					(reg_q616 AND symb_decoder(16#1f#)) OR
 					(reg_q616 AND symb_decoder(16#49#)) OR
 					(reg_q616 AND symb_decoder(16#e3#)) OR
 					(reg_q616 AND symb_decoder(16#d1#)) OR
 					(reg_q616 AND symb_decoder(16#42#)) OR
 					(reg_q616 AND symb_decoder(16#9d#)) OR
 					(reg_q616 AND symb_decoder(16#ba#)) OR
 					(reg_q616 AND symb_decoder(16#0e#)) OR
 					(reg_q616 AND symb_decoder(16#e0#)) OR
 					(reg_q616 AND symb_decoder(16#d0#)) OR
 					(reg_q616 AND symb_decoder(16#e6#)) OR
 					(reg_q616 AND symb_decoder(16#b7#)) OR
 					(reg_q616 AND symb_decoder(16#fb#)) OR
 					(reg_q616 AND symb_decoder(16#23#));
reg_q618_init <= '0' ;
	p_reg_q618: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q618 <= reg_q618_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q618 <= reg_q618_init;
        else
          reg_q618 <= reg_q618_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1359_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1359 AND symb_decoder(16#e5#)) OR
 					(reg_q1359 AND symb_decoder(16#18#)) OR
 					(reg_q1359 AND symb_decoder(16#d2#)) OR
 					(reg_q1359 AND symb_decoder(16#d6#)) OR
 					(reg_q1359 AND symb_decoder(16#de#)) OR
 					(reg_q1359 AND symb_decoder(16#a8#)) OR
 					(reg_q1359 AND symb_decoder(16#57#)) OR
 					(reg_q1359 AND symb_decoder(16#3b#)) OR
 					(reg_q1359 AND symb_decoder(16#fe#)) OR
 					(reg_q1359 AND symb_decoder(16#30#)) OR
 					(reg_q1359 AND symb_decoder(16#e8#)) OR
 					(reg_q1359 AND symb_decoder(16#27#)) OR
 					(reg_q1359 AND symb_decoder(16#12#)) OR
 					(reg_q1359 AND symb_decoder(16#40#)) OR
 					(reg_q1359 AND symb_decoder(16#9f#)) OR
 					(reg_q1359 AND symb_decoder(16#4c#)) OR
 					(reg_q1359 AND symb_decoder(16#b6#)) OR
 					(reg_q1359 AND symb_decoder(16#a1#)) OR
 					(reg_q1359 AND symb_decoder(16#e6#)) OR
 					(reg_q1359 AND symb_decoder(16#65#)) OR
 					(reg_q1359 AND symb_decoder(16#b2#)) OR
 					(reg_q1359 AND symb_decoder(16#72#)) OR
 					(reg_q1359 AND symb_decoder(16#61#)) OR
 					(reg_q1359 AND symb_decoder(16#f5#)) OR
 					(reg_q1359 AND symb_decoder(16#55#)) OR
 					(reg_q1359 AND symb_decoder(16#94#)) OR
 					(reg_q1359 AND symb_decoder(16#9c#)) OR
 					(reg_q1359 AND symb_decoder(16#01#)) OR
 					(reg_q1359 AND symb_decoder(16#4f#)) OR
 					(reg_q1359 AND symb_decoder(16#f8#)) OR
 					(reg_q1359 AND symb_decoder(16#c3#)) OR
 					(reg_q1359 AND symb_decoder(16#ef#)) OR
 					(reg_q1359 AND symb_decoder(16#b8#)) OR
 					(reg_q1359 AND symb_decoder(16#ed#)) OR
 					(reg_q1359 AND symb_decoder(16#76#)) OR
 					(reg_q1359 AND symb_decoder(16#c2#)) OR
 					(reg_q1359 AND symb_decoder(16#b1#)) OR
 					(reg_q1359 AND symb_decoder(16#c8#)) OR
 					(reg_q1359 AND symb_decoder(16#11#)) OR
 					(reg_q1359 AND symb_decoder(16#64#)) OR
 					(reg_q1359 AND symb_decoder(16#69#)) OR
 					(reg_q1359 AND symb_decoder(16#a9#)) OR
 					(reg_q1359 AND symb_decoder(16#3e#)) OR
 					(reg_q1359 AND symb_decoder(16#f9#)) OR
 					(reg_q1359 AND symb_decoder(16#38#)) OR
 					(reg_q1359 AND symb_decoder(16#2e#)) OR
 					(reg_q1359 AND symb_decoder(16#ee#)) OR
 					(reg_q1359 AND symb_decoder(16#88#)) OR
 					(reg_q1359 AND symb_decoder(16#a5#)) OR
 					(reg_q1359 AND symb_decoder(16#d0#)) OR
 					(reg_q1359 AND symb_decoder(16#b7#)) OR
 					(reg_q1359 AND symb_decoder(16#22#)) OR
 					(reg_q1359 AND symb_decoder(16#ad#)) OR
 					(reg_q1359 AND symb_decoder(16#4b#)) OR
 					(reg_q1359 AND symb_decoder(16#bf#)) OR
 					(reg_q1359 AND symb_decoder(16#52#)) OR
 					(reg_q1359 AND symb_decoder(16#02#)) OR
 					(reg_q1359 AND symb_decoder(16#82#)) OR
 					(reg_q1359 AND symb_decoder(16#26#)) OR
 					(reg_q1359 AND symb_decoder(16#2b#)) OR
 					(reg_q1359 AND symb_decoder(16#14#)) OR
 					(reg_q1359 AND symb_decoder(16#5f#)) OR
 					(reg_q1359 AND symb_decoder(16#03#)) OR
 					(reg_q1359 AND symb_decoder(16#37#)) OR
 					(reg_q1359 AND symb_decoder(16#7c#)) OR
 					(reg_q1359 AND symb_decoder(16#d1#)) OR
 					(reg_q1359 AND symb_decoder(16#b3#)) OR
 					(reg_q1359 AND symb_decoder(16#51#)) OR
 					(reg_q1359 AND symb_decoder(16#d3#)) OR
 					(reg_q1359 AND symb_decoder(16#1d#)) OR
 					(reg_q1359 AND symb_decoder(16#aa#)) OR
 					(reg_q1359 AND symb_decoder(16#0f#)) OR
 					(reg_q1359 AND symb_decoder(16#29#)) OR
 					(reg_q1359 AND symb_decoder(16#98#)) OR
 					(reg_q1359 AND symb_decoder(16#46#)) OR
 					(reg_q1359 AND symb_decoder(16#0a#)) OR
 					(reg_q1359 AND symb_decoder(16#83#)) OR
 					(reg_q1359 AND symb_decoder(16#ea#)) OR
 					(reg_q1359 AND symb_decoder(16#a4#)) OR
 					(reg_q1359 AND symb_decoder(16#4a#)) OR
 					(reg_q1359 AND symb_decoder(16#47#)) OR
 					(reg_q1359 AND symb_decoder(16#7f#)) OR
 					(reg_q1359 AND symb_decoder(16#3f#)) OR
 					(reg_q1359 AND symb_decoder(16#c5#)) OR
 					(reg_q1359 AND symb_decoder(16#8b#)) OR
 					(reg_q1359 AND symb_decoder(16#ae#)) OR
 					(reg_q1359 AND symb_decoder(16#f6#)) OR
 					(reg_q1359 AND symb_decoder(16#0c#)) OR
 					(reg_q1359 AND symb_decoder(16#4d#)) OR
 					(reg_q1359 AND symb_decoder(16#56#)) OR
 					(reg_q1359 AND symb_decoder(16#8d#)) OR
 					(reg_q1359 AND symb_decoder(16#42#)) OR
 					(reg_q1359 AND symb_decoder(16#a6#)) OR
 					(reg_q1359 AND symb_decoder(16#e9#)) OR
 					(reg_q1359 AND symb_decoder(16#c6#)) OR
 					(reg_q1359 AND symb_decoder(16#2d#)) OR
 					(reg_q1359 AND symb_decoder(16#97#)) OR
 					(reg_q1359 AND symb_decoder(16#0b#)) OR
 					(reg_q1359 AND symb_decoder(16#28#)) OR
 					(reg_q1359 AND symb_decoder(16#09#)) OR
 					(reg_q1359 AND symb_decoder(16#af#)) OR
 					(reg_q1359 AND symb_decoder(16#15#)) OR
 					(reg_q1359 AND symb_decoder(16#7d#)) OR
 					(reg_q1359 AND symb_decoder(16#9d#)) OR
 					(reg_q1359 AND symb_decoder(16#48#)) OR
 					(reg_q1359 AND symb_decoder(16#35#)) OR
 					(reg_q1359 AND symb_decoder(16#c9#)) OR
 					(reg_q1359 AND symb_decoder(16#5b#)) OR
 					(reg_q1359 AND symb_decoder(16#45#)) OR
 					(reg_q1359 AND symb_decoder(16#7e#)) OR
 					(reg_q1359 AND symb_decoder(16#a2#)) OR
 					(reg_q1359 AND symb_decoder(16#fd#)) OR
 					(reg_q1359 AND symb_decoder(16#ec#)) OR
 					(reg_q1359 AND symb_decoder(16#84#)) OR
 					(reg_q1359 AND symb_decoder(16#75#)) OR
 					(reg_q1359 AND symb_decoder(16#23#)) OR
 					(reg_q1359 AND symb_decoder(16#c1#)) OR
 					(reg_q1359 AND symb_decoder(16#63#)) OR
 					(reg_q1359 AND symb_decoder(16#dc#)) OR
 					(reg_q1359 AND symb_decoder(16#68#)) OR
 					(reg_q1359 AND symb_decoder(16#ce#)) OR
 					(reg_q1359 AND symb_decoder(16#2c#)) OR
 					(reg_q1359 AND symb_decoder(16#66#)) OR
 					(reg_q1359 AND symb_decoder(16#db#)) OR
 					(reg_q1359 AND symb_decoder(16#e4#)) OR
 					(reg_q1359 AND symb_decoder(16#ac#)) OR
 					(reg_q1359 AND symb_decoder(16#3d#)) OR
 					(reg_q1359 AND symb_decoder(16#fa#)) OR
 					(reg_q1359 AND symb_decoder(16#be#)) OR
 					(reg_q1359 AND symb_decoder(16#90#)) OR
 					(reg_q1359 AND symb_decoder(16#ab#)) OR
 					(reg_q1359 AND symb_decoder(16#73#)) OR
 					(reg_q1359 AND symb_decoder(16#50#)) OR
 					(reg_q1359 AND symb_decoder(16#0d#)) OR
 					(reg_q1359 AND symb_decoder(16#16#)) OR
 					(reg_q1359 AND symb_decoder(16#8c#)) OR
 					(reg_q1359 AND symb_decoder(16#bb#)) OR
 					(reg_q1359 AND symb_decoder(16#21#)) OR
 					(reg_q1359 AND symb_decoder(16#dd#)) OR
 					(reg_q1359 AND symb_decoder(16#d9#)) OR
 					(reg_q1359 AND symb_decoder(16#1e#)) OR
 					(reg_q1359 AND symb_decoder(16#2f#)) OR
 					(reg_q1359 AND symb_decoder(16#fc#)) OR
 					(reg_q1359 AND symb_decoder(16#ba#)) OR
 					(reg_q1359 AND symb_decoder(16#67#)) OR
 					(reg_q1359 AND symb_decoder(16#5e#)) OR
 					(reg_q1359 AND symb_decoder(16#24#)) OR
 					(reg_q1359 AND symb_decoder(16#8e#)) OR
 					(reg_q1359 AND symb_decoder(16#f0#)) OR
 					(reg_q1359 AND symb_decoder(16#59#)) OR
 					(reg_q1359 AND symb_decoder(16#19#)) OR
 					(reg_q1359 AND symb_decoder(16#5c#)) OR
 					(reg_q1359 AND symb_decoder(16#c0#)) OR
 					(reg_q1359 AND symb_decoder(16#bd#)) OR
 					(reg_q1359 AND symb_decoder(16#05#)) OR
 					(reg_q1359 AND symb_decoder(16#54#)) OR
 					(reg_q1359 AND symb_decoder(16#9a#)) OR
 					(reg_q1359 AND symb_decoder(16#f2#)) OR
 					(reg_q1359 AND symb_decoder(16#7a#)) OR
 					(reg_q1359 AND symb_decoder(16#10#)) OR
 					(reg_q1359 AND symb_decoder(16#17#)) OR
 					(reg_q1359 AND symb_decoder(16#6d#)) OR
 					(reg_q1359 AND symb_decoder(16#85#)) OR
 					(reg_q1359 AND symb_decoder(16#79#)) OR
 					(reg_q1359 AND symb_decoder(16#74#)) OR
 					(reg_q1359 AND symb_decoder(16#9b#)) OR
 					(reg_q1359 AND symb_decoder(16#df#)) OR
 					(reg_q1359 AND symb_decoder(16#0e#)) OR
 					(reg_q1359 AND symb_decoder(16#43#)) OR
 					(reg_q1359 AND symb_decoder(16#96#)) OR
 					(reg_q1359 AND symb_decoder(16#81#)) OR
 					(reg_q1359 AND symb_decoder(16#07#)) OR
 					(reg_q1359 AND symb_decoder(16#5a#)) OR
 					(reg_q1359 AND symb_decoder(16#cf#)) OR
 					(reg_q1359 AND symb_decoder(16#e3#)) OR
 					(reg_q1359 AND symb_decoder(16#58#)) OR
 					(reg_q1359 AND symb_decoder(16#34#)) OR
 					(reg_q1359 AND symb_decoder(16#92#)) OR
 					(reg_q1359 AND symb_decoder(16#1f#)) OR
 					(reg_q1359 AND symb_decoder(16#2a#)) OR
 					(reg_q1359 AND symb_decoder(16#b5#)) OR
 					(reg_q1359 AND symb_decoder(16#3a#)) OR
 					(reg_q1359 AND symb_decoder(16#87#)) OR
 					(reg_q1359 AND symb_decoder(16#d7#)) OR
 					(reg_q1359 AND symb_decoder(16#6c#)) OR
 					(reg_q1359 AND symb_decoder(16#08#)) OR
 					(reg_q1359 AND symb_decoder(16#71#)) OR
 					(reg_q1359 AND symb_decoder(16#e2#)) OR
 					(reg_q1359 AND symb_decoder(16#62#)) OR
 					(reg_q1359 AND symb_decoder(16#04#)) OR
 					(reg_q1359 AND symb_decoder(16#86#)) OR
 					(reg_q1359 AND symb_decoder(16#b4#)) OR
 					(reg_q1359 AND symb_decoder(16#c4#)) OR
 					(reg_q1359 AND symb_decoder(16#bc#)) OR
 					(reg_q1359 AND symb_decoder(16#32#)) OR
 					(reg_q1359 AND symb_decoder(16#ff#)) OR
 					(reg_q1359 AND symb_decoder(16#d4#)) OR
 					(reg_q1359 AND symb_decoder(16#1c#)) OR
 					(reg_q1359 AND symb_decoder(16#31#)) OR
 					(reg_q1359 AND symb_decoder(16#e7#)) OR
 					(reg_q1359 AND symb_decoder(16#b9#)) OR
 					(reg_q1359 AND symb_decoder(16#6e#)) OR
 					(reg_q1359 AND symb_decoder(16#f7#)) OR
 					(reg_q1359 AND symb_decoder(16#a3#)) OR
 					(reg_q1359 AND symb_decoder(16#53#)) OR
 					(reg_q1359 AND symb_decoder(16#cb#)) OR
 					(reg_q1359 AND symb_decoder(16#91#)) OR
 					(reg_q1359 AND symb_decoder(16#33#)) OR
 					(reg_q1359 AND symb_decoder(16#3c#)) OR
 					(reg_q1359 AND symb_decoder(16#4e#)) OR
 					(reg_q1359 AND symb_decoder(16#f4#)) OR
 					(reg_q1359 AND symb_decoder(16#93#)) OR
 					(reg_q1359 AND symb_decoder(16#20#)) OR
 					(reg_q1359 AND symb_decoder(16#6f#)) OR
 					(reg_q1359 AND symb_decoder(16#80#)) OR
 					(reg_q1359 AND symb_decoder(16#f1#)) OR
 					(reg_q1359 AND symb_decoder(16#8f#)) OR
 					(reg_q1359 AND symb_decoder(16#a7#)) OR
 					(reg_q1359 AND symb_decoder(16#6a#)) OR
 					(reg_q1359 AND symb_decoder(16#c7#)) OR
 					(reg_q1359 AND symb_decoder(16#89#)) OR
 					(reg_q1359 AND symb_decoder(16#d8#)) OR
 					(reg_q1359 AND symb_decoder(16#60#)) OR
 					(reg_q1359 AND symb_decoder(16#36#)) OR
 					(reg_q1359 AND symb_decoder(16#cc#)) OR
 					(reg_q1359 AND symb_decoder(16#ca#)) OR
 					(reg_q1359 AND symb_decoder(16#00#)) OR
 					(reg_q1359 AND symb_decoder(16#49#)) OR
 					(reg_q1359 AND symb_decoder(16#44#)) OR
 					(reg_q1359 AND symb_decoder(16#70#)) OR
 					(reg_q1359 AND symb_decoder(16#e0#)) OR
 					(reg_q1359 AND symb_decoder(16#95#)) OR
 					(reg_q1359 AND symb_decoder(16#d5#)) OR
 					(reg_q1359 AND symb_decoder(16#cd#)) OR
 					(reg_q1359 AND symb_decoder(16#7b#)) OR
 					(reg_q1359 AND symb_decoder(16#77#)) OR
 					(reg_q1359 AND symb_decoder(16#e1#)) OR
 					(reg_q1359 AND symb_decoder(16#99#)) OR
 					(reg_q1359 AND symb_decoder(16#13#)) OR
 					(reg_q1359 AND symb_decoder(16#5d#)) OR
 					(reg_q1359 AND symb_decoder(16#8a#)) OR
 					(reg_q1359 AND symb_decoder(16#b0#)) OR
 					(reg_q1359 AND symb_decoder(16#41#)) OR
 					(reg_q1359 AND symb_decoder(16#39#)) OR
 					(reg_q1359 AND symb_decoder(16#eb#)) OR
 					(reg_q1359 AND symb_decoder(16#25#)) OR
 					(reg_q1359 AND symb_decoder(16#9e#)) OR
 					(reg_q1359 AND symb_decoder(16#da#)) OR
 					(reg_q1359 AND symb_decoder(16#78#)) OR
 					(reg_q1359 AND symb_decoder(16#06#)) OR
 					(reg_q1359 AND symb_decoder(16#fb#)) OR
 					(reg_q1359 AND symb_decoder(16#6b#)) OR
 					(reg_q1359 AND symb_decoder(16#1b#)) OR
 					(reg_q1359 AND symb_decoder(16#a0#)) OR
 					(reg_q1359 AND symb_decoder(16#1a#)) OR
 					(reg_q1359 AND symb_decoder(16#f3#));
reg_q1359_init <= '0' ;
	p_reg_q1359: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1359 <= reg_q1359_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1359 <= reg_q1359_init;
        else
          reg_q1359 <= reg_q1359_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2052_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2052 AND symb_decoder(16#0e#)) OR
 					(reg_q2052 AND symb_decoder(16#af#)) OR
 					(reg_q2052 AND symb_decoder(16#9b#)) OR
 					(reg_q2052 AND symb_decoder(16#ed#)) OR
 					(reg_q2052 AND symb_decoder(16#de#)) OR
 					(reg_q2052 AND symb_decoder(16#37#)) OR
 					(reg_q2052 AND symb_decoder(16#54#)) OR
 					(reg_q2052 AND symb_decoder(16#78#)) OR
 					(reg_q2052 AND symb_decoder(16#c5#)) OR
 					(reg_q2052 AND symb_decoder(16#0f#)) OR
 					(reg_q2052 AND symb_decoder(16#bb#)) OR
 					(reg_q2052 AND symb_decoder(16#79#)) OR
 					(reg_q2052 AND symb_decoder(16#cd#)) OR
 					(reg_q2052 AND symb_decoder(16#b0#)) OR
 					(reg_q2052 AND symb_decoder(16#60#)) OR
 					(reg_q2052 AND symb_decoder(16#d8#)) OR
 					(reg_q2052 AND symb_decoder(16#39#)) OR
 					(reg_q2052 AND symb_decoder(16#4a#)) OR
 					(reg_q2052 AND symb_decoder(16#08#)) OR
 					(reg_q2052 AND symb_decoder(16#ba#)) OR
 					(reg_q2052 AND symb_decoder(16#7f#)) OR
 					(reg_q2052 AND symb_decoder(16#02#)) OR
 					(reg_q2052 AND symb_decoder(16#8e#)) OR
 					(reg_q2052 AND symb_decoder(16#6f#)) OR
 					(reg_q2052 AND symb_decoder(16#e0#)) OR
 					(reg_q2052 AND symb_decoder(16#e7#)) OR
 					(reg_q2052 AND symb_decoder(16#2d#)) OR
 					(reg_q2052 AND symb_decoder(16#10#)) OR
 					(reg_q2052 AND symb_decoder(16#8a#)) OR
 					(reg_q2052 AND symb_decoder(16#8b#)) OR
 					(reg_q2052 AND symb_decoder(16#25#)) OR
 					(reg_q2052 AND symb_decoder(16#5c#)) OR
 					(reg_q2052 AND symb_decoder(16#eb#)) OR
 					(reg_q2052 AND symb_decoder(16#da#)) OR
 					(reg_q2052 AND symb_decoder(16#ee#)) OR
 					(reg_q2052 AND symb_decoder(16#49#)) OR
 					(reg_q2052 AND symb_decoder(16#01#)) OR
 					(reg_q2052 AND symb_decoder(16#f4#)) OR
 					(reg_q2052 AND symb_decoder(16#f1#)) OR
 					(reg_q2052 AND symb_decoder(16#fe#)) OR
 					(reg_q2052 AND symb_decoder(16#9f#)) OR
 					(reg_q2052 AND symb_decoder(16#4d#)) OR
 					(reg_q2052 AND symb_decoder(16#27#)) OR
 					(reg_q2052 AND symb_decoder(16#7d#)) OR
 					(reg_q2052 AND symb_decoder(16#a5#)) OR
 					(reg_q2052 AND symb_decoder(16#b3#)) OR
 					(reg_q2052 AND symb_decoder(16#e3#)) OR
 					(reg_q2052 AND symb_decoder(16#1d#)) OR
 					(reg_q2052 AND symb_decoder(16#2b#)) OR
 					(reg_q2052 AND symb_decoder(16#5b#)) OR
 					(reg_q2052 AND symb_decoder(16#e2#)) OR
 					(reg_q2052 AND symb_decoder(16#1a#)) OR
 					(reg_q2052 AND symb_decoder(16#64#)) OR
 					(reg_q2052 AND symb_decoder(16#2e#)) OR
 					(reg_q2052 AND symb_decoder(16#3a#)) OR
 					(reg_q2052 AND symb_decoder(16#42#)) OR
 					(reg_q2052 AND symb_decoder(16#33#)) OR
 					(reg_q2052 AND symb_decoder(16#77#)) OR
 					(reg_q2052 AND symb_decoder(16#b8#)) OR
 					(reg_q2052 AND symb_decoder(16#53#)) OR
 					(reg_q2052 AND symb_decoder(16#75#)) OR
 					(reg_q2052 AND symb_decoder(16#d2#)) OR
 					(reg_q2052 AND symb_decoder(16#aa#)) OR
 					(reg_q2052 AND symb_decoder(16#d7#)) OR
 					(reg_q2052 AND symb_decoder(16#06#)) OR
 					(reg_q2052 AND symb_decoder(16#52#)) OR
 					(reg_q2052 AND symb_decoder(16#48#)) OR
 					(reg_q2052 AND symb_decoder(16#0c#)) OR
 					(reg_q2052 AND symb_decoder(16#a6#)) OR
 					(reg_q2052 AND symb_decoder(16#a4#)) OR
 					(reg_q2052 AND symb_decoder(16#90#)) OR
 					(reg_q2052 AND symb_decoder(16#68#)) OR
 					(reg_q2052 AND symb_decoder(16#c2#)) OR
 					(reg_q2052 AND symb_decoder(16#71#)) OR
 					(reg_q2052 AND symb_decoder(16#1e#)) OR
 					(reg_q2052 AND symb_decoder(16#2a#)) OR
 					(reg_q2052 AND symb_decoder(16#f8#)) OR
 					(reg_q2052 AND symb_decoder(16#cf#)) OR
 					(reg_q2052 AND symb_decoder(16#12#)) OR
 					(reg_q2052 AND symb_decoder(16#19#)) OR
 					(reg_q2052 AND symb_decoder(16#97#)) OR
 					(reg_q2052 AND symb_decoder(16#a7#)) OR
 					(reg_q2052 AND symb_decoder(16#0d#)) OR
 					(reg_q2052 AND symb_decoder(16#94#)) OR
 					(reg_q2052 AND symb_decoder(16#f7#)) OR
 					(reg_q2052 AND symb_decoder(16#62#)) OR
 					(reg_q2052 AND symb_decoder(16#fa#)) OR
 					(reg_q2052 AND symb_decoder(16#7a#)) OR
 					(reg_q2052 AND symb_decoder(16#cb#)) OR
 					(reg_q2052 AND symb_decoder(16#34#)) OR
 					(reg_q2052 AND symb_decoder(16#7e#)) OR
 					(reg_q2052 AND symb_decoder(16#b5#)) OR
 					(reg_q2052 AND symb_decoder(16#ea#)) OR
 					(reg_q2052 AND symb_decoder(16#61#)) OR
 					(reg_q2052 AND symb_decoder(16#ae#)) OR
 					(reg_q2052 AND symb_decoder(16#8d#)) OR
 					(reg_q2052 AND symb_decoder(16#8f#)) OR
 					(reg_q2052 AND symb_decoder(16#65#)) OR
 					(reg_q2052 AND symb_decoder(16#03#)) OR
 					(reg_q2052 AND symb_decoder(16#87#)) OR
 					(reg_q2052 AND symb_decoder(16#5d#)) OR
 					(reg_q2052 AND symb_decoder(16#ef#)) OR
 					(reg_q2052 AND symb_decoder(16#4c#)) OR
 					(reg_q2052 AND symb_decoder(16#a1#)) OR
 					(reg_q2052 AND symb_decoder(16#c1#)) OR
 					(reg_q2052 AND symb_decoder(16#d0#)) OR
 					(reg_q2052 AND symb_decoder(16#9c#)) OR
 					(reg_q2052 AND symb_decoder(16#e9#)) OR
 					(reg_q2052 AND symb_decoder(16#f0#)) OR
 					(reg_q2052 AND symb_decoder(16#59#)) OR
 					(reg_q2052 AND symb_decoder(16#24#)) OR
 					(reg_q2052 AND symb_decoder(16#3c#)) OR
 					(reg_q2052 AND symb_decoder(16#bc#)) OR
 					(reg_q2052 AND symb_decoder(16#a0#)) OR
 					(reg_q2052 AND symb_decoder(16#50#)) OR
 					(reg_q2052 AND symb_decoder(16#40#)) OR
 					(reg_q2052 AND symb_decoder(16#44#)) OR
 					(reg_q2052 AND symb_decoder(16#3f#)) OR
 					(reg_q2052 AND symb_decoder(16#dd#)) OR
 					(reg_q2052 AND symb_decoder(16#20#)) OR
 					(reg_q2052 AND symb_decoder(16#be#)) OR
 					(reg_q2052 AND symb_decoder(16#6e#)) OR
 					(reg_q2052 AND symb_decoder(16#0a#)) OR
 					(reg_q2052 AND symb_decoder(16#d4#)) OR
 					(reg_q2052 AND symb_decoder(16#91#)) OR
 					(reg_q2052 AND symb_decoder(16#13#)) OR
 					(reg_q2052 AND symb_decoder(16#86#)) OR
 					(reg_q2052 AND symb_decoder(16#09#)) OR
 					(reg_q2052 AND symb_decoder(16#05#)) OR
 					(reg_q2052 AND symb_decoder(16#95#)) OR
 					(reg_q2052 AND symb_decoder(16#04#)) OR
 					(reg_q2052 AND symb_decoder(16#43#)) OR
 					(reg_q2052 AND symb_decoder(16#d9#)) OR
 					(reg_q2052 AND symb_decoder(16#35#)) OR
 					(reg_q2052 AND symb_decoder(16#a2#)) OR
 					(reg_q2052 AND symb_decoder(16#00#)) OR
 					(reg_q2052 AND symb_decoder(16#56#)) OR
 					(reg_q2052 AND symb_decoder(16#46#)) OR
 					(reg_q2052 AND symb_decoder(16#15#)) OR
 					(reg_q2052 AND symb_decoder(16#2c#)) OR
 					(reg_q2052 AND symb_decoder(16#ca#)) OR
 					(reg_q2052 AND symb_decoder(16#f6#)) OR
 					(reg_q2052 AND symb_decoder(16#26#)) OR
 					(reg_q2052 AND symb_decoder(16#ce#)) OR
 					(reg_q2052 AND symb_decoder(16#df#)) OR
 					(reg_q2052 AND symb_decoder(16#88#)) OR
 					(reg_q2052 AND symb_decoder(16#8c#)) OR
 					(reg_q2052 AND symb_decoder(16#36#)) OR
 					(reg_q2052 AND symb_decoder(16#ec#)) OR
 					(reg_q2052 AND symb_decoder(16#3d#)) OR
 					(reg_q2052 AND symb_decoder(16#84#)) OR
 					(reg_q2052 AND symb_decoder(16#0b#)) OR
 					(reg_q2052 AND symb_decoder(16#81#)) OR
 					(reg_q2052 AND symb_decoder(16#a8#)) OR
 					(reg_q2052 AND symb_decoder(16#bd#)) OR
 					(reg_q2052 AND symb_decoder(16#18#)) OR
 					(reg_q2052 AND symb_decoder(16#fd#)) OR
 					(reg_q2052 AND symb_decoder(16#b1#)) OR
 					(reg_q2052 AND symb_decoder(16#b9#)) OR
 					(reg_q2052 AND symb_decoder(16#ac#)) OR
 					(reg_q2052 AND symb_decoder(16#82#)) OR
 					(reg_q2052 AND symb_decoder(16#c9#)) OR
 					(reg_q2052 AND symb_decoder(16#76#)) OR
 					(reg_q2052 AND symb_decoder(16#57#)) OR
 					(reg_q2052 AND symb_decoder(16#96#)) OR
 					(reg_q2052 AND symb_decoder(16#e5#)) OR
 					(reg_q2052 AND symb_decoder(16#bf#)) OR
 					(reg_q2052 AND symb_decoder(16#ff#)) OR
 					(reg_q2052 AND symb_decoder(16#74#)) OR
 					(reg_q2052 AND symb_decoder(16#93#)) OR
 					(reg_q2052 AND symb_decoder(16#99#)) OR
 					(reg_q2052 AND symb_decoder(16#5a#)) OR
 					(reg_q2052 AND symb_decoder(16#72#)) OR
 					(reg_q2052 AND symb_decoder(16#80#)) OR
 					(reg_q2052 AND symb_decoder(16#67#)) OR
 					(reg_q2052 AND symb_decoder(16#e6#)) OR
 					(reg_q2052 AND symb_decoder(16#cc#)) OR
 					(reg_q2052 AND symb_decoder(16#e1#)) OR
 					(reg_q2052 AND symb_decoder(16#6d#)) OR
 					(reg_q2052 AND symb_decoder(16#a3#)) OR
 					(reg_q2052 AND symb_decoder(16#32#)) OR
 					(reg_q2052 AND symb_decoder(16#1b#)) OR
 					(reg_q2052 AND symb_decoder(16#85#)) OR
 					(reg_q2052 AND symb_decoder(16#2f#)) OR
 					(reg_q2052 AND symb_decoder(16#29#)) OR
 					(reg_q2052 AND symb_decoder(16#6c#)) OR
 					(reg_q2052 AND symb_decoder(16#21#)) OR
 					(reg_q2052 AND symb_decoder(16#38#)) OR
 					(reg_q2052 AND symb_decoder(16#92#)) OR
 					(reg_q2052 AND symb_decoder(16#b4#)) OR
 					(reg_q2052 AND symb_decoder(16#07#)) OR
 					(reg_q2052 AND symb_decoder(16#51#)) OR
 					(reg_q2052 AND symb_decoder(16#1f#)) OR
 					(reg_q2052 AND symb_decoder(16#7b#)) OR
 					(reg_q2052 AND symb_decoder(16#9a#)) OR
 					(reg_q2052 AND symb_decoder(16#5e#)) OR
 					(reg_q2052 AND symb_decoder(16#70#)) OR
 					(reg_q2052 AND symb_decoder(16#ad#)) OR
 					(reg_q2052 AND symb_decoder(16#b7#)) OR
 					(reg_q2052 AND symb_decoder(16#fc#)) OR
 					(reg_q2052 AND symb_decoder(16#6b#)) OR
 					(reg_q2052 AND symb_decoder(16#f5#)) OR
 					(reg_q2052 AND symb_decoder(16#7c#)) OR
 					(reg_q2052 AND symb_decoder(16#4e#)) OR
 					(reg_q2052 AND symb_decoder(16#9d#)) OR
 					(reg_q2052 AND symb_decoder(16#dc#)) OR
 					(reg_q2052 AND symb_decoder(16#17#)) OR
 					(reg_q2052 AND symb_decoder(16#30#)) OR
 					(reg_q2052 AND symb_decoder(16#db#)) OR
 					(reg_q2052 AND symb_decoder(16#ab#)) OR
 					(reg_q2052 AND symb_decoder(16#63#)) OR
 					(reg_q2052 AND symb_decoder(16#f3#)) OR
 					(reg_q2052 AND symb_decoder(16#11#)) OR
 					(reg_q2052 AND symb_decoder(16#1c#)) OR
 					(reg_q2052 AND symb_decoder(16#b2#)) OR
 					(reg_q2052 AND symb_decoder(16#fb#)) OR
 					(reg_q2052 AND symb_decoder(16#9e#)) OR
 					(reg_q2052 AND symb_decoder(16#d6#)) OR
 					(reg_q2052 AND symb_decoder(16#83#)) OR
 					(reg_q2052 AND symb_decoder(16#b6#)) OR
 					(reg_q2052 AND symb_decoder(16#28#)) OR
 					(reg_q2052 AND symb_decoder(16#55#)) OR
 					(reg_q2052 AND symb_decoder(16#f9#)) OR
 					(reg_q2052 AND symb_decoder(16#41#)) OR
 					(reg_q2052 AND symb_decoder(16#d1#)) OR
 					(reg_q2052 AND symb_decoder(16#4b#)) OR
 					(reg_q2052 AND symb_decoder(16#14#)) OR
 					(reg_q2052 AND symb_decoder(16#a9#)) OR
 					(reg_q2052 AND symb_decoder(16#3e#)) OR
 					(reg_q2052 AND symb_decoder(16#6a#)) OR
 					(reg_q2052 AND symb_decoder(16#d3#)) OR
 					(reg_q2052 AND symb_decoder(16#c0#)) OR
 					(reg_q2052 AND symb_decoder(16#69#)) OR
 					(reg_q2052 AND symb_decoder(16#16#)) OR
 					(reg_q2052 AND symb_decoder(16#22#)) OR
 					(reg_q2052 AND symb_decoder(16#c3#)) OR
 					(reg_q2052 AND symb_decoder(16#47#)) OR
 					(reg_q2052 AND symb_decoder(16#c6#)) OR
 					(reg_q2052 AND symb_decoder(16#3b#)) OR
 					(reg_q2052 AND symb_decoder(16#c4#)) OR
 					(reg_q2052 AND symb_decoder(16#c8#)) OR
 					(reg_q2052 AND symb_decoder(16#66#)) OR
 					(reg_q2052 AND symb_decoder(16#5f#)) OR
 					(reg_q2052 AND symb_decoder(16#e8#)) OR
 					(reg_q2052 AND symb_decoder(16#45#)) OR
 					(reg_q2052 AND symb_decoder(16#31#)) OR
 					(reg_q2052 AND symb_decoder(16#4f#)) OR
 					(reg_q2052 AND symb_decoder(16#73#)) OR
 					(reg_q2052 AND symb_decoder(16#e4#)) OR
 					(reg_q2052 AND symb_decoder(16#89#)) OR
 					(reg_q2052 AND symb_decoder(16#c7#)) OR
 					(reg_q2052 AND symb_decoder(16#f2#)) OR
 					(reg_q2052 AND symb_decoder(16#23#)) OR
 					(reg_q2052 AND symb_decoder(16#d5#)) OR
 					(reg_q2052 AND symb_decoder(16#58#)) OR
 					(reg_q2052 AND symb_decoder(16#98#));
reg_q2052_init <= '0' ;
	p_reg_q2052: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2052 <= reg_q2052_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2052 <= reg_q2052_init;
        else
          reg_q2052 <= reg_q2052_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q363_in <= (reg_q363 AND symb_decoder(16#0d#)) OR
 					(reg_q363 AND symb_decoder(16#20#)) OR
 					(reg_q363 AND symb_decoder(16#0a#)) OR
 					(reg_q363 AND symb_decoder(16#09#)) OR
 					(reg_q363 AND symb_decoder(16#0c#)) OR
 					(reg_q361 AND symb_decoder(16#20#)) OR
 					(reg_q361 AND symb_decoder(16#0c#)) OR
 					(reg_q361 AND symb_decoder(16#09#)) OR
 					(reg_q361 AND symb_decoder(16#0d#)) OR
 					(reg_q361 AND symb_decoder(16#0a#));
reg_q363_init <= '0' ;
	p_reg_q363: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q363 <= reg_q363_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q363 <= reg_q363_init;
        else
          reg_q363 <= reg_q363_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q365_in <= (reg_q363 AND symb_decoder(16#35#)) OR
 					(reg_q363 AND symb_decoder(16#34#)) OR
 					(reg_q363 AND symb_decoder(16#31#)) OR
 					(reg_q363 AND symb_decoder(16#32#)) OR
 					(reg_q363 AND symb_decoder(16#30#)) OR
 					(reg_q363 AND symb_decoder(16#39#)) OR
 					(reg_q363 AND symb_decoder(16#37#)) OR
 					(reg_q363 AND symb_decoder(16#33#)) OR
 					(reg_q363 AND symb_decoder(16#38#)) OR
 					(reg_q363 AND symb_decoder(16#36#)) OR
 					(reg_q365 AND symb_decoder(16#36#)) OR
 					(reg_q365 AND symb_decoder(16#35#)) OR
 					(reg_q365 AND symb_decoder(16#33#)) OR
 					(reg_q365 AND symb_decoder(16#30#)) OR
 					(reg_q365 AND symb_decoder(16#38#)) OR
 					(reg_q365 AND symb_decoder(16#34#)) OR
 					(reg_q365 AND symb_decoder(16#31#)) OR
 					(reg_q365 AND symb_decoder(16#32#)) OR
 					(reg_q365 AND symb_decoder(16#37#)) OR
 					(reg_q365 AND symb_decoder(16#39#));
reg_q365_init <= '0' ;
	p_reg_q365: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q365 <= reg_q365_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q365 <= reg_q365_init;
        else
          reg_q365 <= reg_q365_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1137_in <= (reg_q1137 AND symb_decoder(16#0d#)) OR
 					(reg_q1137 AND symb_decoder(16#20#)) OR
 					(reg_q1137 AND symb_decoder(16#0c#)) OR
 					(reg_q1137 AND symb_decoder(16#0a#)) OR
 					(reg_q1137 AND symb_decoder(16#09#)) OR
 					(reg_q1135 AND symb_decoder(16#09#)) OR
 					(reg_q1135 AND symb_decoder(16#0a#)) OR
 					(reg_q1135 AND symb_decoder(16#0c#)) OR
 					(reg_q1135 AND symb_decoder(16#20#)) OR
 					(reg_q1135 AND symb_decoder(16#0d#));
reg_q1137_init <= '0' ;
	p_reg_q1137: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1137 <= reg_q1137_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1137 <= reg_q1137_init;
        else
          reg_q1137 <= reg_q1137_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1139_in <= (reg_q1137 AND symb_decoder(16#31#)) OR
 					(reg_q1137 AND symb_decoder(16#33#)) OR
 					(reg_q1137 AND symb_decoder(16#37#)) OR
 					(reg_q1137 AND symb_decoder(16#34#)) OR
 					(reg_q1137 AND symb_decoder(16#39#)) OR
 					(reg_q1137 AND symb_decoder(16#35#)) OR
 					(reg_q1137 AND symb_decoder(16#30#)) OR
 					(reg_q1137 AND symb_decoder(16#32#)) OR
 					(reg_q1137 AND symb_decoder(16#36#)) OR
 					(reg_q1137 AND symb_decoder(16#38#)) OR
 					(reg_q1139 AND symb_decoder(16#36#)) OR
 					(reg_q1139 AND symb_decoder(16#34#)) OR
 					(reg_q1139 AND symb_decoder(16#37#)) OR
 					(reg_q1139 AND symb_decoder(16#33#)) OR
 					(reg_q1139 AND symb_decoder(16#35#)) OR
 					(reg_q1139 AND symb_decoder(16#31#)) OR
 					(reg_q1139 AND symb_decoder(16#30#)) OR
 					(reg_q1139 AND symb_decoder(16#38#)) OR
 					(reg_q1139 AND symb_decoder(16#39#)) OR
 					(reg_q1139 AND symb_decoder(16#32#));
reg_q1139_init <= '0' ;
	p_reg_q1139: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1139 <= reg_q1139_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1139 <= reg_q1139_init;
        else
          reg_q1139 <= reg_q1139_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q696_in <= (reg_q696 AND symb_decoder(16#32#)) OR
 					(reg_q696 AND symb_decoder(16#35#)) OR
 					(reg_q696 AND symb_decoder(16#38#)) OR
 					(reg_q696 AND symb_decoder(16#30#)) OR
 					(reg_q696 AND symb_decoder(16#33#)) OR
 					(reg_q696 AND symb_decoder(16#31#)) OR
 					(reg_q696 AND symb_decoder(16#34#)) OR
 					(reg_q696 AND symb_decoder(16#37#)) OR
 					(reg_q696 AND symb_decoder(16#39#)) OR
 					(reg_q696 AND symb_decoder(16#36#)) OR
 					(reg_q694 AND symb_decoder(16#38#)) OR
 					(reg_q694 AND symb_decoder(16#32#)) OR
 					(reg_q694 AND symb_decoder(16#33#)) OR
 					(reg_q694 AND symb_decoder(16#35#)) OR
 					(reg_q694 AND symb_decoder(16#36#)) OR
 					(reg_q694 AND symb_decoder(16#34#)) OR
 					(reg_q694 AND symb_decoder(16#39#)) OR
 					(reg_q694 AND symb_decoder(16#30#)) OR
 					(reg_q694 AND symb_decoder(16#31#)) OR
 					(reg_q694 AND symb_decoder(16#37#));
reg_q696_init <= '0' ;
	p_reg_q696: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q696 <= reg_q696_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q696 <= reg_q696_init;
        else
          reg_q696 <= reg_q696_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q698_in <= (reg_q696 AND symb_decoder(16#2e#));
reg_q698_init <= '0' ;
	p_reg_q698: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q698 <= reg_q698_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q698 <= reg_q698_init;
        else
          reg_q698 <= reg_q698_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q472_in <= (reg_q470 AND symb_decoder(16#25#));
reg_q472_init <= '0' ;
	p_reg_q472: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q472 <= reg_q472_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q472 <= reg_q472_init;
        else
          reg_q472 <= reg_q472_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q474_in <= (reg_q472 AND symb_decoder(16#32#));
reg_q474_init <= '0' ;
	p_reg_q474: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q474 <= reg_q474_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q474 <= reg_q474_init;
        else
          reg_q474 <= reg_q474_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1816_in <= (reg_q1814 AND symb_decoder(16#0d#)) OR
 					(reg_q1814 AND symb_decoder(16#09#)) OR
 					(reg_q1814 AND symb_decoder(16#0a#)) OR
 					(reg_q1814 AND symb_decoder(16#0c#)) OR
 					(reg_q1814 AND symb_decoder(16#20#)) OR
 					(reg_q1816 AND symb_decoder(16#09#)) OR
 					(reg_q1816 AND symb_decoder(16#0c#)) OR
 					(reg_q1816 AND symb_decoder(16#0a#)) OR
 					(reg_q1816 AND symb_decoder(16#20#)) OR
 					(reg_q1816 AND symb_decoder(16#0d#));
reg_q1816_init <= '0' ;
	p_reg_q1816: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1816 <= reg_q1816_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1816 <= reg_q1816_init;
        else
          reg_q1816 <= reg_q1816_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1818_in <= (reg_q1816 AND symb_decoder(16#76#)) OR
 					(reg_q1816 AND symb_decoder(16#56#));
reg_q1818_init <= '0' ;
	p_reg_q1818: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1818 <= reg_q1818_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1818 <= reg_q1818_init;
        else
          reg_q1818 <= reg_q1818_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1975_in <= (reg_q1973 AND symb_decoder(16#23#));
reg_q1975_init <= '0' ;
	p_reg_q1975: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1975 <= reg_q1975_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1975 <= reg_q1975_init;
        else
          reg_q1975 <= reg_q1975_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q46_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q46 AND symb_decoder(16#56#)) OR
 					(reg_q46 AND symb_decoder(16#04#)) OR
 					(reg_q46 AND symb_decoder(16#f5#)) OR
 					(reg_q46 AND symb_decoder(16#ce#)) OR
 					(reg_q46 AND symb_decoder(16#58#)) OR
 					(reg_q46 AND symb_decoder(16#93#)) OR
 					(reg_q46 AND symb_decoder(16#46#)) OR
 					(reg_q46 AND symb_decoder(16#1a#)) OR
 					(reg_q46 AND symb_decoder(16#34#)) OR
 					(reg_q46 AND symb_decoder(16#32#)) OR
 					(reg_q46 AND symb_decoder(16#e0#)) OR
 					(reg_q46 AND symb_decoder(16#16#)) OR
 					(reg_q46 AND symb_decoder(16#64#)) OR
 					(reg_q46 AND symb_decoder(16#cc#)) OR
 					(reg_q46 AND symb_decoder(16#4d#)) OR
 					(reg_q46 AND symb_decoder(16#72#)) OR
 					(reg_q46 AND symb_decoder(16#1e#)) OR
 					(reg_q46 AND symb_decoder(16#db#)) OR
 					(reg_q46 AND symb_decoder(16#35#)) OR
 					(reg_q46 AND symb_decoder(16#38#)) OR
 					(reg_q46 AND symb_decoder(16#0d#)) OR
 					(reg_q46 AND symb_decoder(16#bc#)) OR
 					(reg_q46 AND symb_decoder(16#84#)) OR
 					(reg_q46 AND symb_decoder(16#2b#)) OR
 					(reg_q46 AND symb_decoder(16#c9#)) OR
 					(reg_q46 AND symb_decoder(16#74#)) OR
 					(reg_q46 AND symb_decoder(16#b6#)) OR
 					(reg_q46 AND symb_decoder(16#4a#)) OR
 					(reg_q46 AND symb_decoder(16#e8#)) OR
 					(reg_q46 AND symb_decoder(16#2a#)) OR
 					(reg_q46 AND symb_decoder(16#03#)) OR
 					(reg_q46 AND symb_decoder(16#6b#)) OR
 					(reg_q46 AND symb_decoder(16#f8#)) OR
 					(reg_q46 AND symb_decoder(16#20#)) OR
 					(reg_q46 AND symb_decoder(16#11#)) OR
 					(reg_q46 AND symb_decoder(16#51#)) OR
 					(reg_q46 AND symb_decoder(16#54#)) OR
 					(reg_q46 AND symb_decoder(16#60#)) OR
 					(reg_q46 AND symb_decoder(16#25#)) OR
 					(reg_q46 AND symb_decoder(16#28#)) OR
 					(reg_q46 AND symb_decoder(16#dd#)) OR
 					(reg_q46 AND symb_decoder(16#07#)) OR
 					(reg_q46 AND symb_decoder(16#d7#)) OR
 					(reg_q46 AND symb_decoder(16#5d#)) OR
 					(reg_q46 AND symb_decoder(16#2e#)) OR
 					(reg_q46 AND symb_decoder(16#86#)) OR
 					(reg_q46 AND symb_decoder(16#9e#)) OR
 					(reg_q46 AND symb_decoder(16#a3#)) OR
 					(reg_q46 AND symb_decoder(16#9d#)) OR
 					(reg_q46 AND symb_decoder(16#3b#)) OR
 					(reg_q46 AND symb_decoder(16#2c#)) OR
 					(reg_q46 AND symb_decoder(16#a7#)) OR
 					(reg_q46 AND symb_decoder(16#e1#)) OR
 					(reg_q46 AND symb_decoder(16#4f#)) OR
 					(reg_q46 AND symb_decoder(16#d5#)) OR
 					(reg_q46 AND symb_decoder(16#c4#)) OR
 					(reg_q46 AND symb_decoder(16#7b#)) OR
 					(reg_q46 AND symb_decoder(16#62#)) OR
 					(reg_q46 AND symb_decoder(16#99#)) OR
 					(reg_q46 AND symb_decoder(16#61#)) OR
 					(reg_q46 AND symb_decoder(16#6d#)) OR
 					(reg_q46 AND symb_decoder(16#7d#)) OR
 					(reg_q46 AND symb_decoder(16#dc#)) OR
 					(reg_q46 AND symb_decoder(16#1c#)) OR
 					(reg_q46 AND symb_decoder(16#cd#)) OR
 					(reg_q46 AND symb_decoder(16#f3#)) OR
 					(reg_q46 AND symb_decoder(16#fa#)) OR
 					(reg_q46 AND symb_decoder(16#42#)) OR
 					(reg_q46 AND symb_decoder(16#88#)) OR
 					(reg_q46 AND symb_decoder(16#9b#)) OR
 					(reg_q46 AND symb_decoder(16#44#)) OR
 					(reg_q46 AND symb_decoder(16#52#)) OR
 					(reg_q46 AND symb_decoder(16#f0#)) OR
 					(reg_q46 AND symb_decoder(16#f1#)) OR
 					(reg_q46 AND symb_decoder(16#96#)) OR
 					(reg_q46 AND symb_decoder(16#0b#)) OR
 					(reg_q46 AND symb_decoder(16#f6#)) OR
 					(reg_q46 AND symb_decoder(16#cf#)) OR
 					(reg_q46 AND symb_decoder(16#8e#)) OR
 					(reg_q46 AND symb_decoder(16#79#)) OR
 					(reg_q46 AND symb_decoder(16#67#)) OR
 					(reg_q46 AND symb_decoder(16#ac#)) OR
 					(reg_q46 AND symb_decoder(16#e7#)) OR
 					(reg_q46 AND symb_decoder(16#94#)) OR
 					(reg_q46 AND symb_decoder(16#a9#)) OR
 					(reg_q46 AND symb_decoder(16#b4#)) OR
 					(reg_q46 AND symb_decoder(16#36#)) OR
 					(reg_q46 AND symb_decoder(16#3f#)) OR
 					(reg_q46 AND symb_decoder(16#37#)) OR
 					(reg_q46 AND symb_decoder(16#26#)) OR
 					(reg_q46 AND symb_decoder(16#22#)) OR
 					(reg_q46 AND symb_decoder(16#b3#)) OR
 					(reg_q46 AND symb_decoder(16#4c#)) OR
 					(reg_q46 AND symb_decoder(16#fb#)) OR
 					(reg_q46 AND symb_decoder(16#2f#)) OR
 					(reg_q46 AND symb_decoder(16#4b#)) OR
 					(reg_q46 AND symb_decoder(16#33#)) OR
 					(reg_q46 AND symb_decoder(16#a1#)) OR
 					(reg_q46 AND symb_decoder(16#2d#)) OR
 					(reg_q46 AND symb_decoder(16#b5#)) OR
 					(reg_q46 AND symb_decoder(16#12#)) OR
 					(reg_q46 AND symb_decoder(16#6f#)) OR
 					(reg_q46 AND symb_decoder(16#a4#)) OR
 					(reg_q46 AND symb_decoder(16#eb#)) OR
 					(reg_q46 AND symb_decoder(16#90#)) OR
 					(reg_q46 AND symb_decoder(16#ee#)) OR
 					(reg_q46 AND symb_decoder(16#69#)) OR
 					(reg_q46 AND symb_decoder(16#4e#)) OR
 					(reg_q46 AND symb_decoder(16#f2#)) OR
 					(reg_q46 AND symb_decoder(16#b7#)) OR
 					(reg_q46 AND symb_decoder(16#d3#)) OR
 					(reg_q46 AND symb_decoder(16#a6#)) OR
 					(reg_q46 AND symb_decoder(16#ec#)) OR
 					(reg_q46 AND symb_decoder(16#e9#)) OR
 					(reg_q46 AND symb_decoder(16#43#)) OR
 					(reg_q46 AND symb_decoder(16#14#)) OR
 					(reg_q46 AND symb_decoder(16#da#)) OR
 					(reg_q46 AND symb_decoder(16#13#)) OR
 					(reg_q46 AND symb_decoder(16#d2#)) OR
 					(reg_q46 AND symb_decoder(16#18#)) OR
 					(reg_q46 AND symb_decoder(16#41#)) OR
 					(reg_q46 AND symb_decoder(16#d1#)) OR
 					(reg_q46 AND symb_decoder(16#70#)) OR
 					(reg_q46 AND symb_decoder(16#31#)) OR
 					(reg_q46 AND symb_decoder(16#30#)) OR
 					(reg_q46 AND symb_decoder(16#06#)) OR
 					(reg_q46 AND symb_decoder(16#48#)) OR
 					(reg_q46 AND symb_decoder(16#ff#)) OR
 					(reg_q46 AND symb_decoder(16#53#)) OR
 					(reg_q46 AND symb_decoder(16#7a#)) OR
 					(reg_q46 AND symb_decoder(16#b1#)) OR
 					(reg_q46 AND symb_decoder(16#85#)) OR
 					(reg_q46 AND symb_decoder(16#24#)) OR
 					(reg_q46 AND symb_decoder(16#57#)) OR
 					(reg_q46 AND symb_decoder(16#23#)) OR
 					(reg_q46 AND symb_decoder(16#b8#)) OR
 					(reg_q46 AND symb_decoder(16#59#)) OR
 					(reg_q46 AND symb_decoder(16#6c#)) OR
 					(reg_q46 AND symb_decoder(16#d9#)) OR
 					(reg_q46 AND symb_decoder(16#08#)) OR
 					(reg_q46 AND symb_decoder(16#09#)) OR
 					(reg_q46 AND symb_decoder(16#6e#)) OR
 					(reg_q46 AND symb_decoder(16#bf#)) OR
 					(reg_q46 AND symb_decoder(16#49#)) OR
 					(reg_q46 AND symb_decoder(16#21#)) OR
 					(reg_q46 AND symb_decoder(16#75#)) OR
 					(reg_q46 AND symb_decoder(16#c2#)) OR
 					(reg_q46 AND symb_decoder(16#8d#)) OR
 					(reg_q46 AND symb_decoder(16#d4#)) OR
 					(reg_q46 AND symb_decoder(16#d6#)) OR
 					(reg_q46 AND symb_decoder(16#3d#)) OR
 					(reg_q46 AND symb_decoder(16#c5#)) OR
 					(reg_q46 AND symb_decoder(16#e4#)) OR
 					(reg_q46 AND symb_decoder(16#55#)) OR
 					(reg_q46 AND symb_decoder(16#98#)) OR
 					(reg_q46 AND symb_decoder(16#3c#)) OR
 					(reg_q46 AND symb_decoder(16#aa#)) OR
 					(reg_q46 AND symb_decoder(16#05#)) OR
 					(reg_q46 AND symb_decoder(16#27#)) OR
 					(reg_q46 AND symb_decoder(16#fd#)) OR
 					(reg_q46 AND symb_decoder(16#29#)) OR
 					(reg_q46 AND symb_decoder(16#fe#)) OR
 					(reg_q46 AND symb_decoder(16#b0#)) OR
 					(reg_q46 AND symb_decoder(16#0a#)) OR
 					(reg_q46 AND symb_decoder(16#0c#)) OR
 					(reg_q46 AND symb_decoder(16#e3#)) OR
 					(reg_q46 AND symb_decoder(16#8c#)) OR
 					(reg_q46 AND symb_decoder(16#73#)) OR
 					(reg_q46 AND symb_decoder(16#8a#)) OR
 					(reg_q46 AND symb_decoder(16#ed#)) OR
 					(reg_q46 AND symb_decoder(16#89#)) OR
 					(reg_q46 AND symb_decoder(16#81#)) OR
 					(reg_q46 AND symb_decoder(16#80#)) OR
 					(reg_q46 AND symb_decoder(16#ad#)) OR
 					(reg_q46 AND symb_decoder(16#ab#)) OR
 					(reg_q46 AND symb_decoder(16#7c#)) OR
 					(reg_q46 AND symb_decoder(16#5e#)) OR
 					(reg_q46 AND symb_decoder(16#9a#)) OR
 					(reg_q46 AND symb_decoder(16#d0#)) OR
 					(reg_q46 AND symb_decoder(16#1b#)) OR
 					(reg_q46 AND symb_decoder(16#87#)) OR
 					(reg_q46 AND symb_decoder(16#b9#)) OR
 					(reg_q46 AND symb_decoder(16#cb#)) OR
 					(reg_q46 AND symb_decoder(16#ae#)) OR
 					(reg_q46 AND symb_decoder(16#02#)) OR
 					(reg_q46 AND symb_decoder(16#40#)) OR
 					(reg_q46 AND symb_decoder(16#de#)) OR
 					(reg_q46 AND symb_decoder(16#c7#)) OR
 					(reg_q46 AND symb_decoder(16#45#)) OR
 					(reg_q46 AND symb_decoder(16#ea#)) OR
 					(reg_q46 AND symb_decoder(16#92#)) OR
 					(reg_q46 AND symb_decoder(16#ca#)) OR
 					(reg_q46 AND symb_decoder(16#95#)) OR
 					(reg_q46 AND symb_decoder(16#3a#)) OR
 					(reg_q46 AND symb_decoder(16#ef#)) OR
 					(reg_q46 AND symb_decoder(16#e5#)) OR
 					(reg_q46 AND symb_decoder(16#6a#)) OR
 					(reg_q46 AND symb_decoder(16#66#)) OR
 					(reg_q46 AND symb_decoder(16#47#)) OR
 					(reg_q46 AND symb_decoder(16#00#)) OR
 					(reg_q46 AND symb_decoder(16#19#)) OR
 					(reg_q46 AND symb_decoder(16#f9#)) OR
 					(reg_q46 AND symb_decoder(16#17#)) OR
 					(reg_q46 AND symb_decoder(16#c0#)) OR
 					(reg_q46 AND symb_decoder(16#c8#)) OR
 					(reg_q46 AND symb_decoder(16#a0#)) OR
 					(reg_q46 AND symb_decoder(16#bb#)) OR
 					(reg_q46 AND symb_decoder(16#9f#)) OR
 					(reg_q46 AND symb_decoder(16#83#)) OR
 					(reg_q46 AND symb_decoder(16#97#)) OR
 					(reg_q46 AND symb_decoder(16#af#)) OR
 					(reg_q46 AND symb_decoder(16#76#)) OR
 					(reg_q46 AND symb_decoder(16#82#)) OR
 					(reg_q46 AND symb_decoder(16#a5#)) OR
 					(reg_q46 AND symb_decoder(16#c6#)) OR
 					(reg_q46 AND symb_decoder(16#10#)) OR
 					(reg_q46 AND symb_decoder(16#f7#)) OR
 					(reg_q46 AND symb_decoder(16#a8#)) OR
 					(reg_q46 AND symb_decoder(16#91#)) OR
 					(reg_q46 AND symb_decoder(16#39#)) OR
 					(reg_q46 AND symb_decoder(16#a2#)) OR
 					(reg_q46 AND symb_decoder(16#5c#)) OR
 					(reg_q46 AND symb_decoder(16#3e#)) OR
 					(reg_q46 AND symb_decoder(16#78#)) OR
 					(reg_q46 AND symb_decoder(16#68#)) OR
 					(reg_q46 AND symb_decoder(16#ba#)) OR
 					(reg_q46 AND symb_decoder(16#9c#)) OR
 					(reg_q46 AND symb_decoder(16#c1#)) OR
 					(reg_q46 AND symb_decoder(16#7e#)) OR
 					(reg_q46 AND symb_decoder(16#65#)) OR
 					(reg_q46 AND symb_decoder(16#0e#)) OR
 					(reg_q46 AND symb_decoder(16#bd#)) OR
 					(reg_q46 AND symb_decoder(16#8b#)) OR
 					(reg_q46 AND symb_decoder(16#5f#)) OR
 					(reg_q46 AND symb_decoder(16#01#)) OR
 					(reg_q46 AND symb_decoder(16#b2#)) OR
 					(reg_q46 AND symb_decoder(16#7f#)) OR
 					(reg_q46 AND symb_decoder(16#8f#)) OR
 					(reg_q46 AND symb_decoder(16#5a#)) OR
 					(reg_q46 AND symb_decoder(16#f4#)) OR
 					(reg_q46 AND symb_decoder(16#be#)) OR
 					(reg_q46 AND symb_decoder(16#df#)) OR
 					(reg_q46 AND symb_decoder(16#50#)) OR
 					(reg_q46 AND symb_decoder(16#1d#)) OR
 					(reg_q46 AND symb_decoder(16#c3#)) OR
 					(reg_q46 AND symb_decoder(16#d8#)) OR
 					(reg_q46 AND symb_decoder(16#fc#)) OR
 					(reg_q46 AND symb_decoder(16#1f#)) OR
 					(reg_q46 AND symb_decoder(16#e6#)) OR
 					(reg_q46 AND symb_decoder(16#5b#)) OR
 					(reg_q46 AND symb_decoder(16#71#)) OR
 					(reg_q46 AND symb_decoder(16#15#)) OR
 					(reg_q46 AND symb_decoder(16#63#)) OR
 					(reg_q46 AND symb_decoder(16#0f#)) OR
 					(reg_q46 AND symb_decoder(16#e2#)) OR
 					(reg_q46 AND symb_decoder(16#77#));
reg_q46_init <= '0' ;
	p_reg_q46: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q46 <= reg_q46_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q46 <= reg_q46_init;
        else
          reg_q46 <= reg_q46_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2461_in <= (reg_q2459 AND symb_decoder(16#23#));
reg_q2461_init <= '0' ;
	p_reg_q2461: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2461 <= reg_q2461_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2461 <= reg_q2461_init;
        else
          reg_q2461 <= reg_q2461_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2463_in <= (reg_q2461 AND symb_decoder(16#46#)) OR
 					(reg_q2461 AND symb_decoder(16#66#));
reg_q2463_init <= '0' ;
	p_reg_q2463: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2463 <= reg_q2463_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2463 <= reg_q2463_init;
        else
          reg_q2463 <= reg_q2463_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q700_in <= (reg_q698 AND symb_decoder(16#34#)) OR
 					(reg_q698 AND symb_decoder(16#38#)) OR
 					(reg_q698 AND symb_decoder(16#37#)) OR
 					(reg_q698 AND symb_decoder(16#35#)) OR
 					(reg_q698 AND symb_decoder(16#39#)) OR
 					(reg_q698 AND symb_decoder(16#36#)) OR
 					(reg_q698 AND symb_decoder(16#31#)) OR
 					(reg_q698 AND symb_decoder(16#33#)) OR
 					(reg_q698 AND symb_decoder(16#30#)) OR
 					(reg_q698 AND symb_decoder(16#32#)) OR
 					(reg_q700 AND symb_decoder(16#38#)) OR
 					(reg_q700 AND symb_decoder(16#30#)) OR
 					(reg_q700 AND symb_decoder(16#34#)) OR
 					(reg_q700 AND symb_decoder(16#39#)) OR
 					(reg_q700 AND symb_decoder(16#37#)) OR
 					(reg_q700 AND symb_decoder(16#35#)) OR
 					(reg_q700 AND symb_decoder(16#32#)) OR
 					(reg_q700 AND symb_decoder(16#33#)) OR
 					(reg_q700 AND symb_decoder(16#36#)) OR
 					(reg_q700 AND symb_decoder(16#31#));
reg_q700_init <= '0' ;
	p_reg_q700: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q700 <= reg_q700_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q700 <= reg_q700_init;
        else
          reg_q700 <= reg_q700_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q58_in <= (reg_q58 AND symb_decoder(16#0c#)) OR
 					(reg_q58 AND symb_decoder(16#0a#)) OR
 					(reg_q58 AND symb_decoder(16#09#)) OR
 					(reg_q58 AND symb_decoder(16#0d#)) OR
 					(reg_q58 AND symb_decoder(16#20#)) OR
 					(reg_q56 AND symb_decoder(16#09#)) OR
 					(reg_q56 AND symb_decoder(16#20#)) OR
 					(reg_q56 AND symb_decoder(16#0a#)) OR
 					(reg_q56 AND symb_decoder(16#0d#)) OR
 					(reg_q56 AND symb_decoder(16#0c#));
reg_q58_init <= '0' ;
	p_reg_q58: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q58 <= reg_q58_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q58 <= reg_q58_init;
        else
          reg_q58 <= reg_q58_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2030_in <= (reg_q2030 AND symb_decoder(16#20#)) OR
 					(reg_q2030 AND symb_decoder(16#09#)) OR
 					(reg_q2030 AND symb_decoder(16#0a#)) OR
 					(reg_q2030 AND symb_decoder(16#0c#)) OR
 					(reg_q2030 AND symb_decoder(16#0d#)) OR
 					(reg_q2028 AND symb_decoder(16#0d#)) OR
 					(reg_q2028 AND symb_decoder(16#09#)) OR
 					(reg_q2028 AND symb_decoder(16#0c#)) OR
 					(reg_q2028 AND symb_decoder(16#0a#)) OR
 					(reg_q2028 AND symb_decoder(16#20#));
reg_q2030_init <= '0' ;
	p_reg_q2030: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2030 <= reg_q2030_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2030 <= reg_q2030_init;
        else
          reg_q2030 <= reg_q2030_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2032_in <= (reg_q2030 AND symb_decoder(16#66#)) OR
 					(reg_q2030 AND symb_decoder(16#46#));
reg_q2032_init <= '0' ;
	p_reg_q2032: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2032 <= reg_q2032_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2032 <= reg_q2032_init;
        else
          reg_q2032 <= reg_q2032_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1926_in <= (reg_q1926 AND symb_decoder(16#0a#)) OR
 					(reg_q1926 AND symb_decoder(16#09#)) OR
 					(reg_q1926 AND symb_decoder(16#0d#)) OR
 					(reg_q1926 AND symb_decoder(16#20#)) OR
 					(reg_q1926 AND symb_decoder(16#0c#)) OR
 					(reg_q1924 AND symb_decoder(16#09#)) OR
 					(reg_q1924 AND symb_decoder(16#0a#)) OR
 					(reg_q1924 AND symb_decoder(16#20#)) OR
 					(reg_q1924 AND symb_decoder(16#0d#)) OR
 					(reg_q1924 AND symb_decoder(16#0c#));
reg_q1926_init <= '0' ;
	p_reg_q1926: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1926 <= reg_q1926_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1926 <= reg_q1926_init;
        else
          reg_q1926 <= reg_q1926_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1246_in <= (reg_q1244 AND symb_decoder(16#72#)) OR
 					(reg_q1244 AND symb_decoder(16#52#));
reg_q1246_init <= '0' ;
	p_reg_q1246: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1246 <= reg_q1246_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1246 <= reg_q1246_init;
        else
          reg_q1246 <= reg_q1246_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1248_in <= (reg_q1246 AND symb_decoder(16#0c#)) OR
 					(reg_q1246 AND symb_decoder(16#20#)) OR
 					(reg_q1246 AND symb_decoder(16#09#)) OR
 					(reg_q1246 AND symb_decoder(16#0d#)) OR
 					(reg_q1246 AND symb_decoder(16#0a#)) OR
 					(reg_q1248 AND symb_decoder(16#0c#)) OR
 					(reg_q1248 AND symb_decoder(16#0a#)) OR
 					(reg_q1248 AND symb_decoder(16#0d#)) OR
 					(reg_q1248 AND symb_decoder(16#09#)) OR
 					(reg_q1248 AND symb_decoder(16#20#));
reg_q1248_init <= '0' ;
	p_reg_q1248: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1248 <= reg_q1248_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1248 <= reg_q1248_init;
        else
          reg_q1248 <= reg_q1248_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q616_in <= (reg_q616 AND symb_decoder(16#38#)) OR
 					(reg_q616 AND symb_decoder(16#32#)) OR
 					(reg_q616 AND symb_decoder(16#33#)) OR
 					(reg_q616 AND symb_decoder(16#35#)) OR
 					(reg_q616 AND symb_decoder(16#30#)) OR
 					(reg_q616 AND symb_decoder(16#36#)) OR
 					(reg_q616 AND symb_decoder(16#39#)) OR
 					(reg_q616 AND symb_decoder(16#31#)) OR
 					(reg_q616 AND symb_decoder(16#37#)) OR
 					(reg_q616 AND symb_decoder(16#34#)) OR
 					(reg_q614 AND symb_decoder(16#36#)) OR
 					(reg_q614 AND symb_decoder(16#35#)) OR
 					(reg_q614 AND symb_decoder(16#32#)) OR
 					(reg_q614 AND symb_decoder(16#30#)) OR
 					(reg_q614 AND symb_decoder(16#38#)) OR
 					(reg_q614 AND symb_decoder(16#37#)) OR
 					(reg_q614 AND symb_decoder(16#34#)) OR
 					(reg_q614 AND symb_decoder(16#39#)) OR
 					(reg_q614 AND symb_decoder(16#33#)) OR
 					(reg_q614 AND symb_decoder(16#31#));
reg_q616_init <= '0' ;
	p_reg_q616: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q616 <= reg_q616_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q616 <= reg_q616_init;
        else
          reg_q616 <= reg_q616_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2411_in <= (reg_q2411 AND symb_decoder(16#09#)) OR
 					(reg_q2411 AND symb_decoder(16#0c#)) OR
 					(reg_q2411 AND symb_decoder(16#0a#)) OR
 					(reg_q2411 AND symb_decoder(16#20#)) OR
 					(reg_q2411 AND symb_decoder(16#0d#)) OR
 					(reg_q2409 AND symb_decoder(16#20#)) OR
 					(reg_q2409 AND symb_decoder(16#0c#)) OR
 					(reg_q2409 AND symb_decoder(16#09#)) OR
 					(reg_q2409 AND symb_decoder(16#0d#)) OR
 					(reg_q2409 AND symb_decoder(16#0a#));
reg_q2411_init <= '0' ;
	p_reg_q2411: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2411 <= reg_q2411_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2411 <= reg_q2411_init;
        else
          reg_q2411 <= reg_q2411_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1770_in <= (reg_q1768 AND symb_decoder(16#09#)) OR
 					(reg_q1768 AND symb_decoder(16#0d#)) OR
 					(reg_q1768 AND symb_decoder(16#0c#)) OR
 					(reg_q1768 AND symb_decoder(16#0a#)) OR
 					(reg_q1768 AND symb_decoder(16#20#));
reg_q1770_init <= '0' ;
	p_reg_q1770: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1770 <= reg_q1770_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1770 <= reg_q1770_init;
        else
          reg_q1770 <= reg_q1770_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1772_in <= (reg_q1770 AND symb_decoder(16#0d#)) OR
 					(reg_q1770 AND symb_decoder(16#0c#)) OR
 					(reg_q1770 AND symb_decoder(16#09#)) OR
 					(reg_q1770 AND symb_decoder(16#0a#)) OR
 					(reg_q1770 AND symb_decoder(16#20#));
reg_q1772_init <= '0' ;
	p_reg_q1772: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1772 <= reg_q1772_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1772 <= reg_q1772_init;
        else
          reg_q1772 <= reg_q1772_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q520_in <= (reg_q518 AND symb_decoder(16#5f#));
reg_q520_init <= '0' ;
	p_reg_q520: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q520 <= reg_q520_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q520 <= reg_q520_init;
        else
          reg_q520 <= reg_q520_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q522_in <= (reg_q520 AND symb_decoder(16#31#)) OR
 					(reg_q520 AND symb_decoder(16#39#)) OR
 					(reg_q520 AND symb_decoder(16#32#)) OR
 					(reg_q520 AND symb_decoder(16#36#)) OR
 					(reg_q520 AND symb_decoder(16#38#)) OR
 					(reg_q520 AND symb_decoder(16#30#)) OR
 					(reg_q520 AND symb_decoder(16#34#)) OR
 					(reg_q520 AND symb_decoder(16#35#)) OR
 					(reg_q520 AND symb_decoder(16#37#)) OR
 					(reg_q520 AND symb_decoder(16#33#)) OR
 					(reg_q522 AND symb_decoder(16#36#)) OR
 					(reg_q522 AND symb_decoder(16#33#)) OR
 					(reg_q522 AND symb_decoder(16#39#)) OR
 					(reg_q522 AND symb_decoder(16#34#)) OR
 					(reg_q522 AND symb_decoder(16#30#)) OR
 					(reg_q522 AND symb_decoder(16#38#)) OR
 					(reg_q522 AND symb_decoder(16#31#)) OR
 					(reg_q522 AND symb_decoder(16#37#)) OR
 					(reg_q522 AND symb_decoder(16#32#)) OR
 					(reg_q522 AND symb_decoder(16#35#));
reg_q522_init <= '0' ;
	p_reg_q522: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q522 <= reg_q522_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q522 <= reg_q522_init;
        else
          reg_q522 <= reg_q522_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2103_in <= (reg_q2103 AND symb_decoder(16#0a#)) OR
 					(reg_q2103 AND symb_decoder(16#09#)) OR
 					(reg_q2103 AND symb_decoder(16#0c#)) OR
 					(reg_q2103 AND symb_decoder(16#0d#)) OR
 					(reg_q2103 AND symb_decoder(16#20#)) OR
 					(reg_q2101 AND symb_decoder(16#09#)) OR
 					(reg_q2101 AND symb_decoder(16#0d#)) OR
 					(reg_q2101 AND symb_decoder(16#20#)) OR
 					(reg_q2101 AND symb_decoder(16#0c#)) OR
 					(reg_q2101 AND symb_decoder(16#0a#));
reg_q2103_init <= '0' ;
	p_reg_q2103: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2103 <= reg_q2103_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2103 <= reg_q2103_init;
        else
          reg_q2103 <= reg_q2103_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2105_in <= (reg_q2103 AND symb_decoder(16#58#)) OR
 					(reg_q2103 AND symb_decoder(16#78#));
reg_q2105_init <= '0' ;
	p_reg_q2105: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2105 <= reg_q2105_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2105 <= reg_q2105_init;
        else
          reg_q2105 <= reg_q2105_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2300_in <= (reg_q2298 AND symb_decoder(16#72#)) OR
 					(reg_q2298 AND symb_decoder(16#52#));
reg_q2300_init <= '0' ;
	p_reg_q2300: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2300 <= reg_q2300_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2300 <= reg_q2300_init;
        else
          reg_q2300 <= reg_q2300_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2302_in <= (reg_q2300 AND symb_decoder(16#09#)) OR
 					(reg_q2300 AND symb_decoder(16#0d#)) OR
 					(reg_q2300 AND symb_decoder(16#20#)) OR
 					(reg_q2300 AND symb_decoder(16#0c#)) OR
 					(reg_q2300 AND symb_decoder(16#0a#)) OR
 					(reg_q2302 AND symb_decoder(16#09#)) OR
 					(reg_q2302 AND symb_decoder(16#0c#)) OR
 					(reg_q2302 AND symb_decoder(16#0a#)) OR
 					(reg_q2302 AND symb_decoder(16#20#)) OR
 					(reg_q2302 AND symb_decoder(16#0d#));
reg_q2302_init <= '0' ;
	p_reg_q2302: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2302 <= reg_q2302_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2302 <= reg_q2302_init;
        else
          reg_q2302 <= reg_q2302_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2130_in <= (reg_q2130 AND symb_decoder(16#09#)) OR
 					(reg_q2130 AND symb_decoder(16#20#)) OR
 					(reg_q2130 AND symb_decoder(16#0c#)) OR
 					(reg_q2130 AND symb_decoder(16#0d#)) OR
 					(reg_q2130 AND symb_decoder(16#0a#)) OR
 					(reg_q2128 AND symb_decoder(16#0d#)) OR
 					(reg_q2128 AND symb_decoder(16#09#)) OR
 					(reg_q2128 AND symb_decoder(16#0c#)) OR
 					(reg_q2128 AND symb_decoder(16#20#)) OR
 					(reg_q2128 AND symb_decoder(16#0a#));
reg_q2130_init <= '0' ;
	p_reg_q2130: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2130 <= reg_q2130_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2130 <= reg_q2130_init;
        else
          reg_q2130 <= reg_q2130_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q22_in <= (reg_q22 AND symb_decoder(16#09#)) OR
 					(reg_q22 AND symb_decoder(16#0c#)) OR
 					(reg_q22 AND symb_decoder(16#0d#)) OR
 					(reg_q22 AND symb_decoder(16#20#)) OR
 					(reg_q22 AND symb_decoder(16#0a#)) OR
 					(reg_q20 AND symb_decoder(16#20#)) OR
 					(reg_q20 AND symb_decoder(16#0c#)) OR
 					(reg_q20 AND symb_decoder(16#09#)) OR
 					(reg_q20 AND symb_decoder(16#0a#)) OR
 					(reg_q20 AND symb_decoder(16#0d#));
reg_q22_init <= '0' ;
	p_reg_q22: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q22 <= reg_q22_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q22 <= reg_q22_init;
        else
          reg_q22 <= reg_q22_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2579_in <= (reg_q2579 AND symb_decoder(16#20#)) OR
 					(reg_q2579 AND symb_decoder(16#0d#)) OR
 					(reg_q2579 AND symb_decoder(16#09#)) OR
 					(reg_q2579 AND symb_decoder(16#0c#)) OR
 					(reg_q2579 AND symb_decoder(16#0a#)) OR
 					(reg_q2577 AND symb_decoder(16#0c#)) OR
 					(reg_q2577 AND symb_decoder(16#0d#)) OR
 					(reg_q2577 AND symb_decoder(16#0a#)) OR
 					(reg_q2577 AND symb_decoder(16#09#)) OR
 					(reg_q2577 AND symb_decoder(16#20#));
reg_q2579_init <= '0' ;
	p_reg_q2579: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2579 <= reg_q2579_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2579 <= reg_q2579_init;
        else
          reg_q2579 <= reg_q2579_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q671_in <= (reg_q669 AND symb_decoder(16#46#)) OR
 					(reg_q669 AND symb_decoder(16#66#));
reg_q671_init <= '0' ;
	p_reg_q671: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q671 <= reg_q671_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q671 <= reg_q671_init;
        else
          reg_q671 <= reg_q671_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q673_in <= (reg_q671 AND symb_decoder(16#73#)) OR
 					(reg_q671 AND symb_decoder(16#48#)) OR
 					(reg_q671 AND symb_decoder(16#70#)) OR
 					(reg_q671 AND symb_decoder(16#72#)) OR
 					(reg_q671 AND symb_decoder(16#59#)) OR
 					(reg_q671 AND symb_decoder(16#4b#)) OR
 					(reg_q671 AND symb_decoder(16#64#)) OR
 					(reg_q671 AND symb_decoder(16#55#)) OR
 					(reg_q671 AND symb_decoder(16#76#)) OR
 					(reg_q671 AND symb_decoder(16#7a#)) OR
 					(reg_q671 AND symb_decoder(16#68#)) OR
 					(reg_q671 AND symb_decoder(16#41#)) OR
 					(reg_q671 AND symb_decoder(16#65#)) OR
 					(reg_q671 AND symb_decoder(16#66#)) OR
 					(reg_q671 AND symb_decoder(16#6f#)) OR
 					(reg_q671 AND symb_decoder(16#62#)) OR
 					(reg_q671 AND symb_decoder(16#4a#)) OR
 					(reg_q671 AND symb_decoder(16#74#)) OR
 					(reg_q671 AND symb_decoder(16#56#)) OR
 					(reg_q671 AND symb_decoder(16#42#)) OR
 					(reg_q671 AND symb_decoder(16#49#)) OR
 					(reg_q671 AND symb_decoder(16#52#)) OR
 					(reg_q671 AND symb_decoder(16#4d#)) OR
 					(reg_q671 AND symb_decoder(16#6e#)) OR
 					(reg_q671 AND symb_decoder(16#67#)) OR
 					(reg_q671 AND symb_decoder(16#6a#)) OR
 					(reg_q671 AND symb_decoder(16#43#)) OR
 					(reg_q671 AND symb_decoder(16#71#)) OR
 					(reg_q671 AND symb_decoder(16#50#)) OR
 					(reg_q671 AND symb_decoder(16#46#)) OR
 					(reg_q671 AND symb_decoder(16#51#)) OR
 					(reg_q671 AND symb_decoder(16#44#)) OR
 					(reg_q671 AND symb_decoder(16#78#)) OR
 					(reg_q671 AND symb_decoder(16#45#)) OR
 					(reg_q671 AND symb_decoder(16#63#)) OR
 					(reg_q671 AND symb_decoder(16#4f#)) OR
 					(reg_q671 AND symb_decoder(16#54#)) OR
 					(reg_q671 AND symb_decoder(16#75#)) OR
 					(reg_q671 AND symb_decoder(16#6d#)) OR
 					(reg_q671 AND symb_decoder(16#6b#)) OR
 					(reg_q671 AND symb_decoder(16#47#)) OR
 					(reg_q671 AND symb_decoder(16#6c#)) OR
 					(reg_q671 AND symb_decoder(16#77#)) OR
 					(reg_q671 AND symb_decoder(16#61#)) OR
 					(reg_q671 AND symb_decoder(16#58#)) OR
 					(reg_q671 AND symb_decoder(16#57#)) OR
 					(reg_q671 AND symb_decoder(16#5a#)) OR
 					(reg_q671 AND symb_decoder(16#4e#)) OR
 					(reg_q671 AND symb_decoder(16#4c#)) OR
 					(reg_q671 AND symb_decoder(16#69#)) OR
 					(reg_q671 AND symb_decoder(16#53#)) OR
 					(reg_q671 AND symb_decoder(16#79#));
reg_q673_init <= '0' ;
	p_reg_q673: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q673 <= reg_q673_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q673 <= reg_q673_init;
        else
          reg_q673 <= reg_q673_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2_in <= (reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q0 AND symb_decoder(16#30#));
reg_q2_init <= '0' ;
	p_reg_q2: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2 <= reg_q2_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2 <= reg_q2_init;
        else
          reg_q2 <= reg_q2_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2323_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2323 AND symb_decoder(16#18#)) OR
 					(reg_q2323 AND symb_decoder(16#f8#)) OR
 					(reg_q2323 AND symb_decoder(16#cc#)) OR
 					(reg_q2323 AND symb_decoder(16#85#)) OR
 					(reg_q2323 AND symb_decoder(16#fc#)) OR
 					(reg_q2323 AND symb_decoder(16#47#)) OR
 					(reg_q2323 AND symb_decoder(16#c9#)) OR
 					(reg_q2323 AND symb_decoder(16#14#)) OR
 					(reg_q2323 AND symb_decoder(16#99#)) OR
 					(reg_q2323 AND symb_decoder(16#32#)) OR
 					(reg_q2323 AND symb_decoder(16#61#)) OR
 					(reg_q2323 AND symb_decoder(16#e8#)) OR
 					(reg_q2323 AND symb_decoder(16#5c#)) OR
 					(reg_q2323 AND symb_decoder(16#46#)) OR
 					(reg_q2323 AND symb_decoder(16#fa#)) OR
 					(reg_q2323 AND symb_decoder(16#c1#)) OR
 					(reg_q2323 AND symb_decoder(16#a8#)) OR
 					(reg_q2323 AND symb_decoder(16#ee#)) OR
 					(reg_q2323 AND symb_decoder(16#c4#)) OR
 					(reg_q2323 AND symb_decoder(16#97#)) OR
 					(reg_q2323 AND symb_decoder(16#e4#)) OR
 					(reg_q2323 AND symb_decoder(16#16#)) OR
 					(reg_q2323 AND symb_decoder(16#02#)) OR
 					(reg_q2323 AND symb_decoder(16#8d#)) OR
 					(reg_q2323 AND symb_decoder(16#f9#)) OR
 					(reg_q2323 AND symb_decoder(16#83#)) OR
 					(reg_q2323 AND symb_decoder(16#40#)) OR
 					(reg_q2323 AND symb_decoder(16#ef#)) OR
 					(reg_q2323 AND symb_decoder(16#60#)) OR
 					(reg_q2323 AND symb_decoder(16#55#)) OR
 					(reg_q2323 AND symb_decoder(16#93#)) OR
 					(reg_q2323 AND symb_decoder(16#26#)) OR
 					(reg_q2323 AND symb_decoder(16#1c#)) OR
 					(reg_q2323 AND symb_decoder(16#3d#)) OR
 					(reg_q2323 AND symb_decoder(16#53#)) OR
 					(reg_q2323 AND symb_decoder(16#ea#)) OR
 					(reg_q2323 AND symb_decoder(16#a5#)) OR
 					(reg_q2323 AND symb_decoder(16#c2#)) OR
 					(reg_q2323 AND symb_decoder(16#0c#)) OR
 					(reg_q2323 AND symb_decoder(16#74#)) OR
 					(reg_q2323 AND symb_decoder(16#ab#)) OR
 					(reg_q2323 AND symb_decoder(16#62#)) OR
 					(reg_q2323 AND symb_decoder(16#d1#)) OR
 					(reg_q2323 AND symb_decoder(16#b0#)) OR
 					(reg_q2323 AND symb_decoder(16#10#)) OR
 					(reg_q2323 AND symb_decoder(16#a7#)) OR
 					(reg_q2323 AND symb_decoder(16#3a#)) OR
 					(reg_q2323 AND symb_decoder(16#4f#)) OR
 					(reg_q2323 AND symb_decoder(16#db#)) OR
 					(reg_q2323 AND symb_decoder(16#f3#)) OR
 					(reg_q2323 AND symb_decoder(16#05#)) OR
 					(reg_q2323 AND symb_decoder(16#12#)) OR
 					(reg_q2323 AND symb_decoder(16#0e#)) OR
 					(reg_q2323 AND symb_decoder(16#d9#)) OR
 					(reg_q2323 AND symb_decoder(16#66#)) OR
 					(reg_q2323 AND symb_decoder(16#e5#)) OR
 					(reg_q2323 AND symb_decoder(16#cd#)) OR
 					(reg_q2323 AND symb_decoder(16#c6#)) OR
 					(reg_q2323 AND symb_decoder(16#aa#)) OR
 					(reg_q2323 AND symb_decoder(16#b2#)) OR
 					(reg_q2323 AND symb_decoder(16#5d#)) OR
 					(reg_q2323 AND symb_decoder(16#3f#)) OR
 					(reg_q2323 AND symb_decoder(16#d0#)) OR
 					(reg_q2323 AND symb_decoder(16#a6#)) OR
 					(reg_q2323 AND symb_decoder(16#8a#)) OR
 					(reg_q2323 AND symb_decoder(16#07#)) OR
 					(reg_q2323 AND symb_decoder(16#1a#)) OR
 					(reg_q2323 AND symb_decoder(16#d7#)) OR
 					(reg_q2323 AND symb_decoder(16#eb#)) OR
 					(reg_q2323 AND symb_decoder(16#fd#)) OR
 					(reg_q2323 AND symb_decoder(16#0a#)) OR
 					(reg_q2323 AND symb_decoder(16#82#)) OR
 					(reg_q2323 AND symb_decoder(16#d8#)) OR
 					(reg_q2323 AND symb_decoder(16#11#)) OR
 					(reg_q2323 AND symb_decoder(16#cf#)) OR
 					(reg_q2323 AND symb_decoder(16#77#)) OR
 					(reg_q2323 AND symb_decoder(16#b9#)) OR
 					(reg_q2323 AND symb_decoder(16#23#)) OR
 					(reg_q2323 AND symb_decoder(16#79#)) OR
 					(reg_q2323 AND symb_decoder(16#03#)) OR
 					(reg_q2323 AND symb_decoder(16#4c#)) OR
 					(reg_q2323 AND symb_decoder(16#1b#)) OR
 					(reg_q2323 AND symb_decoder(16#b7#)) OR
 					(reg_q2323 AND symb_decoder(16#be#)) OR
 					(reg_q2323 AND symb_decoder(16#f7#)) OR
 					(reg_q2323 AND symb_decoder(16#ca#)) OR
 					(reg_q2323 AND symb_decoder(16#88#)) OR
 					(reg_q2323 AND symb_decoder(16#f0#)) OR
 					(reg_q2323 AND symb_decoder(16#2c#)) OR
 					(reg_q2323 AND symb_decoder(16#c0#)) OR
 					(reg_q2323 AND symb_decoder(16#5b#)) OR
 					(reg_q2323 AND symb_decoder(16#98#)) OR
 					(reg_q2323 AND symb_decoder(16#90#)) OR
 					(reg_q2323 AND symb_decoder(16#b4#)) OR
 					(reg_q2323 AND symb_decoder(16#c3#)) OR
 					(reg_q2323 AND symb_decoder(16#57#)) OR
 					(reg_q2323 AND symb_decoder(16#67#)) OR
 					(reg_q2323 AND symb_decoder(16#15#)) OR
 					(reg_q2323 AND symb_decoder(16#e7#)) OR
 					(reg_q2323 AND symb_decoder(16#a9#)) OR
 					(reg_q2323 AND symb_decoder(16#ae#)) OR
 					(reg_q2323 AND symb_decoder(16#09#)) OR
 					(reg_q2323 AND symb_decoder(16#c8#)) OR
 					(reg_q2323 AND symb_decoder(16#28#)) OR
 					(reg_q2323 AND symb_decoder(16#0d#)) OR
 					(reg_q2323 AND symb_decoder(16#d3#)) OR
 					(reg_q2323 AND symb_decoder(16#71#)) OR
 					(reg_q2323 AND symb_decoder(16#24#)) OR
 					(reg_q2323 AND symb_decoder(16#b5#)) OR
 					(reg_q2323 AND symb_decoder(16#f6#)) OR
 					(reg_q2323 AND symb_decoder(16#08#)) OR
 					(reg_q2323 AND symb_decoder(16#58#)) OR
 					(reg_q2323 AND symb_decoder(16#9e#)) OR
 					(reg_q2323 AND symb_decoder(16#35#)) OR
 					(reg_q2323 AND symb_decoder(16#d5#)) OR
 					(reg_q2323 AND symb_decoder(16#e2#)) OR
 					(reg_q2323 AND symb_decoder(16#8b#)) OR
 					(reg_q2323 AND symb_decoder(16#44#)) OR
 					(reg_q2323 AND symb_decoder(16#48#)) OR
 					(reg_q2323 AND symb_decoder(16#73#)) OR
 					(reg_q2323 AND symb_decoder(16#76#)) OR
 					(reg_q2323 AND symb_decoder(16#5a#)) OR
 					(reg_q2323 AND symb_decoder(16#00#)) OR
 					(reg_q2323 AND symb_decoder(16#94#)) OR
 					(reg_q2323 AND symb_decoder(16#8e#)) OR
 					(reg_q2323 AND symb_decoder(16#bf#)) OR
 					(reg_q2323 AND symb_decoder(16#a2#)) OR
 					(reg_q2323 AND symb_decoder(16#4a#)) OR
 					(reg_q2323 AND symb_decoder(16#20#)) OR
 					(reg_q2323 AND symb_decoder(16#0f#)) OR
 					(reg_q2323 AND symb_decoder(16#19#)) OR
 					(reg_q2323 AND symb_decoder(16#2f#)) OR
 					(reg_q2323 AND symb_decoder(16#b8#)) OR
 					(reg_q2323 AND symb_decoder(16#68#)) OR
 					(reg_q2323 AND symb_decoder(16#fe#)) OR
 					(reg_q2323 AND symb_decoder(16#45#)) OR
 					(reg_q2323 AND symb_decoder(16#49#)) OR
 					(reg_q2323 AND symb_decoder(16#13#)) OR
 					(reg_q2323 AND symb_decoder(16#a3#)) OR
 					(reg_q2323 AND symb_decoder(16#ec#)) OR
 					(reg_q2323 AND symb_decoder(16#84#)) OR
 					(reg_q2323 AND symb_decoder(16#d4#)) OR
 					(reg_q2323 AND symb_decoder(16#8f#)) OR
 					(reg_q2323 AND symb_decoder(16#27#)) OR
 					(reg_q2323 AND symb_decoder(16#da#)) OR
 					(reg_q2323 AND symb_decoder(16#9a#)) OR
 					(reg_q2323 AND symb_decoder(16#c5#)) OR
 					(reg_q2323 AND symb_decoder(16#87#)) OR
 					(reg_q2323 AND symb_decoder(16#70#)) OR
 					(reg_q2323 AND symb_decoder(16#b3#)) OR
 					(reg_q2323 AND symb_decoder(16#65#)) OR
 					(reg_q2323 AND symb_decoder(16#3e#)) OR
 					(reg_q2323 AND symb_decoder(16#6c#)) OR
 					(reg_q2323 AND symb_decoder(16#e0#)) OR
 					(reg_q2323 AND symb_decoder(16#3c#)) OR
 					(reg_q2323 AND symb_decoder(16#fb#)) OR
 					(reg_q2323 AND symb_decoder(16#7b#)) OR
 					(reg_q2323 AND symb_decoder(16#7f#)) OR
 					(reg_q2323 AND symb_decoder(16#01#)) OR
 					(reg_q2323 AND symb_decoder(16#8c#)) OR
 					(reg_q2323 AND symb_decoder(16#7d#)) OR
 					(reg_q2323 AND symb_decoder(16#f4#)) OR
 					(reg_q2323 AND symb_decoder(16#ff#)) OR
 					(reg_q2323 AND symb_decoder(16#6b#)) OR
 					(reg_q2323 AND symb_decoder(16#2a#)) OR
 					(reg_q2323 AND symb_decoder(16#81#)) OR
 					(reg_q2323 AND symb_decoder(16#dc#)) OR
 					(reg_q2323 AND symb_decoder(16#34#)) OR
 					(reg_q2323 AND symb_decoder(16#de#)) OR
 					(reg_q2323 AND symb_decoder(16#f5#)) OR
 					(reg_q2323 AND symb_decoder(16#a1#)) OR
 					(reg_q2323 AND symb_decoder(16#80#)) OR
 					(reg_q2323 AND symb_decoder(16#50#)) OR
 					(reg_q2323 AND symb_decoder(16#29#)) OR
 					(reg_q2323 AND symb_decoder(16#9c#)) OR
 					(reg_q2323 AND symb_decoder(16#22#)) OR
 					(reg_q2323 AND symb_decoder(16#e6#)) OR
 					(reg_q2323 AND symb_decoder(16#06#)) OR
 					(reg_q2323 AND symb_decoder(16#bb#)) OR
 					(reg_q2323 AND symb_decoder(16#63#)) OR
 					(reg_q2323 AND symb_decoder(16#f2#)) OR
 					(reg_q2323 AND symb_decoder(16#3b#)) OR
 					(reg_q2323 AND symb_decoder(16#e3#)) OR
 					(reg_q2323 AND symb_decoder(16#cb#)) OR
 					(reg_q2323 AND symb_decoder(16#64#)) OR
 					(reg_q2323 AND symb_decoder(16#37#)) OR
 					(reg_q2323 AND symb_decoder(16#91#)) OR
 					(reg_q2323 AND symb_decoder(16#38#)) OR
 					(reg_q2323 AND symb_decoder(16#7e#)) OR
 					(reg_q2323 AND symb_decoder(16#51#)) OR
 					(reg_q2323 AND symb_decoder(16#78#)) OR
 					(reg_q2323 AND symb_decoder(16#ac#)) OR
 					(reg_q2323 AND symb_decoder(16#41#)) OR
 					(reg_q2323 AND symb_decoder(16#21#)) OR
 					(reg_q2323 AND symb_decoder(16#df#)) OR
 					(reg_q2323 AND symb_decoder(16#4d#)) OR
 					(reg_q2323 AND symb_decoder(16#56#)) OR
 					(reg_q2323 AND symb_decoder(16#86#)) OR
 					(reg_q2323 AND symb_decoder(16#89#)) OR
 					(reg_q2323 AND symb_decoder(16#92#)) OR
 					(reg_q2323 AND symb_decoder(16#6f#)) OR
 					(reg_q2323 AND symb_decoder(16#4b#)) OR
 					(reg_q2323 AND symb_decoder(16#96#)) OR
 					(reg_q2323 AND symb_decoder(16#43#)) OR
 					(reg_q2323 AND symb_decoder(16#75#)) OR
 					(reg_q2323 AND symb_decoder(16#2e#)) OR
 					(reg_q2323 AND symb_decoder(16#52#)) OR
 					(reg_q2323 AND symb_decoder(16#59#)) OR
 					(reg_q2323 AND symb_decoder(16#ad#)) OR
 					(reg_q2323 AND symb_decoder(16#39#)) OR
 					(reg_q2323 AND symb_decoder(16#72#)) OR
 					(reg_q2323 AND symb_decoder(16#e9#)) OR
 					(reg_q2323 AND symb_decoder(16#04#)) OR
 					(reg_q2323 AND symb_decoder(16#ed#)) OR
 					(reg_q2323 AND symb_decoder(16#dd#)) OR
 					(reg_q2323 AND symb_decoder(16#17#)) OR
 					(reg_q2323 AND symb_decoder(16#b6#)) OR
 					(reg_q2323 AND symb_decoder(16#5e#)) OR
 					(reg_q2323 AND symb_decoder(16#5f#)) OR
 					(reg_q2323 AND symb_decoder(16#69#)) OR
 					(reg_q2323 AND symb_decoder(16#bc#)) OR
 					(reg_q2323 AND symb_decoder(16#ce#)) OR
 					(reg_q2323 AND symb_decoder(16#31#)) OR
 					(reg_q2323 AND symb_decoder(16#c7#)) OR
 					(reg_q2323 AND symb_decoder(16#1d#)) OR
 					(reg_q2323 AND symb_decoder(16#9b#)) OR
 					(reg_q2323 AND symb_decoder(16#54#)) OR
 					(reg_q2323 AND symb_decoder(16#a0#)) OR
 					(reg_q2323 AND symb_decoder(16#33#)) OR
 					(reg_q2323 AND symb_decoder(16#6e#)) OR
 					(reg_q2323 AND symb_decoder(16#2d#)) OR
 					(reg_q2323 AND symb_decoder(16#6d#)) OR
 					(reg_q2323 AND symb_decoder(16#30#)) OR
 					(reg_q2323 AND symb_decoder(16#d2#)) OR
 					(reg_q2323 AND symb_decoder(16#0b#)) OR
 					(reg_q2323 AND symb_decoder(16#6a#)) OR
 					(reg_q2323 AND symb_decoder(16#af#)) OR
 					(reg_q2323 AND symb_decoder(16#d6#)) OR
 					(reg_q2323 AND symb_decoder(16#a4#)) OR
 					(reg_q2323 AND symb_decoder(16#7a#)) OR
 					(reg_q2323 AND symb_decoder(16#9f#)) OR
 					(reg_q2323 AND symb_decoder(16#1f#)) OR
 					(reg_q2323 AND symb_decoder(16#4e#)) OR
 					(reg_q2323 AND symb_decoder(16#9d#)) OR
 					(reg_q2323 AND symb_decoder(16#e1#)) OR
 					(reg_q2323 AND symb_decoder(16#2b#)) OR
 					(reg_q2323 AND symb_decoder(16#b1#)) OR
 					(reg_q2323 AND symb_decoder(16#f1#)) OR
 					(reg_q2323 AND symb_decoder(16#ba#)) OR
 					(reg_q2323 AND symb_decoder(16#25#)) OR
 					(reg_q2323 AND symb_decoder(16#7c#)) OR
 					(reg_q2323 AND symb_decoder(16#42#)) OR
 					(reg_q2323 AND symb_decoder(16#36#)) OR
 					(reg_q2323 AND symb_decoder(16#bd#)) OR
 					(reg_q2323 AND symb_decoder(16#1e#)) OR
 					(reg_q2323 AND symb_decoder(16#95#));
reg_q2323_init <= '0' ;
	p_reg_q2323: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2323 <= reg_q2323_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2323 <= reg_q2323_init;
        else
          reg_q2323 <= reg_q2323_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2128_in <= (reg_q2126 AND symb_decoder(16#65#)) OR
 					(reg_q2126 AND symb_decoder(16#45#));
reg_q2128_init <= '0' ;
	p_reg_q2128: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2128 <= reg_q2128_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2128 <= reg_q2128_init;
        else
          reg_q2128 <= reg_q2128_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2254_in <= (reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2253 AND symb_decoder(16#21#));
reg_q2254_init <= '0' ;
	p_reg_q2254: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2254 <= reg_q2254_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2254 <= reg_q2254_init;
        else
          reg_q2254 <= reg_q2254_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2256_in <= (reg_q2254 AND symb_decoder(16#21#));
reg_q2256_init <= '0' ;
	p_reg_q2256: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2256 <= reg_q2256_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2256 <= reg_q2256_init;
        else
          reg_q2256 <= reg_q2256_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q351_in <= (reg_q349 AND symb_decoder(16#53#)) OR
 					(reg_q349 AND symb_decoder(16#73#));
reg_q351_init <= '0' ;
	p_reg_q351: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q351 <= reg_q351_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q351 <= reg_q351_init;
        else
          reg_q351 <= reg_q351_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q353_in <= (reg_q351 AND symb_decoder(16#45#)) OR
 					(reg_q351 AND symb_decoder(16#65#));
reg_q353_init <= '0' ;
	p_reg_q353: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q353 <= reg_q353_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q353 <= reg_q353_init;
        else
          reg_q353 <= reg_q353_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2601_in <= (reg_q2601 AND symb_decoder(16#20#)) OR
 					(reg_q2601 AND symb_decoder(16#09#)) OR
 					(reg_q2601 AND symb_decoder(16#0d#)) OR
 					(reg_q2601 AND symb_decoder(16#0a#)) OR
 					(reg_q2601 AND symb_decoder(16#0c#)) OR
 					(reg_q2599 AND symb_decoder(16#0a#)) OR
 					(reg_q2599 AND symb_decoder(16#0d#)) OR
 					(reg_q2599 AND symb_decoder(16#20#)) OR
 					(reg_q2599 AND symb_decoder(16#0c#)) OR
 					(reg_q2599 AND symb_decoder(16#09#));
reg_q2601_init <= '0' ;
	p_reg_q2601: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2601 <= reg_q2601_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2601 <= reg_q2601_init;
        else
          reg_q2601 <= reg_q2601_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1393_in <= (reg_q1391 AND symb_decoder(16#3a#));
reg_q1393_init <= '0' ;
	p_reg_q1393: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1393 <= reg_q1393_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1393 <= reg_q1393_init;
        else
          reg_q1393 <= reg_q1393_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1395_in <= (reg_q1393 AND symb_decoder(16#0a#)) OR
 					(reg_q1393 AND symb_decoder(16#0c#)) OR
 					(reg_q1393 AND symb_decoder(16#20#)) OR
 					(reg_q1393 AND symb_decoder(16#0d#)) OR
 					(reg_q1393 AND symb_decoder(16#09#)) OR
 					(reg_q1395 AND symb_decoder(16#0d#)) OR
 					(reg_q1395 AND symb_decoder(16#0a#)) OR
 					(reg_q1395 AND symb_decoder(16#0c#)) OR
 					(reg_q1395 AND symb_decoder(16#20#)) OR
 					(reg_q1395 AND symb_decoder(16#09#));
reg_q1395_init <= '0' ;
	p_reg_q1395: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1395 <= reg_q1395_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1395 <= reg_q1395_init;
        else
          reg_q1395 <= reg_q1395_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q876_in <= (reg_q874 AND symb_decoder(16#5d#));
reg_q876_init <= '0' ;
	p_reg_q876: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q876 <= reg_q876_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q876 <= reg_q876_init;
        else
          reg_q876 <= reg_q876_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q878_in <= (reg_q876 AND symb_decoder(16#36#)) OR
 					(reg_q876 AND symb_decoder(16#30#)) OR
 					(reg_q876 AND symb_decoder(16#31#)) OR
 					(reg_q876 AND symb_decoder(16#35#)) OR
 					(reg_q876 AND symb_decoder(16#33#)) OR
 					(reg_q876 AND symb_decoder(16#34#)) OR
 					(reg_q876 AND symb_decoder(16#38#)) OR
 					(reg_q876 AND symb_decoder(16#37#)) OR
 					(reg_q876 AND symb_decoder(16#32#)) OR
 					(reg_q876 AND symb_decoder(16#39#));
reg_q878_init <= '0' ;
	p_reg_q878: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q878 <= reg_q878_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q878 <= reg_q878_init;
        else
          reg_q878 <= reg_q878_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1535_in <= (reg_q1535 AND symb_decoder(16#20#)) OR
 					(reg_q1535 AND symb_decoder(16#09#)) OR
 					(reg_q1535 AND symb_decoder(16#0c#)) OR
 					(reg_q1535 AND symb_decoder(16#0a#)) OR
 					(reg_q1535 AND symb_decoder(16#0d#)) OR
 					(reg_q1533 AND symb_decoder(16#20#)) OR
 					(reg_q1533 AND symb_decoder(16#0d#)) OR
 					(reg_q1533 AND symb_decoder(16#0a#)) OR
 					(reg_q1533 AND symb_decoder(16#09#)) OR
 					(reg_q1533 AND symb_decoder(16#0c#));
reg_q1535_init <= '0' ;
	p_reg_q1535: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1535 <= reg_q1535_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1535 <= reg_q1535_init;
        else
          reg_q1535 <= reg_q1535_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1537_in <= (reg_q1535 AND symb_decoder(16#37#)) OR
 					(reg_q1535 AND symb_decoder(16#39#)) OR
 					(reg_q1535 AND symb_decoder(16#36#)) OR
 					(reg_q1535 AND symb_decoder(16#35#)) OR
 					(reg_q1535 AND symb_decoder(16#33#)) OR
 					(reg_q1535 AND symb_decoder(16#32#)) OR
 					(reg_q1535 AND symb_decoder(16#30#)) OR
 					(reg_q1535 AND symb_decoder(16#34#)) OR
 					(reg_q1535 AND symb_decoder(16#31#)) OR
 					(reg_q1535 AND symb_decoder(16#38#)) OR
 					(reg_q1537 AND symb_decoder(16#37#)) OR
 					(reg_q1537 AND symb_decoder(16#38#)) OR
 					(reg_q1537 AND symb_decoder(16#30#)) OR
 					(reg_q1537 AND symb_decoder(16#35#)) OR
 					(reg_q1537 AND symb_decoder(16#32#)) OR
 					(reg_q1537 AND symb_decoder(16#36#)) OR
 					(reg_q1537 AND symb_decoder(16#33#)) OR
 					(reg_q1537 AND symb_decoder(16#39#)) OR
 					(reg_q1537 AND symb_decoder(16#34#)) OR
 					(reg_q1537 AND symb_decoder(16#31#));
reg_q1537_init <= '0' ;
	p_reg_q1537: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1537 <= reg_q1537_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1537 <= reg_q1537_init;
        else
          reg_q1537 <= reg_q1537_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q844_in <= (reg_q844 AND symb_decoder(16#33#)) OR
 					(reg_q844 AND symb_decoder(16#32#)) OR
 					(reg_q844 AND symb_decoder(16#36#)) OR
 					(reg_q844 AND symb_decoder(16#38#)) OR
 					(reg_q844 AND symb_decoder(16#39#)) OR
 					(reg_q844 AND symb_decoder(16#31#)) OR
 					(reg_q844 AND symb_decoder(16#30#)) OR
 					(reg_q844 AND symb_decoder(16#34#)) OR
 					(reg_q844 AND symb_decoder(16#35#)) OR
 					(reg_q844 AND symb_decoder(16#37#)) OR
 					(reg_q842 AND symb_decoder(16#32#)) OR
 					(reg_q842 AND symb_decoder(16#37#)) OR
 					(reg_q842 AND symb_decoder(16#30#)) OR
 					(reg_q842 AND symb_decoder(16#31#)) OR
 					(reg_q842 AND symb_decoder(16#34#)) OR
 					(reg_q842 AND symb_decoder(16#33#)) OR
 					(reg_q842 AND symb_decoder(16#38#)) OR
 					(reg_q842 AND symb_decoder(16#39#)) OR
 					(reg_q842 AND symb_decoder(16#36#)) OR
 					(reg_q842 AND symb_decoder(16#35#));
reg_q844_init <= '0' ;
	p_reg_q844: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q844 <= reg_q844_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q844 <= reg_q844_init;
        else
          reg_q844 <= reg_q844_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q257_in <= (reg_q257 AND symb_decoder(16#34#)) OR
 					(reg_q257 AND symb_decoder(16#30#)) OR
 					(reg_q257 AND symb_decoder(16#32#)) OR
 					(reg_q257 AND symb_decoder(16#35#)) OR
 					(reg_q257 AND symb_decoder(16#37#)) OR
 					(reg_q257 AND symb_decoder(16#36#)) OR
 					(reg_q257 AND symb_decoder(16#31#)) OR
 					(reg_q257 AND symb_decoder(16#39#)) OR
 					(reg_q257 AND symb_decoder(16#38#)) OR
 					(reg_q257 AND symb_decoder(16#33#)) OR
 					(reg_q255 AND symb_decoder(16#37#)) OR
 					(reg_q255 AND symb_decoder(16#34#)) OR
 					(reg_q255 AND symb_decoder(16#39#)) OR
 					(reg_q255 AND symb_decoder(16#32#)) OR
 					(reg_q255 AND symb_decoder(16#35#)) OR
 					(reg_q255 AND symb_decoder(16#36#)) OR
 					(reg_q255 AND symb_decoder(16#31#)) OR
 					(reg_q255 AND symb_decoder(16#38#)) OR
 					(reg_q255 AND symb_decoder(16#30#)) OR
 					(reg_q255 AND symb_decoder(16#33#));
reg_q257_init <= '0' ;
	p_reg_q257: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q257 <= reg_q257_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q257 <= reg_q257_init;
        else
          reg_q257 <= reg_q257_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1313_in <= (reg_q1311 AND symb_decoder(16#65#)) OR
 					(reg_q1311 AND symb_decoder(16#45#));
reg_q1313_init <= '0' ;
	p_reg_q1313: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1313 <= reg_q1313_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1313 <= reg_q1313_init;
        else
          reg_q1313 <= reg_q1313_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1315_in <= (reg_q1313 AND symb_decoder(16#6e#)) OR
 					(reg_q1313 AND symb_decoder(16#4e#));
reg_q1315_init <= '0' ;
	p_reg_q1315: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1315 <= reg_q1315_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1315 <= reg_q1315_init;
        else
          reg_q1315 <= reg_q1315_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q880_in <= (reg_q878 AND symb_decoder(16#00#)) OR
 					(reg_q887 AND symb_decoder(16#00#)) OR
 					(reg_q884 AND symb_decoder(16#00#)) OR
 					(reg_q886 AND symb_decoder(16#00#));
reg_q880_init <= '0' ;
	p_reg_q880: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q880 <= reg_q880_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q880 <= reg_q880_init;
        else
          reg_q880 <= reg_q880_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q882_in <= (reg_q880 AND symb_decoder(16#62#)) OR
 					(reg_q880 AND symb_decoder(16#63#)) OR
 					(reg_q880 AND symb_decoder(16#68#)) OR
 					(reg_q880 AND symb_decoder(16#44#)) OR
 					(reg_q880 AND symb_decoder(16#64#)) OR
 					(reg_q880 AND symb_decoder(16#75#)) OR
 					(reg_q880 AND symb_decoder(16#65#)) OR
 					(reg_q880 AND symb_decoder(16#4d#)) OR
 					(reg_q880 AND symb_decoder(16#57#)) OR
 					(reg_q880 AND symb_decoder(16#7a#)) OR
 					(reg_q880 AND symb_decoder(16#6b#)) OR
 					(reg_q880 AND symb_decoder(16#56#)) OR
 					(reg_q880 AND symb_decoder(16#6a#)) OR
 					(reg_q880 AND symb_decoder(16#47#)) OR
 					(reg_q880 AND symb_decoder(16#41#)) OR
 					(reg_q880 AND symb_decoder(16#79#)) OR
 					(reg_q880 AND symb_decoder(16#45#)) OR
 					(reg_q880 AND symb_decoder(16#4b#)) OR
 					(reg_q880 AND symb_decoder(16#51#)) OR
 					(reg_q880 AND symb_decoder(16#50#)) OR
 					(reg_q880 AND symb_decoder(16#70#)) OR
 					(reg_q880 AND symb_decoder(16#55#)) OR
 					(reg_q880 AND symb_decoder(16#76#)) OR
 					(reg_q880 AND symb_decoder(16#52#)) OR
 					(reg_q880 AND symb_decoder(16#67#)) OR
 					(reg_q880 AND symb_decoder(16#4f#)) OR
 					(reg_q880 AND symb_decoder(16#6e#)) OR
 					(reg_q880 AND symb_decoder(16#73#)) OR
 					(reg_q880 AND symb_decoder(16#43#)) OR
 					(reg_q880 AND symb_decoder(16#59#)) OR
 					(reg_q880 AND symb_decoder(16#53#)) OR
 					(reg_q880 AND symb_decoder(16#54#)) OR
 					(reg_q880 AND symb_decoder(16#46#)) OR
 					(reg_q880 AND symb_decoder(16#5a#)) OR
 					(reg_q880 AND symb_decoder(16#42#)) OR
 					(reg_q880 AND symb_decoder(16#66#)) OR
 					(reg_q880 AND symb_decoder(16#6d#)) OR
 					(reg_q880 AND symb_decoder(16#72#)) OR
 					(reg_q880 AND symb_decoder(16#49#)) OR
 					(reg_q880 AND symb_decoder(16#6c#)) OR
 					(reg_q880 AND symb_decoder(16#4a#)) OR
 					(reg_q880 AND symb_decoder(16#61#)) OR
 					(reg_q880 AND symb_decoder(16#4e#)) OR
 					(reg_q880 AND symb_decoder(16#77#)) OR
 					(reg_q880 AND symb_decoder(16#6f#)) OR
 					(reg_q880 AND symb_decoder(16#4c#)) OR
 					(reg_q880 AND symb_decoder(16#78#)) OR
 					(reg_q880 AND symb_decoder(16#58#)) OR
 					(reg_q880 AND symb_decoder(16#71#)) OR
 					(reg_q880 AND symb_decoder(16#74#)) OR
 					(reg_q880 AND symb_decoder(16#48#)) OR
 					(reg_q880 AND symb_decoder(16#69#));
reg_q882_init <= '0' ;
	p_reg_q882: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q882 <= reg_q882_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q882 <= reg_q882_init;
        else
          reg_q882 <= reg_q882_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q807_in <= (reg_q805 AND symb_decoder(16#2e#));
reg_q807_init <= '0' ;
	p_reg_q807: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q807 <= reg_q807_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q807 <= reg_q807_init;
        else
          reg_q807 <= reg_q807_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q809_in <= (reg_q807 AND symb_decoder(16#34#)) OR
 					(reg_q807 AND symb_decoder(16#33#)) OR
 					(reg_q807 AND symb_decoder(16#39#)) OR
 					(reg_q807 AND symb_decoder(16#32#)) OR
 					(reg_q807 AND symb_decoder(16#38#)) OR
 					(reg_q807 AND symb_decoder(16#35#)) OR
 					(reg_q807 AND symb_decoder(16#37#)) OR
 					(reg_q807 AND symb_decoder(16#30#)) OR
 					(reg_q807 AND symb_decoder(16#31#)) OR
 					(reg_q807 AND symb_decoder(16#36#)) OR
 					(reg_q809 AND symb_decoder(16#35#)) OR
 					(reg_q809 AND symb_decoder(16#37#)) OR
 					(reg_q809 AND symb_decoder(16#33#)) OR
 					(reg_q809 AND symb_decoder(16#38#)) OR
 					(reg_q809 AND symb_decoder(16#34#)) OR
 					(reg_q809 AND symb_decoder(16#36#)) OR
 					(reg_q809 AND symb_decoder(16#31#)) OR
 					(reg_q809 AND symb_decoder(16#30#)) OR
 					(reg_q809 AND symb_decoder(16#39#)) OR
 					(reg_q809 AND symb_decoder(16#32#));
reg_q809_init <= '0' ;
	p_reg_q809: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q809 <= reg_q809_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q809 <= reg_q809_init;
        else
          reg_q809 <= reg_q809_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q379_in <= (reg_q377 AND symb_decoder(16#45#)) OR
 					(reg_q377 AND symb_decoder(16#65#));
reg_q379_init <= '0' ;
	p_reg_q379: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q379 <= reg_q379_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q379 <= reg_q379_init;
        else
          reg_q379 <= reg_q379_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q381_in <= (reg_q379 AND symb_decoder(16#0d#)) OR
 					(reg_q379 AND symb_decoder(16#0a#)) OR
 					(reg_q379 AND symb_decoder(16#09#)) OR
 					(reg_q379 AND symb_decoder(16#0c#)) OR
 					(reg_q379 AND symb_decoder(16#20#)) OR
 					(reg_q381 AND symb_decoder(16#0a#)) OR
 					(reg_q381 AND symb_decoder(16#09#)) OR
 					(reg_q381 AND symb_decoder(16#20#)) OR
 					(reg_q381 AND symb_decoder(16#0d#)) OR
 					(reg_q381 AND symb_decoder(16#0c#));
reg_q381_init <= '0' ;
	p_reg_q381: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q381 <= reg_q381_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q381 <= reg_q381_init;
        else
          reg_q381 <= reg_q381_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q832_in <= (reg_q828 AND symb_decoder(16#30#)) OR
 					(reg_q828 AND symb_decoder(16#34#)) OR
 					(reg_q828 AND symb_decoder(16#35#)) OR
 					(reg_q828 AND symb_decoder(16#39#)) OR
 					(reg_q828 AND symb_decoder(16#33#)) OR
 					(reg_q828 AND symb_decoder(16#37#)) OR
 					(reg_q828 AND symb_decoder(16#31#)) OR
 					(reg_q828 AND symb_decoder(16#36#)) OR
 					(reg_q828 AND symb_decoder(16#38#)) OR
 					(reg_q828 AND symb_decoder(16#32#)) OR
 					(reg_q848 AND symb_decoder(16#38#)) OR
 					(reg_q848 AND symb_decoder(16#35#)) OR
 					(reg_q848 AND symb_decoder(16#32#)) OR
 					(reg_q848 AND symb_decoder(16#30#)) OR
 					(reg_q848 AND symb_decoder(16#34#)) OR
 					(reg_q848 AND symb_decoder(16#33#)) OR
 					(reg_q848 AND symb_decoder(16#31#)) OR
 					(reg_q848 AND symb_decoder(16#36#)) OR
 					(reg_q848 AND symb_decoder(16#39#)) OR
 					(reg_q848 AND symb_decoder(16#37#)) OR
 					(reg_q832 AND symb_decoder(16#33#)) OR
 					(reg_q832 AND symb_decoder(16#36#)) OR
 					(reg_q832 AND symb_decoder(16#32#)) OR
 					(reg_q832 AND symb_decoder(16#31#)) OR
 					(reg_q832 AND symb_decoder(16#34#)) OR
 					(reg_q832 AND symb_decoder(16#30#)) OR
 					(reg_q832 AND symb_decoder(16#39#)) OR
 					(reg_q832 AND symb_decoder(16#38#)) OR
 					(reg_q832 AND symb_decoder(16#37#)) OR
 					(reg_q832 AND symb_decoder(16#35#));
reg_q832_init <= '0' ;
	p_reg_q832: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q832 <= reg_q832_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q832 <= reg_q832_init;
        else
          reg_q832 <= reg_q832_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q945_in <= (reg_q943 AND symb_decoder(16#2e#));
reg_q945_init <= '0' ;
	p_reg_q945: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q945 <= reg_q945_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q945 <= reg_q945_init;
        else
          reg_q945 <= reg_q945_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q947_in <= (reg_q945 AND symb_decoder(16#31#)) OR
 					(reg_q945 AND symb_decoder(16#34#)) OR
 					(reg_q945 AND symb_decoder(16#32#)) OR
 					(reg_q945 AND symb_decoder(16#30#)) OR
 					(reg_q945 AND symb_decoder(16#35#)) OR
 					(reg_q945 AND symb_decoder(16#33#)) OR
 					(reg_q945 AND symb_decoder(16#39#)) OR
 					(reg_q945 AND symb_decoder(16#36#)) OR
 					(reg_q945 AND symb_decoder(16#37#)) OR
 					(reg_q945 AND symb_decoder(16#38#)) OR
 					(reg_q947 AND symb_decoder(16#38#)) OR
 					(reg_q947 AND symb_decoder(16#32#)) OR
 					(reg_q947 AND symb_decoder(16#34#)) OR
 					(reg_q947 AND symb_decoder(16#35#)) OR
 					(reg_q947 AND symb_decoder(16#30#)) OR
 					(reg_q947 AND symb_decoder(16#31#)) OR
 					(reg_q947 AND symb_decoder(16#36#)) OR
 					(reg_q947 AND symb_decoder(16#39#)) OR
 					(reg_q947 AND symb_decoder(16#37#)) OR
 					(reg_q947 AND symb_decoder(16#33#));
reg_q947_init <= '0' ;
	p_reg_q947: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q947 <= reg_q947_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q947 <= reg_q947_init;
        else
          reg_q947 <= reg_q947_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2395_in <= (reg_q2393 AND symb_decoder(16#4f#)) OR
 					(reg_q2393 AND symb_decoder(16#6f#));
reg_q2395_init <= '0' ;
	p_reg_q2395: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2395 <= reg_q2395_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2395 <= reg_q2395_init;
        else
          reg_q2395 <= reg_q2395_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2397_in <= (reg_q2395 AND symb_decoder(16#4d#)) OR
 					(reg_q2395 AND symb_decoder(16#6d#));
reg_q2397_init <= '0' ;
	p_reg_q2397: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2397 <= reg_q2397_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2397 <= reg_q2397_init;
        else
          reg_q2397 <= reg_q2397_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1345_in <= (reg_q1345 AND symb_decoder(16#0c#)) OR
 					(reg_q1345 AND symb_decoder(16#09#)) OR
 					(reg_q1345 AND symb_decoder(16#0d#)) OR
 					(reg_q1345 AND symb_decoder(16#0a#)) OR
 					(reg_q1345 AND symb_decoder(16#20#)) OR
 					(reg_q1343 AND symb_decoder(16#0d#)) OR
 					(reg_q1343 AND symb_decoder(16#20#)) OR
 					(reg_q1343 AND symb_decoder(16#0c#)) OR
 					(reg_q1343 AND symb_decoder(16#0a#)) OR
 					(reg_q1343 AND symb_decoder(16#09#));
reg_q1345_init <= '0' ;
	p_reg_q1345: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1345 <= reg_q1345_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1345 <= reg_q1345_init;
        else
          reg_q1345 <= reg_q1345_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q566_in <= (reg_q564 AND symb_decoder(16#3d#));
reg_q566_init <= '0' ;
	p_reg_q566: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q566 <= reg_q566_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q566 <= reg_q566_init;
        else
          reg_q566 <= reg_q566_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q568_in <= (reg_q566 AND symb_decoder(16#25#));
reg_q568_init <= '0' ;
	p_reg_q568: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q568 <= reg_q568_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q568 <= reg_q568_init;
        else
          reg_q568 <= reg_q568_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2514_in <= (reg_q2512 AND symb_decoder(16#2a#));
reg_q2514_init <= '0' ;
	p_reg_q2514: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2514 <= reg_q2514_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2514 <= reg_q2514_init;
        else
          reg_q2514 <= reg_q2514_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2516_in <= (reg_q2514 AND symb_decoder(16#33#)) OR
 					(reg_q2514 AND symb_decoder(16#38#)) OR
 					(reg_q2514 AND symb_decoder(16#32#)) OR
 					(reg_q2514 AND symb_decoder(16#36#)) OR
 					(reg_q2514 AND symb_decoder(16#30#)) OR
 					(reg_q2514 AND symb_decoder(16#39#)) OR
 					(reg_q2514 AND symb_decoder(16#34#)) OR
 					(reg_q2514 AND symb_decoder(16#37#)) OR
 					(reg_q2514 AND symb_decoder(16#31#)) OR
 					(reg_q2514 AND symb_decoder(16#35#)) OR
 					(reg_q2516 AND symb_decoder(16#38#)) OR
 					(reg_q2516 AND symb_decoder(16#34#)) OR
 					(reg_q2516 AND symb_decoder(16#30#)) OR
 					(reg_q2516 AND symb_decoder(16#37#)) OR
 					(reg_q2516 AND symb_decoder(16#32#)) OR
 					(reg_q2516 AND symb_decoder(16#36#)) OR
 					(reg_q2516 AND symb_decoder(16#35#)) OR
 					(reg_q2516 AND symb_decoder(16#31#)) OR
 					(reg_q2516 AND symb_decoder(16#33#)) OR
 					(reg_q2516 AND symb_decoder(16#39#));
reg_q2516_init <= '0' ;
	p_reg_q2516: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2516 <= reg_q2516_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2516 <= reg_q2516_init;
        else
          reg_q2516 <= reg_q2516_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2530_in <= (reg_q2530 AND symb_decoder(16#30#)) OR
 					(reg_q2530 AND symb_decoder(16#33#)) OR
 					(reg_q2530 AND symb_decoder(16#34#)) OR
 					(reg_q2530 AND symb_decoder(16#36#)) OR
 					(reg_q2530 AND symb_decoder(16#38#)) OR
 					(reg_q2530 AND symb_decoder(16#32#)) OR
 					(reg_q2530 AND symb_decoder(16#31#)) OR
 					(reg_q2530 AND symb_decoder(16#35#)) OR
 					(reg_q2530 AND symb_decoder(16#37#)) OR
 					(reg_q2530 AND symb_decoder(16#39#)) OR
 					(reg_q2528 AND symb_decoder(16#39#)) OR
 					(reg_q2528 AND symb_decoder(16#37#)) OR
 					(reg_q2528 AND symb_decoder(16#32#)) OR
 					(reg_q2528 AND symb_decoder(16#38#)) OR
 					(reg_q2528 AND symb_decoder(16#34#)) OR
 					(reg_q2528 AND symb_decoder(16#33#)) OR
 					(reg_q2528 AND symb_decoder(16#35#)) OR
 					(reg_q2528 AND symb_decoder(16#31#)) OR
 					(reg_q2528 AND symb_decoder(16#30#)) OR
 					(reg_q2528 AND symb_decoder(16#36#));
reg_q2530_init <= '0' ;
	p_reg_q2530: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2530 <= reg_q2530_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2530 <= reg_q2530_init;
        else
          reg_q2530 <= reg_q2530_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q56_in <= (reg_q54 AND symb_decoder(16#6b#)) OR
 					(reg_q54 AND symb_decoder(16#4b#));
reg_q56_init <= '0' ;
	p_reg_q56: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q56 <= reg_q56_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q56 <= reg_q56_init;
        else
          reg_q56 <= reg_q56_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q530_in <= (reg_q530 AND symb_decoder(16#36#)) OR
 					(reg_q530 AND symb_decoder(16#33#)) OR
 					(reg_q530 AND symb_decoder(16#35#)) OR
 					(reg_q530 AND symb_decoder(16#38#)) OR
 					(reg_q530 AND symb_decoder(16#39#)) OR
 					(reg_q530 AND symb_decoder(16#30#)) OR
 					(reg_q530 AND symb_decoder(16#34#)) OR
 					(reg_q530 AND symb_decoder(16#37#)) OR
 					(reg_q530 AND symb_decoder(16#31#)) OR
 					(reg_q530 AND symb_decoder(16#32#)) OR
 					(reg_q528 AND symb_decoder(16#39#)) OR
 					(reg_q528 AND symb_decoder(16#35#)) OR
 					(reg_q528 AND symb_decoder(16#38#)) OR
 					(reg_q528 AND symb_decoder(16#36#)) OR
 					(reg_q528 AND symb_decoder(16#34#)) OR
 					(reg_q528 AND symb_decoder(16#32#)) OR
 					(reg_q528 AND symb_decoder(16#33#)) OR
 					(reg_q528 AND symb_decoder(16#31#)) OR
 					(reg_q528 AND symb_decoder(16#37#)) OR
 					(reg_q528 AND symb_decoder(16#30#));
reg_q530_init <= '0' ;
	p_reg_q530: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q530 <= reg_q530_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q530 <= reg_q530_init;
        else
          reg_q530 <= reg_q530_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1603_in <= (reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q1603 AND symb_decoder(16#d6#)) OR
 					(reg_q1603 AND symb_decoder(16#75#)) OR
 					(reg_q1603 AND symb_decoder(16#b9#)) OR
 					(reg_q1603 AND symb_decoder(16#c3#)) OR
 					(reg_q1603 AND symb_decoder(16#b2#)) OR
 					(reg_q1603 AND symb_decoder(16#dd#)) OR
 					(reg_q1603 AND symb_decoder(16#7c#)) OR
 					(reg_q1603 AND symb_decoder(16#d0#)) OR
 					(reg_q1603 AND symb_decoder(16#8a#)) OR
 					(reg_q1603 AND symb_decoder(16#fd#)) OR
 					(reg_q1603 AND symb_decoder(16#e2#)) OR
 					(reg_q1603 AND symb_decoder(16#91#)) OR
 					(reg_q1603 AND symb_decoder(16#ff#)) OR
 					(reg_q1603 AND symb_decoder(16#4b#)) OR
 					(reg_q1603 AND symb_decoder(16#c5#)) OR
 					(reg_q1603 AND symb_decoder(16#3b#)) OR
 					(reg_q1603 AND symb_decoder(16#5f#)) OR
 					(reg_q1603 AND symb_decoder(16#8f#)) OR
 					(reg_q1603 AND symb_decoder(16#0d#)) OR
 					(reg_q1603 AND symb_decoder(16#72#)) OR
 					(reg_q1603 AND symb_decoder(16#34#)) OR
 					(reg_q1603 AND symb_decoder(16#30#)) OR
 					(reg_q1603 AND symb_decoder(16#ac#)) OR
 					(reg_q1603 AND symb_decoder(16#f7#)) OR
 					(reg_q1603 AND symb_decoder(16#5e#)) OR
 					(reg_q1603 AND symb_decoder(16#77#)) OR
 					(reg_q1603 AND symb_decoder(16#d8#)) OR
 					(reg_q1603 AND symb_decoder(16#48#)) OR
 					(reg_q1603 AND symb_decoder(16#61#)) OR
 					(reg_q1603 AND symb_decoder(16#1f#)) OR
 					(reg_q1603 AND symb_decoder(16#bf#)) OR
 					(reg_q1603 AND symb_decoder(16#cf#)) OR
 					(reg_q1603 AND symb_decoder(16#8d#)) OR
 					(reg_q1603 AND symb_decoder(16#99#)) OR
 					(reg_q1603 AND symb_decoder(16#81#)) OR
 					(reg_q1603 AND symb_decoder(16#59#)) OR
 					(reg_q1603 AND symb_decoder(16#b1#)) OR
 					(reg_q1603 AND symb_decoder(16#c6#)) OR
 					(reg_q1603 AND symb_decoder(16#a4#)) OR
 					(reg_q1603 AND symb_decoder(16#bb#)) OR
 					(reg_q1603 AND symb_decoder(16#32#)) OR
 					(reg_q1603 AND symb_decoder(16#07#)) OR
 					(reg_q1603 AND symb_decoder(16#44#)) OR
 					(reg_q1603 AND symb_decoder(16#06#)) OR
 					(reg_q1603 AND symb_decoder(16#62#)) OR
 					(reg_q1603 AND symb_decoder(16#19#)) OR
 					(reg_q1603 AND symb_decoder(16#94#)) OR
 					(reg_q1603 AND symb_decoder(16#ba#)) OR
 					(reg_q1603 AND symb_decoder(16#14#)) OR
 					(reg_q1603 AND symb_decoder(16#6f#)) OR
 					(reg_q1603 AND symb_decoder(16#2c#)) OR
 					(reg_q1603 AND symb_decoder(16#82#)) OR
 					(reg_q1603 AND symb_decoder(16#53#)) OR
 					(reg_q1603 AND symb_decoder(16#55#)) OR
 					(reg_q1603 AND symb_decoder(16#a5#)) OR
 					(reg_q1603 AND symb_decoder(16#fa#)) OR
 					(reg_q1603 AND symb_decoder(16#4e#)) OR
 					(reg_q1603 AND symb_decoder(16#1c#)) OR
 					(reg_q1603 AND symb_decoder(16#7d#)) OR
 					(reg_q1603 AND symb_decoder(16#e3#)) OR
 					(reg_q1603 AND symb_decoder(16#f8#)) OR
 					(reg_q1603 AND symb_decoder(16#cb#)) OR
 					(reg_q1603 AND symb_decoder(16#a8#)) OR
 					(reg_q1603 AND symb_decoder(16#56#)) OR
 					(reg_q1603 AND symb_decoder(16#31#)) OR
 					(reg_q1603 AND symb_decoder(16#3c#)) OR
 					(reg_q1603 AND symb_decoder(16#28#)) OR
 					(reg_q1603 AND symb_decoder(16#3f#)) OR
 					(reg_q1603 AND symb_decoder(16#25#)) OR
 					(reg_q1603 AND symb_decoder(16#b3#)) OR
 					(reg_q1603 AND symb_decoder(16#58#)) OR
 					(reg_q1603 AND symb_decoder(16#96#)) OR
 					(reg_q1603 AND symb_decoder(16#54#)) OR
 					(reg_q1603 AND symb_decoder(16#7f#)) OR
 					(reg_q1603 AND symb_decoder(16#79#)) OR
 					(reg_q1603 AND symb_decoder(16#4d#)) OR
 					(reg_q1603 AND symb_decoder(16#e7#)) OR
 					(reg_q1603 AND symb_decoder(16#c9#)) OR
 					(reg_q1603 AND symb_decoder(16#76#)) OR
 					(reg_q1603 AND symb_decoder(16#bd#)) OR
 					(reg_q1603 AND symb_decoder(16#83#)) OR
 					(reg_q1603 AND symb_decoder(16#d3#)) OR
 					(reg_q1603 AND symb_decoder(16#84#)) OR
 					(reg_q1603 AND symb_decoder(16#45#)) OR
 					(reg_q1603 AND symb_decoder(16#6a#)) OR
 					(reg_q1603 AND symb_decoder(16#20#)) OR
 					(reg_q1603 AND symb_decoder(16#90#)) OR
 					(reg_q1603 AND symb_decoder(16#fc#)) OR
 					(reg_q1603 AND symb_decoder(16#33#)) OR
 					(reg_q1603 AND symb_decoder(16#ef#)) OR
 					(reg_q1603 AND symb_decoder(16#71#)) OR
 					(reg_q1603 AND symb_decoder(16#c1#)) OR
 					(reg_q1603 AND symb_decoder(16#70#)) OR
 					(reg_q1603 AND symb_decoder(16#b5#)) OR
 					(reg_q1603 AND symb_decoder(16#f9#)) OR
 					(reg_q1603 AND symb_decoder(16#65#)) OR
 					(reg_q1603 AND symb_decoder(16#92#)) OR
 					(reg_q1603 AND symb_decoder(16#8b#)) OR
 					(reg_q1603 AND symb_decoder(16#c4#)) OR
 					(reg_q1603 AND symb_decoder(16#89#)) OR
 					(reg_q1603 AND symb_decoder(16#9f#)) OR
 					(reg_q1603 AND symb_decoder(16#2b#)) OR
 					(reg_q1603 AND symb_decoder(16#12#)) OR
 					(reg_q1603 AND symb_decoder(16#d5#)) OR
 					(reg_q1603 AND symb_decoder(16#ee#)) OR
 					(reg_q1603 AND symb_decoder(16#b8#)) OR
 					(reg_q1603 AND symb_decoder(16#0a#)) OR
 					(reg_q1603 AND symb_decoder(16#52#)) OR
 					(reg_q1603 AND symb_decoder(16#f0#)) OR
 					(reg_q1603 AND symb_decoder(16#d9#)) OR
 					(reg_q1603 AND symb_decoder(16#1e#)) OR
 					(reg_q1603 AND symb_decoder(16#3e#)) OR
 					(reg_q1603 AND symb_decoder(16#c0#)) OR
 					(reg_q1603 AND symb_decoder(16#13#)) OR
 					(reg_q1603 AND symb_decoder(16#49#)) OR
 					(reg_q1603 AND symb_decoder(16#57#)) OR
 					(reg_q1603 AND symb_decoder(16#4c#)) OR
 					(reg_q1603 AND symb_decoder(16#67#)) OR
 					(reg_q1603 AND symb_decoder(16#9c#)) OR
 					(reg_q1603 AND symb_decoder(16#c7#)) OR
 					(reg_q1603 AND symb_decoder(16#a9#)) OR
 					(reg_q1603 AND symb_decoder(16#47#)) OR
 					(reg_q1603 AND symb_decoder(16#2d#)) OR
 					(reg_q1603 AND symb_decoder(16#ae#)) OR
 					(reg_q1603 AND symb_decoder(16#ad#)) OR
 					(reg_q1603 AND symb_decoder(16#97#)) OR
 					(reg_q1603 AND symb_decoder(16#0e#)) OR
 					(reg_q1603 AND symb_decoder(16#08#)) OR
 					(reg_q1603 AND symb_decoder(16#98#)) OR
 					(reg_q1603 AND symb_decoder(16#00#)) OR
 					(reg_q1603 AND symb_decoder(16#a0#)) OR
 					(reg_q1603 AND symb_decoder(16#17#)) OR
 					(reg_q1603 AND symb_decoder(16#43#)) OR
 					(reg_q1603 AND symb_decoder(16#f1#)) OR
 					(reg_q1603 AND symb_decoder(16#fb#)) OR
 					(reg_q1603 AND symb_decoder(16#c8#)) OR
 					(reg_q1603 AND symb_decoder(16#39#)) OR
 					(reg_q1603 AND symb_decoder(16#35#)) OR
 					(reg_q1603 AND symb_decoder(16#6e#)) OR
 					(reg_q1603 AND symb_decoder(16#8e#)) OR
 					(reg_q1603 AND symb_decoder(16#e1#)) OR
 					(reg_q1603 AND symb_decoder(16#ec#)) OR
 					(reg_q1603 AND symb_decoder(16#d4#)) OR
 					(reg_q1603 AND symb_decoder(16#1a#)) OR
 					(reg_q1603 AND symb_decoder(16#a7#)) OR
 					(reg_q1603 AND symb_decoder(16#37#)) OR
 					(reg_q1603 AND symb_decoder(16#7e#)) OR
 					(reg_q1603 AND symb_decoder(16#bc#)) OR
 					(reg_q1603 AND symb_decoder(16#e4#)) OR
 					(reg_q1603 AND symb_decoder(16#64#)) OR
 					(reg_q1603 AND symb_decoder(16#6c#)) OR
 					(reg_q1603 AND symb_decoder(16#21#)) OR
 					(reg_q1603 AND symb_decoder(16#d2#)) OR
 					(reg_q1603 AND symb_decoder(16#38#)) OR
 					(reg_q1603 AND symb_decoder(16#36#)) OR
 					(reg_q1603 AND symb_decoder(16#7b#)) OR
 					(reg_q1603 AND symb_decoder(16#9a#)) OR
 					(reg_q1603 AND symb_decoder(16#26#)) OR
 					(reg_q1603 AND symb_decoder(16#6d#)) OR
 					(reg_q1603 AND symb_decoder(16#2f#)) OR
 					(reg_q1603 AND symb_decoder(16#74#)) OR
 					(reg_q1603 AND symb_decoder(16#e9#)) OR
 					(reg_q1603 AND symb_decoder(16#95#)) OR
 					(reg_q1603 AND symb_decoder(16#23#)) OR
 					(reg_q1603 AND symb_decoder(16#ab#)) OR
 					(reg_q1603 AND symb_decoder(16#24#)) OR
 					(reg_q1603 AND symb_decoder(16#df#)) OR
 					(reg_q1603 AND symb_decoder(16#c2#)) OR
 					(reg_q1603 AND symb_decoder(16#e5#)) OR
 					(reg_q1603 AND symb_decoder(16#a2#)) OR
 					(reg_q1603 AND symb_decoder(16#02#)) OR
 					(reg_q1603 AND symb_decoder(16#68#)) OR
 					(reg_q1603 AND symb_decoder(16#69#)) OR
 					(reg_q1603 AND symb_decoder(16#cc#)) OR
 					(reg_q1603 AND symb_decoder(16#af#)) OR
 					(reg_q1603 AND symb_decoder(16#03#)) OR
 					(reg_q1603 AND symb_decoder(16#0c#)) OR
 					(reg_q1603 AND symb_decoder(16#09#)) OR
 					(reg_q1603 AND symb_decoder(16#88#)) OR
 					(reg_q1603 AND symb_decoder(16#41#)) OR
 					(reg_q1603 AND symb_decoder(16#11#)) OR
 					(reg_q1603 AND symb_decoder(16#5c#)) OR
 					(reg_q1603 AND symb_decoder(16#f2#)) OR
 					(reg_q1603 AND symb_decoder(16#db#)) OR
 					(reg_q1603 AND symb_decoder(16#66#)) OR
 					(reg_q1603 AND symb_decoder(16#50#)) OR
 					(reg_q1603 AND symb_decoder(16#fe#)) OR
 					(reg_q1603 AND symb_decoder(16#2e#)) OR
 					(reg_q1603 AND symb_decoder(16#3d#)) OR
 					(reg_q1603 AND symb_decoder(16#3a#)) OR
 					(reg_q1603 AND symb_decoder(16#e6#)) OR
 					(reg_q1603 AND symb_decoder(16#51#)) OR
 					(reg_q1603 AND symb_decoder(16#0b#)) OR
 					(reg_q1603 AND symb_decoder(16#da#)) OR
 					(reg_q1603 AND symb_decoder(16#80#)) OR
 					(reg_q1603 AND symb_decoder(16#d1#)) OR
 					(reg_q1603 AND symb_decoder(16#29#)) OR
 					(reg_q1603 AND symb_decoder(16#4a#)) OR
 					(reg_q1603 AND symb_decoder(16#01#)) OR
 					(reg_q1603 AND symb_decoder(16#5a#)) OR
 					(reg_q1603 AND symb_decoder(16#87#)) OR
 					(reg_q1603 AND symb_decoder(16#1d#)) OR
 					(reg_q1603 AND symb_decoder(16#46#)) OR
 					(reg_q1603 AND symb_decoder(16#40#)) OR
 					(reg_q1603 AND symb_decoder(16#f4#)) OR
 					(reg_q1603 AND symb_decoder(16#9e#)) OR
 					(reg_q1603 AND symb_decoder(16#8c#)) OR
 					(reg_q1603 AND symb_decoder(16#b7#)) OR
 					(reg_q1603 AND symb_decoder(16#f5#)) OR
 					(reg_q1603 AND symb_decoder(16#42#)) OR
 					(reg_q1603 AND symb_decoder(16#ca#)) OR
 					(reg_q1603 AND symb_decoder(16#15#)) OR
 					(reg_q1603 AND symb_decoder(16#f6#)) OR
 					(reg_q1603 AND symb_decoder(16#ce#)) OR
 					(reg_q1603 AND symb_decoder(16#9d#)) OR
 					(reg_q1603 AND symb_decoder(16#a1#)) OR
 					(reg_q1603 AND symb_decoder(16#e0#)) OR
 					(reg_q1603 AND symb_decoder(16#04#)) OR
 					(reg_q1603 AND symb_decoder(16#f3#)) OR
 					(reg_q1603 AND symb_decoder(16#eb#)) OR
 					(reg_q1603 AND symb_decoder(16#dc#)) OR
 					(reg_q1603 AND symb_decoder(16#18#)) OR
 					(reg_q1603 AND symb_decoder(16#0f#)) OR
 					(reg_q1603 AND symb_decoder(16#78#)) OR
 					(reg_q1603 AND symb_decoder(16#85#)) OR
 					(reg_q1603 AND symb_decoder(16#a6#)) OR
 					(reg_q1603 AND symb_decoder(16#a3#)) OR
 					(reg_q1603 AND symb_decoder(16#e8#)) OR
 					(reg_q1603 AND symb_decoder(16#93#)) OR
 					(reg_q1603 AND symb_decoder(16#4f#)) OR
 					(reg_q1603 AND symb_decoder(16#ed#)) OR
 					(reg_q1603 AND symb_decoder(16#de#)) OR
 					(reg_q1603 AND symb_decoder(16#5d#)) OR
 					(reg_q1603 AND symb_decoder(16#63#)) OR
 					(reg_q1603 AND symb_decoder(16#16#)) OR
 					(reg_q1603 AND symb_decoder(16#60#)) OR
 					(reg_q1603 AND symb_decoder(16#05#)) OR
 					(reg_q1603 AND symb_decoder(16#86#)) OR
 					(reg_q1603 AND symb_decoder(16#10#)) OR
 					(reg_q1603 AND symb_decoder(16#d7#)) OR
 					(reg_q1603 AND symb_decoder(16#2a#)) OR
 					(reg_q1603 AND symb_decoder(16#5b#)) OR
 					(reg_q1603 AND symb_decoder(16#be#)) OR
 					(reg_q1603 AND symb_decoder(16#aa#)) OR
 					(reg_q1603 AND symb_decoder(16#b4#)) OR
 					(reg_q1603 AND symb_decoder(16#b6#)) OR
 					(reg_q1603 AND symb_decoder(16#9b#)) OR
 					(reg_q1603 AND symb_decoder(16#1b#)) OR
 					(reg_q1603 AND symb_decoder(16#6b#)) OR
 					(reg_q1603 AND symb_decoder(16#b0#)) OR
 					(reg_q1603 AND symb_decoder(16#cd#)) OR
 					(reg_q1603 AND symb_decoder(16#22#)) OR
 					(reg_q1603 AND symb_decoder(16#7a#)) OR
 					(reg_q1603 AND symb_decoder(16#ea#)) OR
 					(reg_q1603 AND symb_decoder(16#27#)) OR
 					(reg_q1603 AND symb_decoder(16#73#));
reg_q1603_init <= '0' ;
	p_reg_q1603: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1603 <= reg_q1603_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1603 <= reg_q1603_init;
        else
          reg_q1603 <= reg_q1603_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q907_in <= (reg_q905 AND symb_decoder(16#4a#)) OR
 					(reg_q905 AND symb_decoder(16#6a#));
reg_q907_init <= '0' ;
	p_reg_q907: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q907 <= reg_q907_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q907 <= reg_q907_init;
        else
          reg_q907 <= reg_q907_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q909_in <= (reg_q907 AND symb_decoder(16#55#)) OR
 					(reg_q907 AND symb_decoder(16#75#));
reg_q909_init <= '0' ;
	p_reg_q909: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q909 <= reg_q909_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q909 <= reg_q909_init;
        else
          reg_q909 <= reg_q909_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q610_in <= (reg_q608 AND symb_decoder(16#25#));
reg_q610_init <= '0' ;
	p_reg_q610: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q610 <= reg_q610_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q610 <= reg_q610_init;
        else
          reg_q610 <= reg_q610_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q612_in <= (reg_q610 AND symb_decoder(16#32#));
reg_q612_init <= '0' ;
	p_reg_q612: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q612 <= reg_q612_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q612 <= reg_q612_init;
        else
          reg_q612 <= reg_q612_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1462_in <= (reg_q1462 AND symb_decoder(16#20#)) OR
 					(reg_q1462 AND symb_decoder(16#0c#)) OR
 					(reg_q1462 AND symb_decoder(16#09#)) OR
 					(reg_q1462 AND symb_decoder(16#0a#)) OR
 					(reg_q1462 AND symb_decoder(16#0d#)) OR
 					(reg_q1460 AND symb_decoder(16#09#)) OR
 					(reg_q1460 AND symb_decoder(16#0a#)) OR
 					(reg_q1460 AND symb_decoder(16#0d#)) OR
 					(reg_q1460 AND symb_decoder(16#20#)) OR
 					(reg_q1460 AND symb_decoder(16#0c#));
reg_q1462_init <= '0' ;
	p_reg_q1462: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1462 <= reg_q1462_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1462 <= reg_q1462_init;
        else
          reg_q1462 <= reg_q1462_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q123_in <= (reg_q121 AND symb_decoder(16#35#)) OR
 					(reg_q121 AND symb_decoder(16#32#)) OR
 					(reg_q121 AND symb_decoder(16#38#)) OR
 					(reg_q121 AND symb_decoder(16#31#)) OR
 					(reg_q121 AND symb_decoder(16#30#)) OR
 					(reg_q121 AND symb_decoder(16#36#)) OR
 					(reg_q121 AND symb_decoder(16#39#)) OR
 					(reg_q121 AND symb_decoder(16#33#)) OR
 					(reg_q121 AND symb_decoder(16#37#)) OR
 					(reg_q121 AND symb_decoder(16#34#)) OR
 					(reg_q123 AND symb_decoder(16#31#)) OR
 					(reg_q123 AND symb_decoder(16#34#)) OR
 					(reg_q123 AND symb_decoder(16#38#)) OR
 					(reg_q123 AND symb_decoder(16#39#)) OR
 					(reg_q123 AND symb_decoder(16#30#)) OR
 					(reg_q123 AND symb_decoder(16#36#)) OR
 					(reg_q123 AND symb_decoder(16#32#)) OR
 					(reg_q123 AND symb_decoder(16#33#)) OR
 					(reg_q123 AND symb_decoder(16#35#)) OR
 					(reg_q123 AND symb_decoder(16#37#));
reg_q123_init <= '0' ;
	p_reg_q123: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q123 <= reg_q123_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q123 <= reg_q123_init;
        else
          reg_q123 <= reg_q123_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2213_in <= (reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2212 AND symb_decoder(16#77#)) OR
 					(reg_q2212 AND symb_decoder(16#57#));
reg_q2213_init <= '0' ;
	p_reg_q2213: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2213 <= reg_q2213_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2213 <= reg_q2213_init;
        else
          reg_q2213 <= reg_q2213_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q426_in <= (reg_q426 AND symb_decoder(16#20#)) OR
 					(reg_q426 AND symb_decoder(16#0a#)) OR
 					(reg_q426 AND symb_decoder(16#0c#)) OR
 					(reg_q426 AND symb_decoder(16#0d#)) OR
 					(reg_q426 AND symb_decoder(16#09#)) OR
 					(reg_q424 AND symb_decoder(16#0c#)) OR
 					(reg_q424 AND symb_decoder(16#0a#)) OR
 					(reg_q424 AND symb_decoder(16#20#)) OR
 					(reg_q424 AND symb_decoder(16#09#)) OR
 					(reg_q424 AND symb_decoder(16#0d#));
reg_q426_init <= '0' ;
	p_reg_q426: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q426 <= reg_q426_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q426 <= reg_q426_init;
        else
          reg_q426 <= reg_q426_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2405_in <= (reg_q2403 AND symb_decoder(16#62#)) OR
 					(reg_q2403 AND symb_decoder(16#42#));
reg_q2405_init <= '0' ;
	p_reg_q2405: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2405 <= reg_q2405_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2405 <= reg_q2405_init;
        else
          reg_q2405 <= reg_q2405_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2407_in <= (reg_q2405 AND symb_decoder(16#61#)) OR
 					(reg_q2405 AND symb_decoder(16#41#));
reg_q2407_init <= '0' ;
	p_reg_q2407: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2407 <= reg_q2407_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2407 <= reg_q2407_init;
        else
          reg_q2407 <= reg_q2407_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1470_in <= (reg_q1470 AND symb_decoder(16#0d#)) OR
 					(reg_q1470 AND symb_decoder(16#0a#)) OR
 					(reg_q1470 AND symb_decoder(16#09#)) OR
 					(reg_q1470 AND symb_decoder(16#20#)) OR
 					(reg_q1470 AND symb_decoder(16#0c#)) OR
 					(reg_q1468 AND symb_decoder(16#0c#)) OR
 					(reg_q1468 AND symb_decoder(16#20#)) OR
 					(reg_q1468 AND symb_decoder(16#0a#)) OR
 					(reg_q1468 AND symb_decoder(16#09#)) OR
 					(reg_q1468 AND symb_decoder(16#0d#));
reg_q1470_init <= '0' ;
	p_reg_q1470: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1470 <= reg_q1470_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1470 <= reg_q1470_init;
        else
          reg_q1470 <= reg_q1470_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2028_in <= (reg_q2026 AND symb_decoder(16#47#)) OR
 					(reg_q2026 AND symb_decoder(16#67#));
reg_q2028_init <= '0' ;
	p_reg_q2028: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2028 <= reg_q2028_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2028 <= reg_q2028_init;
        else
          reg_q2028 <= reg_q2028_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1217_in <= (reg_q1215 AND symb_decoder(16#65#)) OR
 					(reg_q1215 AND symb_decoder(16#45#));
reg_q1217_init <= '0' ;
	p_reg_q1217: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1217 <= reg_q1217_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1217 <= reg_q1217_init;
        else
          reg_q1217 <= reg_q1217_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1219_in <= (reg_q1217 AND symb_decoder(16#31#)) OR
 					(reg_q1217 AND symb_decoder(16#33#)) OR
 					(reg_q1217 AND symb_decoder(16#34#)) OR
 					(reg_q1217 AND symb_decoder(16#37#)) OR
 					(reg_q1217 AND symb_decoder(16#32#)) OR
 					(reg_q1217 AND symb_decoder(16#39#)) OR
 					(reg_q1217 AND symb_decoder(16#35#)) OR
 					(reg_q1217 AND symb_decoder(16#38#)) OR
 					(reg_q1217 AND symb_decoder(16#36#)) OR
 					(reg_q1217 AND symb_decoder(16#30#)) OR
 					(reg_q1219 AND symb_decoder(16#38#)) OR
 					(reg_q1219 AND symb_decoder(16#36#)) OR
 					(reg_q1219 AND symb_decoder(16#35#)) OR
 					(reg_q1219 AND symb_decoder(16#33#)) OR
 					(reg_q1219 AND symb_decoder(16#39#)) OR
 					(reg_q1219 AND symb_decoder(16#34#)) OR
 					(reg_q1219 AND symb_decoder(16#32#)) OR
 					(reg_q1219 AND symb_decoder(16#31#)) OR
 					(reg_q1219 AND symb_decoder(16#37#)) OR
 					(reg_q1219 AND symb_decoder(16#30#));
reg_q1219_init <= '0' ;
	p_reg_q1219: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1219 <= reg_q1219_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1219 <= reg_q1219_init;
        else
          reg_q1219 <= reg_q1219_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q241_in <= (reg_q241 AND symb_decoder(16#38#)) OR
 					(reg_q241 AND symb_decoder(16#31#)) OR
 					(reg_q241 AND symb_decoder(16#39#)) OR
 					(reg_q241 AND symb_decoder(16#30#)) OR
 					(reg_q241 AND symb_decoder(16#34#)) OR
 					(reg_q241 AND symb_decoder(16#33#)) OR
 					(reg_q241 AND symb_decoder(16#32#)) OR
 					(reg_q241 AND symb_decoder(16#35#)) OR
 					(reg_q241 AND symb_decoder(16#37#)) OR
 					(reg_q241 AND symb_decoder(16#36#)) OR
 					(reg_q239 AND symb_decoder(16#30#)) OR
 					(reg_q239 AND symb_decoder(16#38#)) OR
 					(reg_q239 AND symb_decoder(16#35#)) OR
 					(reg_q239 AND symb_decoder(16#31#)) OR
 					(reg_q239 AND symb_decoder(16#33#)) OR
 					(reg_q239 AND symb_decoder(16#34#)) OR
 					(reg_q239 AND symb_decoder(16#32#)) OR
 					(reg_q239 AND symb_decoder(16#39#)) OR
 					(reg_q239 AND symb_decoder(16#36#)) OR
 					(reg_q239 AND symb_decoder(16#37#));
reg_q241_init <= '0' ;
	p_reg_q241: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q241 <= reg_q241_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q241 <= reg_q241_init;
        else
          reg_q241 <= reg_q241_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1088_in <= (reg_q1086 AND symb_decoder(16#2e#));
reg_q1088_init <= '0' ;
	p_reg_q1088: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1088 <= reg_q1088_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1088 <= reg_q1088_init;
        else
          reg_q1088 <= reg_q1088_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1090_in <= (reg_q1088 AND symb_decoder(16#31#)) OR
 					(reg_q1088 AND symb_decoder(16#33#)) OR
 					(reg_q1088 AND symb_decoder(16#36#)) OR
 					(reg_q1088 AND symb_decoder(16#39#)) OR
 					(reg_q1088 AND symb_decoder(16#38#)) OR
 					(reg_q1088 AND symb_decoder(16#35#)) OR
 					(reg_q1088 AND symb_decoder(16#32#)) OR
 					(reg_q1088 AND symb_decoder(16#37#)) OR
 					(reg_q1088 AND symb_decoder(16#34#)) OR
 					(reg_q1088 AND symb_decoder(16#30#)) OR
 					(reg_q1090 AND symb_decoder(16#38#)) OR
 					(reg_q1090 AND symb_decoder(16#30#)) OR
 					(reg_q1090 AND symb_decoder(16#39#)) OR
 					(reg_q1090 AND symb_decoder(16#32#)) OR
 					(reg_q1090 AND symb_decoder(16#34#)) OR
 					(reg_q1090 AND symb_decoder(16#36#)) OR
 					(reg_q1090 AND symb_decoder(16#37#)) OR
 					(reg_q1090 AND symb_decoder(16#35#)) OR
 					(reg_q1090 AND symb_decoder(16#33#)) OR
 					(reg_q1090 AND symb_decoder(16#31#));
reg_q1090_init <= '0' ;
	p_reg_q1090: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1090 <= reg_q1090_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1090 <= reg_q1090_init;
        else
          reg_q1090 <= reg_q1090_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1991_in <= (reg_q1989 AND symb_decoder(16#2e#));
reg_q1991_init <= '0' ;
	p_reg_q1991: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1991 <= reg_q1991_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1991 <= reg_q1991_init;
        else
          reg_q1991 <= reg_q1991_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1993_in <= (reg_q1991 AND symb_decoder(16#33#)) OR
 					(reg_q1991 AND symb_decoder(16#32#)) OR
 					(reg_q1991 AND symb_decoder(16#34#)) OR
 					(reg_q1991 AND symb_decoder(16#36#)) OR
 					(reg_q1991 AND symb_decoder(16#31#)) OR
 					(reg_q1991 AND symb_decoder(16#37#)) OR
 					(reg_q1991 AND symb_decoder(16#39#)) OR
 					(reg_q1991 AND symb_decoder(16#30#)) OR
 					(reg_q1991 AND symb_decoder(16#35#)) OR
 					(reg_q1991 AND symb_decoder(16#38#)) OR
 					(reg_q1993 AND symb_decoder(16#30#)) OR
 					(reg_q1993 AND symb_decoder(16#38#)) OR
 					(reg_q1993 AND symb_decoder(16#35#)) OR
 					(reg_q1993 AND symb_decoder(16#37#)) OR
 					(reg_q1993 AND symb_decoder(16#34#)) OR
 					(reg_q1993 AND symb_decoder(16#32#)) OR
 					(reg_q1993 AND symb_decoder(16#39#)) OR
 					(reg_q1993 AND symb_decoder(16#36#)) OR
 					(reg_q1993 AND symb_decoder(16#31#)) OR
 					(reg_q1993 AND symb_decoder(16#33#));
reg_q1993_init <= '0' ;
	p_reg_q1993: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1993 <= reg_q1993_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1993 <= reg_q1993_init;
        else
          reg_q1993 <= reg_q1993_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1145_in <= (reg_q1143 AND symb_decoder(16#2e#));
reg_q1145_init <= '0' ;
	p_reg_q1145: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1145 <= reg_q1145_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1145 <= reg_q1145_init;
        else
          reg_q1145 <= reg_q1145_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1147_in <= (reg_q1145 AND symb_decoder(16#37#)) OR
 					(reg_q1145 AND symb_decoder(16#32#)) OR
 					(reg_q1145 AND symb_decoder(16#30#)) OR
 					(reg_q1145 AND symb_decoder(16#36#)) OR
 					(reg_q1145 AND symb_decoder(16#35#)) OR
 					(reg_q1145 AND symb_decoder(16#39#)) OR
 					(reg_q1145 AND symb_decoder(16#34#)) OR
 					(reg_q1145 AND symb_decoder(16#38#)) OR
 					(reg_q1145 AND symb_decoder(16#31#)) OR
 					(reg_q1145 AND symb_decoder(16#33#)) OR
 					(reg_q1147 AND symb_decoder(16#33#)) OR
 					(reg_q1147 AND symb_decoder(16#37#)) OR
 					(reg_q1147 AND symb_decoder(16#36#)) OR
 					(reg_q1147 AND symb_decoder(16#38#)) OR
 					(reg_q1147 AND symb_decoder(16#35#)) OR
 					(reg_q1147 AND symb_decoder(16#30#)) OR
 					(reg_q1147 AND symb_decoder(16#31#)) OR
 					(reg_q1147 AND symb_decoder(16#34#)) OR
 					(reg_q1147 AND symb_decoder(16#39#)) OR
 					(reg_q1147 AND symb_decoder(16#32#));
reg_q1147_init <= '0' ;
	p_reg_q1147: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1147 <= reg_q1147_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1147 <= reg_q1147_init;
        else
          reg_q1147 <= reg_q1147_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1967_in <= (reg_q1965 AND symb_decoder(16#52#)) OR
 					(reg_q1965 AND symb_decoder(16#72#));
reg_q1967_init <= '0' ;
	p_reg_q1967: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1967 <= reg_q1967_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1967 <= reg_q1967_init;
        else
          reg_q1967 <= reg_q1967_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1969_in <= (reg_q1967 AND symb_decoder(16#76#)) OR
 					(reg_q1967 AND symb_decoder(16#56#));
reg_q1969_init <= '0' ;
	p_reg_q1969: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1969 <= reg_q1969_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1969 <= reg_q1969_init;
        else
          reg_q1969 <= reg_q1969_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1106_in <= (reg_q1106 AND symb_decoder(16#0c#)) OR
 					(reg_q1106 AND symb_decoder(16#09#)) OR
 					(reg_q1106 AND symb_decoder(16#0d#)) OR
 					(reg_q1106 AND symb_decoder(16#0a#)) OR
 					(reg_q1106 AND symb_decoder(16#20#)) OR
 					(reg_q1104 AND symb_decoder(16#0d#)) OR
 					(reg_q1104 AND symb_decoder(16#20#)) OR
 					(reg_q1104 AND symb_decoder(16#0c#)) OR
 					(reg_q1104 AND symb_decoder(16#09#)) OR
 					(reg_q1104 AND symb_decoder(16#0a#));
reg_q1106_init <= '0' ;
	p_reg_q1106: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1106 <= reg_q1106_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1106 <= reg_q1106_init;
        else
          reg_q1106 <= reg_q1106_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1205_in <= (reg_q1203 AND symb_decoder(16#6e#)) OR
 					(reg_q1203 AND symb_decoder(16#4e#));
reg_q1205_init <= '0' ;
	p_reg_q1205: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1205 <= reg_q1205_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1205 <= reg_q1205_init;
        else
          reg_q1205 <= reg_q1205_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q524_in <= (reg_q522 AND symb_decoder(16#2e#));
reg_q524_init <= '0' ;
	p_reg_q524: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q524 <= reg_q524_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q524 <= reg_q524_init;
        else
          reg_q524 <= reg_q524_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q526_in <= (reg_q524 AND symb_decoder(16#35#)) OR
 					(reg_q524 AND symb_decoder(16#33#)) OR
 					(reg_q524 AND symb_decoder(16#30#)) OR
 					(reg_q524 AND symb_decoder(16#32#)) OR
 					(reg_q524 AND symb_decoder(16#31#)) OR
 					(reg_q524 AND symb_decoder(16#34#)) OR
 					(reg_q524 AND symb_decoder(16#37#)) OR
 					(reg_q524 AND symb_decoder(16#39#)) OR
 					(reg_q524 AND symb_decoder(16#36#)) OR
 					(reg_q524 AND symb_decoder(16#38#)) OR
 					(reg_q526 AND symb_decoder(16#31#)) OR
 					(reg_q526 AND symb_decoder(16#37#)) OR
 					(reg_q526 AND symb_decoder(16#34#)) OR
 					(reg_q526 AND symb_decoder(16#39#)) OR
 					(reg_q526 AND symb_decoder(16#38#)) OR
 					(reg_q526 AND symb_decoder(16#36#)) OR
 					(reg_q526 AND symb_decoder(16#30#)) OR
 					(reg_q526 AND symb_decoder(16#32#)) OR
 					(reg_q526 AND symb_decoder(16#35#)) OR
 					(reg_q526 AND symb_decoder(16#33#));
reg_q526_init <= '0' ;
	p_reg_q526: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q526 <= reg_q526_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q526 <= reg_q526_init;
        else
          reg_q526 <= reg_q526_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1468_in <= (reg_q1466 AND symb_decoder(16#45#)) OR
 					(reg_q1466 AND symb_decoder(16#65#));
reg_q1468_init <= '0' ;
	p_reg_q1468: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1468 <= reg_q1468_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1468 <= reg_q1468_init;
        else
          reg_q1468 <= reg_q1468_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1672_in <= (reg_q1670 AND symb_decoder(16#3b#));
reg_q1672_init <= '0' ;
	p_reg_q1672: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1672 <= reg_q1672_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1672 <= reg_q1672_init;
        else
          reg_q1672 <= reg_q1672_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1674_in <= (reg_q1672 AND symb_decoder(16#0d#)) OR
 					(reg_q1672 AND symb_decoder(16#20#)) OR
 					(reg_q1672 AND symb_decoder(16#0a#)) OR
 					(reg_q1672 AND symb_decoder(16#09#)) OR
 					(reg_q1672 AND symb_decoder(16#0c#)) OR
 					(reg_q1674 AND symb_decoder(16#0d#)) OR
 					(reg_q1674 AND symb_decoder(16#0a#)) OR
 					(reg_q1674 AND symb_decoder(16#20#)) OR
 					(reg_q1674 AND symb_decoder(16#0c#)) OR
 					(reg_q1674 AND symb_decoder(16#09#));
reg_q1674_init <= '0' ;
	p_reg_q1674: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1674 <= reg_q1674_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1674 <= reg_q1674_init;
        else
          reg_q1674 <= reg_q1674_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2375_in <= (reg_q2373 AND symb_decoder(16#2e#));
reg_q2375_init <= '0' ;
	p_reg_q2375: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2375 <= reg_q2375_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2375 <= reg_q2375_init;
        else
          reg_q2375 <= reg_q2375_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2377_in <= (reg_q2375 AND symb_decoder(16#34#)) OR
 					(reg_q2375 AND symb_decoder(16#39#)) OR
 					(reg_q2375 AND symb_decoder(16#35#)) OR
 					(reg_q2375 AND symb_decoder(16#33#)) OR
 					(reg_q2375 AND symb_decoder(16#32#)) OR
 					(reg_q2375 AND symb_decoder(16#31#)) OR
 					(reg_q2375 AND symb_decoder(16#38#)) OR
 					(reg_q2375 AND symb_decoder(16#30#)) OR
 					(reg_q2375 AND symb_decoder(16#36#)) OR
 					(reg_q2375 AND symb_decoder(16#37#)) OR
 					(reg_q2377 AND symb_decoder(16#31#)) OR
 					(reg_q2377 AND symb_decoder(16#32#)) OR
 					(reg_q2377 AND symb_decoder(16#36#)) OR
 					(reg_q2377 AND symb_decoder(16#30#)) OR
 					(reg_q2377 AND symb_decoder(16#38#)) OR
 					(reg_q2377 AND symb_decoder(16#35#)) OR
 					(reg_q2377 AND symb_decoder(16#33#)) OR
 					(reg_q2377 AND symb_decoder(16#39#)) OR
 					(reg_q2377 AND symb_decoder(16#34#)) OR
 					(reg_q2377 AND symb_decoder(16#37#));
reg_q2377_init <= '0' ;
	p_reg_q2377: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2377 <= reg_q2377_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2377 <= reg_q2377_init;
        else
          reg_q2377 <= reg_q2377_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q173_in <= (reg_q171 AND symb_decoder(16#79#)) OR
 					(reg_q171 AND symb_decoder(16#59#));
reg_q173_init <= '0' ;
	p_reg_q173: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q173 <= reg_q173_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q173 <= reg_q173_init;
        else
          reg_q173 <= reg_q173_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q175_in <= (reg_q173 AND symb_decoder(16#21#));
reg_q175_init <= '0' ;
	p_reg_q175: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q175 <= reg_q175_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q175 <= reg_q175_init;
        else
          reg_q175 <= reg_q175_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q309_in <= (reg_q307 AND symb_decoder(16#73#)) OR
 					(reg_q307 AND symb_decoder(16#53#));
reg_q309_init <= '0' ;
	p_reg_q309: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q309 <= reg_q309_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q309 <= reg_q309_init;
        else
          reg_q309 <= reg_q309_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q311_in <= (reg_q309 AND symb_decoder(16#57#)) OR
 					(reg_q309 AND symb_decoder(16#77#));
reg_q311_init <= '0' ;
	p_reg_q311: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q311 <= reg_q311_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q311 <= reg_q311_init;
        else
          reg_q311 <= reg_q311_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1421_in <= (reg_q1419 AND symb_decoder(16#70#)) OR
 					(reg_q1419 AND symb_decoder(16#50#));
reg_q1421_init <= '0' ;
	p_reg_q1421: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1421 <= reg_q1421_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1421 <= reg_q1421_init;
        else
          reg_q1421 <= reg_q1421_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1423_in <= (reg_q1421 AND symb_decoder(16#45#)) OR
 					(reg_q1421 AND symb_decoder(16#65#));
reg_q1423_init <= '0' ;
	p_reg_q1423: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1423 <= reg_q1423_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1423 <= reg_q1423_init;
        else
          reg_q1423 <= reg_q1423_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q803_in <= (reg_q801 AND symb_decoder(16#2e#));
reg_q803_init <= '0' ;
	p_reg_q803: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q803 <= reg_q803_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q803 <= reg_q803_init;
        else
          reg_q803 <= reg_q803_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q805_in <= (reg_q803 AND symb_decoder(16#38#)) OR
 					(reg_q803 AND symb_decoder(16#32#)) OR
 					(reg_q803 AND symb_decoder(16#36#)) OR
 					(reg_q803 AND symb_decoder(16#30#)) OR
 					(reg_q803 AND symb_decoder(16#34#)) OR
 					(reg_q803 AND symb_decoder(16#33#)) OR
 					(reg_q803 AND symb_decoder(16#39#)) OR
 					(reg_q803 AND symb_decoder(16#31#)) OR
 					(reg_q803 AND symb_decoder(16#37#)) OR
 					(reg_q803 AND symb_decoder(16#35#)) OR
 					(reg_q805 AND symb_decoder(16#30#)) OR
 					(reg_q805 AND symb_decoder(16#34#)) OR
 					(reg_q805 AND symb_decoder(16#39#)) OR
 					(reg_q805 AND symb_decoder(16#38#)) OR
 					(reg_q805 AND symb_decoder(16#36#)) OR
 					(reg_q805 AND symb_decoder(16#32#)) OR
 					(reg_q805 AND symb_decoder(16#31#)) OR
 					(reg_q805 AND symb_decoder(16#35#)) OR
 					(reg_q805 AND symb_decoder(16#37#)) OR
 					(reg_q805 AND symb_decoder(16#33#));
reg_q805_init <= '0' ;
	p_reg_q805: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q805 <= reg_q805_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q805 <= reg_q805_init;
        else
          reg_q805 <= reg_q805_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1335_in <= (reg_q1335 AND symb_decoder(16#35#)) OR
 					(reg_q1335 AND symb_decoder(16#39#)) OR
 					(reg_q1335 AND symb_decoder(16#32#)) OR
 					(reg_q1335 AND symb_decoder(16#34#)) OR
 					(reg_q1335 AND symb_decoder(16#30#)) OR
 					(reg_q1335 AND symb_decoder(16#36#)) OR
 					(reg_q1335 AND symb_decoder(16#33#)) OR
 					(reg_q1335 AND symb_decoder(16#37#)) OR
 					(reg_q1335 AND symb_decoder(16#38#)) OR
 					(reg_q1335 AND symb_decoder(16#31#)) OR
 					(reg_q1333 AND symb_decoder(16#38#)) OR
 					(reg_q1333 AND symb_decoder(16#35#)) OR
 					(reg_q1333 AND symb_decoder(16#31#)) OR
 					(reg_q1333 AND symb_decoder(16#39#)) OR
 					(reg_q1333 AND symb_decoder(16#32#)) OR
 					(reg_q1333 AND symb_decoder(16#33#)) OR
 					(reg_q1333 AND symb_decoder(16#34#)) OR
 					(reg_q1333 AND symb_decoder(16#37#)) OR
 					(reg_q1333 AND symb_decoder(16#30#)) OR
 					(reg_q1333 AND symb_decoder(16#36#));
reg_q1335_init <= '0' ;
	p_reg_q1335: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1335 <= reg_q1335_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1335 <= reg_q1335_init;
        else
          reg_q1335 <= reg_q1335_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2229_in <= (reg_q2229 AND symb_decoder(16#0c#)) OR
 					(reg_q2229 AND symb_decoder(16#0a#)) OR
 					(reg_q2229 AND symb_decoder(16#20#)) OR
 					(reg_q2229 AND symb_decoder(16#0d#)) OR
 					(reg_q2229 AND symb_decoder(16#09#)) OR
 					(reg_q2227 AND symb_decoder(16#20#)) OR
 					(reg_q2227 AND symb_decoder(16#0a#)) OR
 					(reg_q2227 AND symb_decoder(16#09#)) OR
 					(reg_q2227 AND symb_decoder(16#0c#)) OR
 					(reg_q2227 AND symb_decoder(16#0d#));
reg_q2229_init <= '0' ;
	p_reg_q2229: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2229 <= reg_q2229_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2229 <= reg_q2229_init;
        else
          reg_q2229 <= reg_q2229_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2093_in <= (reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2092 AND symb_decoder(16#55#)) OR
 					(reg_q2092 AND symb_decoder(16#75#));
reg_q2093_init <= '0' ;
	p_reg_q2093: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2093 <= reg_q2093_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2093 <= reg_q2093_init;
        else
          reg_q2093 <= reg_q2093_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1983_in <= (reg_q1981 AND symb_decoder(16#2e#));
reg_q1983_init <= '0' ;
	p_reg_q1983: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1983 <= reg_q1983_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1983 <= reg_q1983_init;
        else
          reg_q1983 <= reg_q1983_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1985_in <= (reg_q1983 AND symb_decoder(16#30#)) OR
 					(reg_q1983 AND symb_decoder(16#33#)) OR
 					(reg_q1983 AND symb_decoder(16#37#)) OR
 					(reg_q1983 AND symb_decoder(16#35#)) OR
 					(reg_q1983 AND symb_decoder(16#39#)) OR
 					(reg_q1983 AND symb_decoder(16#38#)) OR
 					(reg_q1983 AND symb_decoder(16#36#)) OR
 					(reg_q1983 AND symb_decoder(16#34#)) OR
 					(reg_q1983 AND symb_decoder(16#31#)) OR
 					(reg_q1983 AND symb_decoder(16#32#)) OR
 					(reg_q1985 AND symb_decoder(16#38#)) OR
 					(reg_q1985 AND symb_decoder(16#37#)) OR
 					(reg_q1985 AND symb_decoder(16#36#)) OR
 					(reg_q1985 AND symb_decoder(16#31#)) OR
 					(reg_q1985 AND symb_decoder(16#32#)) OR
 					(reg_q1985 AND symb_decoder(16#35#)) OR
 					(reg_q1985 AND symb_decoder(16#34#)) OR
 					(reg_q1985 AND symb_decoder(16#30#)) OR
 					(reg_q1985 AND symb_decoder(16#39#)) OR
 					(reg_q1985 AND symb_decoder(16#33#));
reg_q1985_init <= '0' ;
	p_reg_q1985: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1985 <= reg_q1985_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1985 <= reg_q1985_init;
        else
          reg_q1985 <= reg_q1985_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1425_in <= (reg_q1423 AND symb_decoder(16#72#)) OR
 					(reg_q1423 AND symb_decoder(16#52#));
reg_q1425_init <= '0' ;
	p_reg_q1425: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1425 <= reg_q1425_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1425 <= reg_q1425_init;
        else
          reg_q1425 <= reg_q1425_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q129_in <= (reg_q127 AND symb_decoder(16#0c#)) OR
 					(reg_q127 AND symb_decoder(16#09#)) OR
 					(reg_q127 AND symb_decoder(16#20#)) OR
 					(reg_q127 AND symb_decoder(16#0d#)) OR
 					(reg_q127 AND symb_decoder(16#0a#)) OR
 					(reg_q129 AND symb_decoder(16#0c#)) OR
 					(reg_q129 AND symb_decoder(16#0d#)) OR
 					(reg_q129 AND symb_decoder(16#20#)) OR
 					(reg_q129 AND symb_decoder(16#0a#)) OR
 					(reg_q129 AND symb_decoder(16#09#));
reg_q129_init <= '0' ;
	p_reg_q129: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q129 <= reg_q129_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q129 <= reg_q129_init;
        else
          reg_q129 <= reg_q129_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1866_in <= (reg_q1864 AND symb_decoder(16#2e#));
reg_q1866_init <= '0' ;
	p_reg_q1866: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1866 <= reg_q1866_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1866 <= reg_q1866_init;
        else
          reg_q1866 <= reg_q1866_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1868_in <= (reg_q1866 AND symb_decoder(16#0a#)) OR
 					(reg_q1866 AND symb_decoder(16#0c#)) OR
 					(reg_q1866 AND symb_decoder(16#0d#)) OR
 					(reg_q1866 AND symb_decoder(16#20#)) OR
 					(reg_q1866 AND symb_decoder(16#09#)) OR
 					(reg_q1868 AND symb_decoder(16#0a#)) OR
 					(reg_q1868 AND symb_decoder(16#0c#)) OR
 					(reg_q1868 AND symb_decoder(16#0d#)) OR
 					(reg_q1868 AND symb_decoder(16#09#)) OR
 					(reg_q1868 AND symb_decoder(16#20#));
reg_q1868_init <= '0' ;
	p_reg_q1868: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1868 <= reg_q1868_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1868 <= reg_q1868_init;
        else
          reg_q1868 <= reg_q1868_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2066_in <= (reg_q2066 AND symb_decoder(16#09#)) OR
 					(reg_q2066 AND symb_decoder(16#0a#)) OR
 					(reg_q2066 AND symb_decoder(16#0d#)) OR
 					(reg_q2066 AND symb_decoder(16#0c#)) OR
 					(reg_q2066 AND symb_decoder(16#20#)) OR
 					(reg_q2064 AND symb_decoder(16#20#)) OR
 					(reg_q2064 AND symb_decoder(16#09#)) OR
 					(reg_q2064 AND symb_decoder(16#0d#)) OR
 					(reg_q2064 AND symb_decoder(16#0a#)) OR
 					(reg_q2064 AND symb_decoder(16#0c#));
reg_q2066_init <= '0' ;
	p_reg_q2066: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2066 <= reg_q2066_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2066 <= reg_q2066_init;
        else
          reg_q2066 <= reg_q2066_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1341_in <= (reg_q1341 AND symb_decoder(16#0a#)) OR
 					(reg_q1341 AND symb_decoder(16#0d#)) OR
 					(reg_q1341 AND symb_decoder(16#0c#)) OR
 					(reg_q1341 AND symb_decoder(16#20#)) OR
 					(reg_q1341 AND symb_decoder(16#09#)) OR
 					(reg_q1339 AND symb_decoder(16#09#)) OR
 					(reg_q1339 AND symb_decoder(16#0a#)) OR
 					(reg_q1339 AND symb_decoder(16#0d#)) OR
 					(reg_q1339 AND symb_decoder(16#0c#)) OR
 					(reg_q1339 AND symb_decoder(16#20#));
reg_q1341_init <= '0' ;
	p_reg_q1341: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1341 <= reg_q1341_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1341 <= reg_q1341_init;
        else
          reg_q1341 <= reg_q1341_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2215_in <= (reg_q2213 AND symb_decoder(16#69#)) OR
 					(reg_q2213 AND symb_decoder(16#49#));
reg_q2215_init <= '0' ;
	p_reg_q2215: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2215 <= reg_q2215_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2215 <= reg_q2215_init;
        else
          reg_q2215 <= reg_q2215_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q622_in <= (reg_q620 AND symb_decoder(16#45#)) OR
 					(reg_q620 AND symb_decoder(16#65#));
reg_q622_init <= '0' ;
	p_reg_q622: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q622 <= reg_q622_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q622 <= reg_q622_init;
        else
          reg_q622 <= reg_q622_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q624_in <= (reg_q622 AND symb_decoder(16#52#)) OR
 					(reg_q622 AND symb_decoder(16#72#));
reg_q624_init <= '0' ;
	p_reg_q624: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q624 <= reg_q624_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q624 <= reg_q624_init;
        else
          reg_q624 <= reg_q624_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1840_in <= (reg_q1838 AND symb_decoder(16#44#)) OR
 					(reg_q1838 AND symb_decoder(16#64#));
reg_q1840_init <= '0' ;
	p_reg_q1840: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1840 <= reg_q1840_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1840 <= reg_q1840_init;
        else
          reg_q1840 <= reg_q1840_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1842_in <= (reg_q1840 AND symb_decoder(16#6c#)) OR
 					(reg_q1840 AND symb_decoder(16#4c#));
reg_q1842_init <= '0' ;
	p_reg_q1842: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1842 <= reg_q1842_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1842 <= reg_q1842_init;
        else
          reg_q1842 <= reg_q1842_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q86_in <= (reg_q86 AND symb_decoder(16#20#)) OR
 					(reg_q86 AND symb_decoder(16#0d#)) OR
 					(reg_q86 AND symb_decoder(16#09#)) OR
 					(reg_q86 AND symb_decoder(16#0a#)) OR
 					(reg_q86 AND symb_decoder(16#0c#)) OR
 					(reg_q84 AND symb_decoder(16#0c#)) OR
 					(reg_q84 AND symb_decoder(16#09#)) OR
 					(reg_q84 AND symb_decoder(16#0d#)) OR
 					(reg_q84 AND symb_decoder(16#0a#)) OR
 					(reg_q84 AND symb_decoder(16#20#));
reg_q86_init <= '0' ;
	p_reg_q86: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q86 <= reg_q86_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q86 <= reg_q86_init;
        else
          reg_q86 <= reg_q86_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1522_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1521 AND symb_decoder(16#0d#)) OR
 					(reg_q1521 AND symb_decoder(16#0a#));
reg_q1522_init <= '0' ;
	p_reg_q1522: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1522 <= reg_q1522_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1522 <= reg_q1522_init;
        else
          reg_q1522 <= reg_q1522_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1523_in <= (reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q1522 AND symb_decoder(16#6e#)) OR
 					(reg_q1522 AND symb_decoder(16#4e#));
reg_q1523_init <= '0' ;
	p_reg_q1523: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1523 <= reg_q1523_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1523 <= reg_q1523_init;
        else
          reg_q1523 <= reg_q1523_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1403_in <= (reg_q1401 AND symb_decoder(16#65#)) OR
 					(reg_q1401 AND symb_decoder(16#45#));
reg_q1403_init <= '0' ;
	p_reg_q1403: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1403 <= reg_q1403_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1403 <= reg_q1403_init;
        else
          reg_q1403 <= reg_q1403_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1405_in <= (reg_q1403 AND symb_decoder(16#52#)) OR
 					(reg_q1403 AND symb_decoder(16#72#));
reg_q1405_init <= '0' ;
	p_reg_q1405: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1405 <= reg_q1405_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1405 <= reg_q1405_init;
        else
          reg_q1405 <= reg_q1405_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2054_in <= (reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2052 AND symb_decoder(16#54#));
reg_q2054_init <= '0' ;
	p_reg_q2054: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2054 <= reg_q2054_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2054 <= reg_q2054_init;
        else
          reg_q2054 <= reg_q2054_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1541_in <= (reg_q1541 AND symb_decoder(16#32#)) OR
 					(reg_q1541 AND symb_decoder(16#38#)) OR
 					(reg_q1541 AND symb_decoder(16#37#)) OR
 					(reg_q1541 AND symb_decoder(16#30#)) OR
 					(reg_q1541 AND symb_decoder(16#33#)) OR
 					(reg_q1541 AND symb_decoder(16#39#)) OR
 					(reg_q1541 AND symb_decoder(16#36#)) OR
 					(reg_q1541 AND symb_decoder(16#34#)) OR
 					(reg_q1541 AND symb_decoder(16#35#)) OR
 					(reg_q1541 AND symb_decoder(16#31#)) OR
 					(reg_q1539 AND symb_decoder(16#38#)) OR
 					(reg_q1539 AND symb_decoder(16#35#)) OR
 					(reg_q1539 AND symb_decoder(16#37#)) OR
 					(reg_q1539 AND symb_decoder(16#33#)) OR
 					(reg_q1539 AND symb_decoder(16#39#)) OR
 					(reg_q1539 AND symb_decoder(16#34#)) OR
 					(reg_q1539 AND symb_decoder(16#31#)) OR
 					(reg_q1539 AND symb_decoder(16#30#)) OR
 					(reg_q1539 AND symb_decoder(16#32#)) OR
 					(reg_q1539 AND symb_decoder(16#36#));
reg_q1541_init <= '0' ;
	p_reg_q1541: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1541 <= reg_q1541_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1541 <= reg_q1541_init;
        else
          reg_q1541 <= reg_q1541_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2684_in <= (reg_q2682 AND symb_decoder(16#74#)) OR
 					(reg_q2682 AND symb_decoder(16#54#));
reg_q2684_init <= '0' ;
	p_reg_q2684: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2684 <= reg_q2684_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2684 <= reg_q2684_init;
        else
          reg_q2684 <= reg_q2684_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2686_in <= (reg_q2684 AND symb_decoder(16#45#)) OR
 					(reg_q2684 AND symb_decoder(16#65#));
reg_q2686_init <= '0' ;
	p_reg_q2686: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2686 <= reg_q2686_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2686 <= reg_q2686_init;
        else
          reg_q2686 <= reg_q2686_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1784_in <= (reg_q1782 AND symb_decoder(16#09#)) OR
 					(reg_q1782 AND symb_decoder(16#0a#)) OR
 					(reg_q1782 AND symb_decoder(16#0d#)) OR
 					(reg_q1782 AND symb_decoder(16#0c#)) OR
 					(reg_q1782 AND symb_decoder(16#20#));
reg_q1784_init <= '0' ;
	p_reg_q1784: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1784 <= reg_q1784_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1784 <= reg_q1784_init;
        else
          reg_q1784 <= reg_q1784_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1786_in <= (reg_q1784 AND symb_decoder(16#0d#)) OR
 					(reg_q1784 AND symb_decoder(16#0c#)) OR
 					(reg_q1784 AND symb_decoder(16#09#)) OR
 					(reg_q1784 AND symb_decoder(16#0a#)) OR
 					(reg_q1784 AND symb_decoder(16#20#));
reg_q1786_init <= '0' ;
	p_reg_q1786: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1786 <= reg_q1786_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1786 <= reg_q1786_init;
        else
          reg_q1786 <= reg_q1786_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2499_in <= (reg_q2499 AND symb_decoder(16#37#)) OR
 					(reg_q2499 AND symb_decoder(16#39#)) OR
 					(reg_q2499 AND symb_decoder(16#34#)) OR
 					(reg_q2499 AND symb_decoder(16#36#)) OR
 					(reg_q2499 AND symb_decoder(16#32#)) OR
 					(reg_q2499 AND symb_decoder(16#38#)) OR
 					(reg_q2499 AND symb_decoder(16#30#)) OR
 					(reg_q2499 AND symb_decoder(16#35#)) OR
 					(reg_q2499 AND symb_decoder(16#31#)) OR
 					(reg_q2499 AND symb_decoder(16#33#)) OR
 					(reg_q2497 AND symb_decoder(16#39#)) OR
 					(reg_q2497 AND symb_decoder(16#34#)) OR
 					(reg_q2497 AND symb_decoder(16#33#)) OR
 					(reg_q2497 AND symb_decoder(16#38#)) OR
 					(reg_q2497 AND symb_decoder(16#32#)) OR
 					(reg_q2497 AND symb_decoder(16#37#)) OR
 					(reg_q2497 AND symb_decoder(16#31#)) OR
 					(reg_q2497 AND symb_decoder(16#30#)) OR
 					(reg_q2497 AND symb_decoder(16#36#)) OR
 					(reg_q2497 AND symb_decoder(16#35#));
reg_q2499_init <= '0' ;
	p_reg_q2499: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2499 <= reg_q2499_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2499 <= reg_q2499_init;
        else
          reg_q2499 <= reg_q2499_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1906_in <= (reg_q1904 AND symb_decoder(16#52#)) OR
 					(reg_q1904 AND symb_decoder(16#72#));
reg_q1906_init <= '0' ;
	p_reg_q1906: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1906 <= reg_q1906_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1906 <= reg_q1906_init;
        else
          reg_q1906 <= reg_q1906_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1908_in <= (reg_q1906 AND symb_decoder(16#65#)) OR
 					(reg_q1906 AND symb_decoder(16#45#));
reg_q1908_init <= '0' ;
	p_reg_q1908: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1908 <= reg_q1908_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1908 <= reg_q1908_init;
        else
          reg_q1908 <= reg_q1908_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q744_in <= (reg_q742 AND symb_decoder(16#65#)) OR
 					(reg_q742 AND symb_decoder(16#45#));
reg_q744_init <= '0' ;
	p_reg_q744: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q744 <= reg_q744_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q744 <= reg_q744_init;
        else
          reg_q744 <= reg_q744_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q746_in <= (reg_q744 AND symb_decoder(16#4e#)) OR
 					(reg_q744 AND symb_decoder(16#6e#));
reg_q746_init <= '0' ;
	p_reg_q746: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q746 <= reg_q746_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q746 <= reg_q746_init;
        else
          reg_q746 <= reg_q746_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1131_in <= (reg_q1129 AND symb_decoder(16#74#)) OR
 					(reg_q1129 AND symb_decoder(16#54#));
reg_q1131_init <= '0' ;
	p_reg_q1131: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1131 <= reg_q1131_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1131 <= reg_q1131_init;
        else
          reg_q1131 <= reg_q1131_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1133_in <= (reg_q1131 AND symb_decoder(16#52#)) OR
 					(reg_q1131 AND symb_decoder(16#72#));
reg_q1133_init <= '0' ;
	p_reg_q1133: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1133 <= reg_q1133_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1133 <= reg_q1133_init;
        else
          reg_q1133 <= reg_q1133_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1454_in <= (reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q1453 AND symb_decoder(16#68#)) OR
 					(reg_q1453 AND symb_decoder(16#48#));
reg_q1454_init <= '0' ;
	p_reg_q1454: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1454 <= reg_q1454_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1454 <= reg_q1454_init;
        else
          reg_q1454 <= reg_q1454_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1000_in <= (reg_q998 AND symb_decoder(16#70#)) OR
 					(reg_q998 AND symb_decoder(16#50#));
reg_q1000_init <= '0' ;
	p_reg_q1000: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1000 <= reg_q1000_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1000 <= reg_q1000_init;
        else
          reg_q1000 <= reg_q1000_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1002_in <= (reg_q1000 AND symb_decoder(16#0a#)) OR
 					(reg_q1000 AND symb_decoder(16#09#)) OR
 					(reg_q1000 AND symb_decoder(16#0d#)) OR
 					(reg_q1000 AND symb_decoder(16#0c#)) OR
 					(reg_q1000 AND symb_decoder(16#20#)) OR
 					(reg_q1002 AND symb_decoder(16#20#)) OR
 					(reg_q1002 AND symb_decoder(16#0a#)) OR
 					(reg_q1002 AND symb_decoder(16#09#)) OR
 					(reg_q1002 AND symb_decoder(16#0d#)) OR
 					(reg_q1002 AND symb_decoder(16#0c#));
reg_q1002_init <= '0' ;
	p_reg_q1002: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1002 <= reg_q1002_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1002 <= reg_q1002_init;
        else
          reg_q1002 <= reg_q1002_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1918_in <= (reg_q1918 AND symb_decoder(16#20#)) OR
 					(reg_q1918 AND symb_decoder(16#09#)) OR
 					(reg_q1918 AND symb_decoder(16#0c#)) OR
 					(reg_q1918 AND symb_decoder(16#0a#)) OR
 					(reg_q1918 AND symb_decoder(16#0d#)) OR
 					(reg_q1916 AND symb_decoder(16#0a#)) OR
 					(reg_q1916 AND symb_decoder(16#20#)) OR
 					(reg_q1916 AND symb_decoder(16#09#)) OR
 					(reg_q1916 AND symb_decoder(16#0d#)) OR
 					(reg_q1916 AND symb_decoder(16#0c#));
reg_q1918_init <= '0' ;
	p_reg_q1918: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1918 <= reg_q1918_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1918 <= reg_q1918_init;
        else
          reg_q1918 <= reg_q1918_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2280_in <= (reg_q2278 AND symb_decoder(16#76#)) OR
 					(reg_q2278 AND symb_decoder(16#56#));
reg_q2280_init <= '0' ;
	p_reg_q2280: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2280 <= reg_q2280_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2280 <= reg_q2280_init;
        else
          reg_q2280 <= reg_q2280_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2282_in <= (reg_q2280 AND symb_decoder(16#36#)) OR
 					(reg_q2280 AND symb_decoder(16#34#)) OR
 					(reg_q2280 AND symb_decoder(16#39#)) OR
 					(reg_q2280 AND symb_decoder(16#35#)) OR
 					(reg_q2280 AND symb_decoder(16#32#)) OR
 					(reg_q2280 AND symb_decoder(16#37#)) OR
 					(reg_q2280 AND symb_decoder(16#31#)) OR
 					(reg_q2280 AND symb_decoder(16#38#)) OR
 					(reg_q2280 AND symb_decoder(16#30#)) OR
 					(reg_q2280 AND symb_decoder(16#33#)) OR
 					(reg_q2282 AND symb_decoder(16#36#)) OR
 					(reg_q2282 AND symb_decoder(16#35#)) OR
 					(reg_q2282 AND symb_decoder(16#31#)) OR
 					(reg_q2282 AND symb_decoder(16#33#)) OR
 					(reg_q2282 AND symb_decoder(16#34#)) OR
 					(reg_q2282 AND symb_decoder(16#32#)) OR
 					(reg_q2282 AND symb_decoder(16#37#)) OR
 					(reg_q2282 AND symb_decoder(16#38#)) OR
 					(reg_q2282 AND symb_decoder(16#39#)) OR
 					(reg_q2282 AND symb_decoder(16#30#));
reg_q2282_init <= '0' ;
	p_reg_q2282: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2282 <= reg_q2282_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2282 <= reg_q2282_init;
        else
          reg_q2282 <= reg_q2282_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q239_in <= (reg_q237 AND symb_decoder(16#ff#));
reg_q239_init <= '0' ;
	p_reg_q239: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q239 <= reg_q239_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q239 <= reg_q239_init;
        else
          reg_q239 <= reg_q239_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2620_in <= (reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2619 AND symb_decoder(16#c0#));
reg_q2620_init <= '0' ;
	p_reg_q2620: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2620 <= reg_q2620_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2620 <= reg_q2620_init;
        else
          reg_q2620 <= reg_q2620_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2622_in <= (reg_q2620 AND symb_decoder(16#73#)) OR
 					(reg_q2620 AND symb_decoder(16#53#));
reg_q2622_init <= '0' ;
	p_reg_q2622: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2622 <= reg_q2622_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2622 <= reg_q2622_init;
        else
          reg_q2622 <= reg_q2622_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2569_in <= (reg_q2567 AND symb_decoder(16#57#)) OR
 					(reg_q2567 AND symb_decoder(16#77#));
reg_q2569_init <= '0' ;
	p_reg_q2569: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2569 <= reg_q2569_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2569 <= reg_q2569_init;
        else
          reg_q2569 <= reg_q2569_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2571_in <= (reg_q2569 AND symb_decoder(16#4e#)) OR
 					(reg_q2569 AND symb_decoder(16#6e#));
reg_q2571_init <= '0' ;
	p_reg_q2571: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2571 <= reg_q2571_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2571 <= reg_q2571_init;
        else
          reg_q2571 <= reg_q2571_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2072_in <= (reg_q2070 AND symb_decoder(16#50#));
reg_q2072_init <= '0' ;
	p_reg_q2072: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2072 <= reg_q2072_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2072 <= reg_q2072_init;
        else
          reg_q2072 <= reg_q2072_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2074_in <= (reg_q2072 AND symb_decoder(16#0c#)) OR
 					(reg_q2072 AND symb_decoder(16#0a#)) OR
 					(reg_q2072 AND symb_decoder(16#0d#)) OR
 					(reg_q2072 AND symb_decoder(16#20#)) OR
 					(reg_q2072 AND symb_decoder(16#09#)) OR
 					(reg_q2074 AND symb_decoder(16#0a#)) OR
 					(reg_q2074 AND symb_decoder(16#09#)) OR
 					(reg_q2074 AND symb_decoder(16#0d#)) OR
 					(reg_q2074 AND symb_decoder(16#20#)) OR
 					(reg_q2074 AND symb_decoder(16#0c#));
reg_q2074_init <= '0' ;
	p_reg_q2074: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2074 <= reg_q2074_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2074 <= reg_q2074_init;
        else
          reg_q2074 <= reg_q2074_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1060_in <= (reg_q1058 AND symb_decoder(16#4f#)) OR
 					(reg_q1058 AND symb_decoder(16#6f#));
reg_q1060_init <= '0' ;
	p_reg_q1060: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1060 <= reg_q1060_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1060 <= reg_q1060_init;
        else
          reg_q1060 <= reg_q1060_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1062_in <= (reg_q1060 AND symb_decoder(16#49#)) OR
 					(reg_q1060 AND symb_decoder(16#69#));
reg_q1062_init <= '0' ;
	p_reg_q1062: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1062 <= reg_q1062_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1062 <= reg_q1062_init;
        else
          reg_q1062 <= reg_q1062_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q133_in <= (reg_q131 AND symb_decoder(16#6f#)) OR
 					(reg_q131 AND symb_decoder(16#4f#));
reg_q133_init <= '0' ;
	p_reg_q133: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q133 <= reg_q133_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q133 <= reg_q133_init;
        else
          reg_q133 <= reg_q133_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q135_in <= (reg_q133 AND symb_decoder(16#6e#)) OR
 					(reg_q133 AND symb_decoder(16#4e#));
reg_q135_init <= '0' ;
	p_reg_q135: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q135 <= reg_q135_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q135 <= reg_q135_init;
        else
          reg_q135 <= reg_q135_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q341_in <= (reg_q339 AND symb_decoder(16#74#)) OR
 					(reg_q339 AND symb_decoder(16#54#));
reg_q341_init <= '0' ;
	p_reg_q341: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q341 <= reg_q341_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q341 <= reg_q341_init;
        else
          reg_q341 <= reg_q341_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q343_in <= (reg_q341 AND symb_decoder(16#72#)) OR
 					(reg_q341 AND symb_decoder(16#52#));
reg_q343_init <= '0' ;
	p_reg_q343: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q343 <= reg_q343_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q343 <= reg_q343_init;
        else
          reg_q343 <= reg_q343_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q797_in <= (reg_q797 AND symb_decoder(16#32#)) OR
 					(reg_q797 AND symb_decoder(16#30#)) OR
 					(reg_q797 AND symb_decoder(16#39#)) OR
 					(reg_q797 AND symb_decoder(16#36#)) OR
 					(reg_q797 AND symb_decoder(16#33#)) OR
 					(reg_q797 AND symb_decoder(16#35#)) OR
 					(reg_q797 AND symb_decoder(16#37#)) OR
 					(reg_q797 AND symb_decoder(16#38#)) OR
 					(reg_q797 AND symb_decoder(16#31#)) OR
 					(reg_q797 AND symb_decoder(16#34#)) OR
 					(reg_q795 AND symb_decoder(16#35#)) OR
 					(reg_q795 AND symb_decoder(16#34#)) OR
 					(reg_q795 AND symb_decoder(16#39#)) OR
 					(reg_q795 AND symb_decoder(16#30#)) OR
 					(reg_q795 AND symb_decoder(16#36#)) OR
 					(reg_q795 AND symb_decoder(16#31#)) OR
 					(reg_q795 AND symb_decoder(16#38#)) OR
 					(reg_q795 AND symb_decoder(16#37#)) OR
 					(reg_q795 AND symb_decoder(16#33#)) OR
 					(reg_q795 AND symb_decoder(16#32#));
reg_q797_init <= '0' ;
	p_reg_q797: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q797 <= reg_q797_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q797 <= reg_q797_init;
        else
          reg_q797 <= reg_q797_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1301_in <= (reg_q1299 AND symb_decoder(16#69#)) OR
 					(reg_q1299 AND symb_decoder(16#49#));
reg_q1301_init <= '0' ;
	p_reg_q1301: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1301 <= reg_q1301_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1301 <= reg_q1301_init;
        else
          reg_q1301 <= reg_q1301_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1303_in <= (reg_q1301 AND symb_decoder(16#72#)) OR
 					(reg_q1301 AND symb_decoder(16#52#));
reg_q1303_init <= '0' ;
	p_reg_q1303: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1303 <= reg_q1303_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1303 <= reg_q1303_init;
        else
          reg_q1303 <= reg_q1303_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q80_in <= (reg_q78 AND symb_decoder(16#76#)) OR
 					(reg_q78 AND symb_decoder(16#56#));
reg_q80_init <= '0' ;
	p_reg_q80: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q80 <= reg_q80_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q80 <= reg_q80_init;
        else
          reg_q80 <= reg_q80_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q82_in <= (reg_q80 AND symb_decoder(16#65#)) OR
 					(reg_q80 AND symb_decoder(16#45#));
reg_q82_init <= '0' ;
	p_reg_q82: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q82 <= reg_q82_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q82 <= reg_q82_init;
        else
          reg_q82 <= reg_q82_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q233_in <= (reg_q233 AND symb_decoder(16#33#)) OR
 					(reg_q233 AND symb_decoder(16#39#)) OR
 					(reg_q233 AND symb_decoder(16#35#)) OR
 					(reg_q233 AND symb_decoder(16#38#)) OR
 					(reg_q233 AND symb_decoder(16#32#)) OR
 					(reg_q233 AND symb_decoder(16#34#)) OR
 					(reg_q233 AND symb_decoder(16#36#)) OR
 					(reg_q233 AND symb_decoder(16#31#)) OR
 					(reg_q233 AND symb_decoder(16#30#)) OR
 					(reg_q233 AND symb_decoder(16#37#)) OR
 					(reg_q231 AND symb_decoder(16#34#)) OR
 					(reg_q231 AND symb_decoder(16#31#)) OR
 					(reg_q231 AND symb_decoder(16#36#)) OR
 					(reg_q231 AND symb_decoder(16#39#)) OR
 					(reg_q231 AND symb_decoder(16#32#)) OR
 					(reg_q231 AND symb_decoder(16#30#)) OR
 					(reg_q231 AND symb_decoder(16#33#)) OR
 					(reg_q231 AND symb_decoder(16#38#)) OR
 					(reg_q231 AND symb_decoder(16#37#)) OR
 					(reg_q231 AND symb_decoder(16#35#));
reg_q233_init <= '0' ;
	p_reg_q233: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q233 <= reg_q233_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q233 <= reg_q233_init;
        else
          reg_q233 <= reg_q233_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q840_in <= (reg_q840 AND symb_decoder(16#34#)) OR
 					(reg_q840 AND symb_decoder(16#35#)) OR
 					(reg_q840 AND symb_decoder(16#30#)) OR
 					(reg_q840 AND symb_decoder(16#36#)) OR
 					(reg_q840 AND symb_decoder(16#39#)) OR
 					(reg_q840 AND symb_decoder(16#37#)) OR
 					(reg_q840 AND symb_decoder(16#38#)) OR
 					(reg_q840 AND symb_decoder(16#31#)) OR
 					(reg_q840 AND symb_decoder(16#32#)) OR
 					(reg_q840 AND symb_decoder(16#33#)) OR
 					(reg_q838 AND symb_decoder(16#31#)) OR
 					(reg_q838 AND symb_decoder(16#35#)) OR
 					(reg_q838 AND symb_decoder(16#37#)) OR
 					(reg_q838 AND symb_decoder(16#32#)) OR
 					(reg_q838 AND symb_decoder(16#30#)) OR
 					(reg_q838 AND symb_decoder(16#39#)) OR
 					(reg_q838 AND symb_decoder(16#38#)) OR
 					(reg_q838 AND symb_decoder(16#33#)) OR
 					(reg_q838 AND symb_decoder(16#36#)) OR
 					(reg_q838 AND symb_decoder(16#34#));
reg_q840_init <= '0' ;
	p_reg_q840: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q840 <= reg_q840_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q840 <= reg_q840_init;
        else
          reg_q840 <= reg_q840_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q14_in <= (reg_q12 AND symb_decoder(16#65#)) OR
 					(reg_q12 AND symb_decoder(16#45#));
reg_q14_init <= '0' ;
	p_reg_q14: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q14 <= reg_q14_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q14 <= reg_q14_init;
        else
          reg_q14 <= reg_q14_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q16_in <= (reg_q14 AND symb_decoder(16#09#)) OR
 					(reg_q14 AND symb_decoder(16#0d#)) OR
 					(reg_q14 AND symb_decoder(16#20#)) OR
 					(reg_q14 AND symb_decoder(16#0a#)) OR
 					(reg_q14 AND symb_decoder(16#0c#)) OR
 					(reg_q16 AND symb_decoder(16#0c#)) OR
 					(reg_q16 AND symb_decoder(16#0a#)) OR
 					(reg_q16 AND symb_decoder(16#20#)) OR
 					(reg_q16 AND symb_decoder(16#0d#)) OR
 					(reg_q16 AND symb_decoder(16#09#));
reg_q16_init <= '0' ;
	p_reg_q16: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q16 <= reg_q16_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q16 <= reg_q16_init;
        else
          reg_q16 <= reg_q16_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1333_in <= (reg_q1333 AND symb_decoder(16#09#)) OR
 					(reg_q1333 AND symb_decoder(16#0d#)) OR
 					(reg_q1333 AND symb_decoder(16#20#)) OR
 					(reg_q1333 AND symb_decoder(16#0a#)) OR
 					(reg_q1333 AND symb_decoder(16#0c#)) OR
 					(reg_q1331 AND symb_decoder(16#09#)) OR
 					(reg_q1331 AND symb_decoder(16#0d#)) OR
 					(reg_q1331 AND symb_decoder(16#0a#)) OR
 					(reg_q1331 AND symb_decoder(16#0c#)) OR
 					(reg_q1331 AND symb_decoder(16#20#));
reg_q1333_init <= '0' ;
	p_reg_q1333: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1333 <= reg_q1333_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1333 <= reg_q1333_init;
        else
          reg_q1333 <= reg_q1333_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2367_in <= (reg_q2365 AND symb_decoder(16#22#));
reg_q2367_init <= '0' ;
	p_reg_q2367: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2367 <= reg_q2367_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2367 <= reg_q2367_init;
        else
          reg_q2367 <= reg_q2367_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2369_in <= (reg_q2367 AND symb_decoder(16#0a#)) OR
 					(reg_q2367 AND symb_decoder(16#20#)) OR
 					(reg_q2367 AND symb_decoder(16#0d#)) OR
 					(reg_q2367 AND symb_decoder(16#09#)) OR
 					(reg_q2367 AND symb_decoder(16#0c#)) OR
 					(reg_q2369 AND symb_decoder(16#0c#)) OR
 					(reg_q2369 AND symb_decoder(16#09#)) OR
 					(reg_q2369 AND symb_decoder(16#0d#)) OR
 					(reg_q2369 AND symb_decoder(16#20#)) OR
 					(reg_q2369 AND symb_decoder(16#0a#));
reg_q2369_init <= '0' ;
	p_reg_q2369: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2369 <= reg_q2369_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2369 <= reg_q2369_init;
        else
          reg_q2369 <= reg_q2369_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1068_in <= (reg_q1066 AND symb_decoder(16#52#)) OR
 					(reg_q1066 AND symb_decoder(16#72#));
reg_q1068_init <= '0' ;
	p_reg_q1068: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1068 <= reg_q1068_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1068 <= reg_q1068_init;
        else
          reg_q1068 <= reg_q1068_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1070_in <= (reg_q1068 AND symb_decoder(16#09#)) OR
 					(reg_q1068 AND symb_decoder(16#20#)) OR
 					(reg_q1068 AND symb_decoder(16#0a#)) OR
 					(reg_q1068 AND symb_decoder(16#0c#)) OR
 					(reg_q1068 AND symb_decoder(16#0d#)) OR
 					(reg_q1070 AND symb_decoder(16#0c#)) OR
 					(reg_q1070 AND symb_decoder(16#0d#)) OR
 					(reg_q1070 AND symb_decoder(16#20#)) OR
 					(reg_q1070 AND symb_decoder(16#0a#)) OR
 					(reg_q1070 AND symb_decoder(16#09#));
reg_q1070_init <= '0' ;
	p_reg_q1070: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1070 <= reg_q1070_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1070 <= reg_q1070_init;
        else
          reg_q1070 <= reg_q1070_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q732_in <= (reg_q730 AND symb_decoder(16#67#)) OR
 					(reg_q730 AND symb_decoder(16#47#));
reg_q732_init <= '0' ;
	p_reg_q732: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q732 <= reg_q732_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q732 <= reg_q732_init;
        else
          reg_q732 <= reg_q732_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q734_in <= (reg_q732 AND symb_decoder(16#09#)) OR
 					(reg_q732 AND symb_decoder(16#20#)) OR
 					(reg_q732 AND symb_decoder(16#0c#)) OR
 					(reg_q732 AND symb_decoder(16#0a#)) OR
 					(reg_q732 AND symb_decoder(16#0d#)) OR
 					(reg_q734 AND symb_decoder(16#20#)) OR
 					(reg_q734 AND symb_decoder(16#0a#)) OR
 					(reg_q734 AND symb_decoder(16#0d#)) OR
 					(reg_q734 AND symb_decoder(16#09#)) OR
 					(reg_q734 AND symb_decoder(16#0c#));
reg_q734_init <= '0' ;
	p_reg_q734: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q734 <= reg_q734_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q734 <= reg_q734_init;
        else
          reg_q734 <= reg_q734_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1762_in <= (reg_q1760 AND symb_decoder(16#0a#)) OR
 					(reg_q1760 AND symb_decoder(16#20#)) OR
 					(reg_q1760 AND symb_decoder(16#09#)) OR
 					(reg_q1760 AND symb_decoder(16#0d#)) OR
 					(reg_q1760 AND symb_decoder(16#0c#));
reg_q1762_init <= '0' ;
	p_reg_q1762: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1762 <= reg_q1762_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1762 <= reg_q1762_init;
        else
          reg_q1762 <= reg_q1762_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1764_in <= (reg_q1762 AND symb_decoder(16#09#)) OR
 					(reg_q1762 AND symb_decoder(16#0a#)) OR
 					(reg_q1762 AND symb_decoder(16#0c#)) OR
 					(reg_q1762 AND symb_decoder(16#20#)) OR
 					(reg_q1762 AND symb_decoder(16#0d#));
reg_q1764_init <= '0' ;
	p_reg_q1764: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1764 <= reg_q1764_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1764 <= reg_q1764_init;
        else
          reg_q1764 <= reg_q1764_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1250_in <= (reg_q1248 AND symb_decoder(16#56#)) OR
 					(reg_q1248 AND symb_decoder(16#76#));
reg_q1250_init <= '0' ;
	p_reg_q1250: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1250 <= reg_q1250_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1250 <= reg_q1250_init;
        else
          reg_q1250 <= reg_q1250_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1252_in <= (reg_q1250 AND symb_decoder(16#33#)) OR
 					(reg_q1250 AND symb_decoder(16#37#)) OR
 					(reg_q1250 AND symb_decoder(16#36#)) OR
 					(reg_q1250 AND symb_decoder(16#31#)) OR
 					(reg_q1250 AND symb_decoder(16#34#)) OR
 					(reg_q1250 AND symb_decoder(16#30#)) OR
 					(reg_q1250 AND symb_decoder(16#39#)) OR
 					(reg_q1250 AND symb_decoder(16#38#)) OR
 					(reg_q1250 AND symb_decoder(16#32#)) OR
 					(reg_q1250 AND symb_decoder(16#35#)) OR
 					(reg_q1252 AND symb_decoder(16#39#)) OR
 					(reg_q1252 AND symb_decoder(16#30#)) OR
 					(reg_q1252 AND symb_decoder(16#38#)) OR
 					(reg_q1252 AND symb_decoder(16#32#)) OR
 					(reg_q1252 AND symb_decoder(16#33#)) OR
 					(reg_q1252 AND symb_decoder(16#31#)) OR
 					(reg_q1252 AND symb_decoder(16#35#)) OR
 					(reg_q1252 AND symb_decoder(16#36#)) OR
 					(reg_q1252 AND symb_decoder(16#34#)) OR
 					(reg_q1252 AND symb_decoder(16#37#));
reg_q1252_init <= '0' ;
	p_reg_q1252: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1252 <= reg_q1252_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1252 <= reg_q1252_init;
        else
          reg_q1252 <= reg_q1252_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1666_in <= (reg_q1666 AND symb_decoder(16#39#)) OR
 					(reg_q1666 AND symb_decoder(16#33#)) OR
 					(reg_q1666 AND symb_decoder(16#35#)) OR
 					(reg_q1666 AND symb_decoder(16#37#)) OR
 					(reg_q1666 AND symb_decoder(16#38#)) OR
 					(reg_q1666 AND symb_decoder(16#32#)) OR
 					(reg_q1666 AND symb_decoder(16#34#)) OR
 					(reg_q1666 AND symb_decoder(16#30#)) OR
 					(reg_q1666 AND symb_decoder(16#31#)) OR
 					(reg_q1666 AND symb_decoder(16#36#)) OR
 					(reg_q1664 AND symb_decoder(16#30#)) OR
 					(reg_q1664 AND symb_decoder(16#38#)) OR
 					(reg_q1664 AND symb_decoder(16#37#)) OR
 					(reg_q1664 AND symb_decoder(16#35#)) OR
 					(reg_q1664 AND symb_decoder(16#33#)) OR
 					(reg_q1664 AND symb_decoder(16#31#)) OR
 					(reg_q1664 AND symb_decoder(16#34#)) OR
 					(reg_q1664 AND symb_decoder(16#39#)) OR
 					(reg_q1664 AND symb_decoder(16#36#)) OR
 					(reg_q1664 AND symb_decoder(16#32#));
reg_q1666_init <= '0' ;
	p_reg_q1666: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1666 <= reg_q1666_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1666 <= reg_q1666_init;
        else
          reg_q1666 <= reg_q1666_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1127_in <= (reg_q1125 AND symb_decoder(16#45#)) OR
 					(reg_q1125 AND symb_decoder(16#65#));
reg_q1127_init <= '0' ;
	p_reg_q1127: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1127 <= reg_q1127_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1127 <= reg_q1127_init;
        else
          reg_q1127 <= reg_q1127_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1129_in <= (reg_q1127 AND symb_decoder(16#6e#)) OR
 					(reg_q1127 AND symb_decoder(16#4e#));
reg_q1129_init <= '0' ;
	p_reg_q1129: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1129 <= reg_q1129_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1129 <= reg_q1129_init;
        else
          reg_q1129 <= reg_q1129_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q558_in <= (reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q556 AND symb_decoder(16#42#)) OR
 					(reg_q556 AND symb_decoder(16#62#));
reg_q558_init <= '0' ;
	p_reg_q558: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q558 <= reg_q558_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q558 <= reg_q558_init;
        else
          reg_q558 <= reg_q558_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q560_in <= (reg_q558 AND symb_decoder(16#4f#)) OR
 					(reg_q558 AND symb_decoder(16#6f#));
reg_q560_init <= '0' ;
	p_reg_q560: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q560 <= reg_q560_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q560 <= reg_q560_init;
        else
          reg_q560 <= reg_q560_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2415_in <= (reg_q2413 AND symb_decoder(16#69#)) OR
 					(reg_q2413 AND symb_decoder(16#49#));
reg_q2415_init <= '0' ;
	p_reg_q2415: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2415 <= reg_q2415_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2415 <= reg_q2415_init;
        else
          reg_q2415 <= reg_q2415_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2417_in <= (reg_q2415 AND symb_decoder(16#0d#)) OR
 					(reg_q2415 AND symb_decoder(16#09#)) OR
 					(reg_q2415 AND symb_decoder(16#0c#)) OR
 					(reg_q2415 AND symb_decoder(16#0a#)) OR
 					(reg_q2415 AND symb_decoder(16#20#)) OR
 					(reg_q2417 AND symb_decoder(16#0a#)) OR
 					(reg_q2417 AND symb_decoder(16#0c#)) OR
 					(reg_q2417 AND symb_decoder(16#20#)) OR
 					(reg_q2417 AND symb_decoder(16#0d#)) OR
 					(reg_q2417 AND symb_decoder(16#09#));
reg_q2417_init <= '0' ;
	p_reg_q2417: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2417 <= reg_q2417_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2417 <= reg_q2417_init;
        else
          reg_q2417 <= reg_q2417_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q781_in <= (reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q780 AND symb_decoder(16#64#)) OR
 					(reg_q780 AND symb_decoder(16#44#));
reg_q781_init <= '0' ;
	p_reg_q781: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q781 <= reg_q781_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q781 <= reg_q781_init;
        else
          reg_q781 <= reg_q781_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q397_in <= (reg_q397 AND symb_decoder(16#09#)) OR
 					(reg_q397 AND symb_decoder(16#20#)) OR
 					(reg_q397 AND symb_decoder(16#0d#)) OR
 					(reg_q397 AND symb_decoder(16#0c#)) OR
 					(reg_q397 AND symb_decoder(16#0a#)) OR
 					(reg_q395 AND symb_decoder(16#0c#)) OR
 					(reg_q395 AND symb_decoder(16#0a#)) OR
 					(reg_q395 AND symb_decoder(16#09#)) OR
 					(reg_q395 AND symb_decoder(16#20#)) OR
 					(reg_q395 AND symb_decoder(16#0d#));
reg_q397_init <= '0' ;
	p_reg_q397: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q397 <= reg_q397_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q397 <= reg_q397_init;
        else
          reg_q397 <= reg_q397_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q742_in <= (reg_q740 AND symb_decoder(16#54#)) OR
 					(reg_q740 AND symb_decoder(16#74#));
reg_q742_init <= '0' ;
	p_reg_q742: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q742 <= reg_q742_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q742 <= reg_q742_init;
        else
          reg_q742 <= reg_q742_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2241_in <= (reg_q2239 AND symb_decoder(16#72#)) OR
 					(reg_q2239 AND symb_decoder(16#52#));
reg_q2241_init <= '0' ;
	p_reg_q2241: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2241 <= reg_q2241_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2241 <= reg_q2241_init;
        else
          reg_q2241 <= reg_q2241_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2243_in <= (reg_q2241 AND symb_decoder(16#0a#)) OR
 					(reg_q2241 AND symb_decoder(16#0d#)) OR
 					(reg_q2241 AND symb_decoder(16#0c#)) OR
 					(reg_q2241 AND symb_decoder(16#20#)) OR
 					(reg_q2241 AND symb_decoder(16#09#)) OR
 					(reg_q2243 AND symb_decoder(16#20#)) OR
 					(reg_q2243 AND symb_decoder(16#09#)) OR
 					(reg_q2243 AND symb_decoder(16#0c#)) OR
 					(reg_q2243 AND symb_decoder(16#0d#)) OR
 					(reg_q2243 AND symb_decoder(16#0a#));
reg_q2243_init <= '0' ;
	p_reg_q2243: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2243 <= reg_q2243_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2243 <= reg_q2243_init;
        else
          reg_q2243 <= reg_q2243_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q251_in <= (reg_q249 AND symb_decoder(16#ff#));
reg_q251_init <= '0' ;
	p_reg_q251: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q251 <= reg_q251_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q251 <= reg_q251_init;
        else
          reg_q251 <= reg_q251_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q253_in <= (reg_q251 AND symb_decoder(16#38#)) OR
 					(reg_q251 AND symb_decoder(16#34#)) OR
 					(reg_q251 AND symb_decoder(16#36#)) OR
 					(reg_q251 AND symb_decoder(16#37#)) OR
 					(reg_q251 AND symb_decoder(16#33#)) OR
 					(reg_q251 AND symb_decoder(16#30#)) OR
 					(reg_q251 AND symb_decoder(16#39#)) OR
 					(reg_q251 AND symb_decoder(16#32#)) OR
 					(reg_q251 AND symb_decoder(16#31#)) OR
 					(reg_q251 AND symb_decoder(16#35#)) OR
 					(reg_q253 AND symb_decoder(16#30#)) OR
 					(reg_q253 AND symb_decoder(16#32#)) OR
 					(reg_q253 AND symb_decoder(16#38#)) OR
 					(reg_q253 AND symb_decoder(16#33#)) OR
 					(reg_q253 AND symb_decoder(16#35#)) OR
 					(reg_q253 AND symb_decoder(16#39#)) OR
 					(reg_q253 AND symb_decoder(16#31#)) OR
 					(reg_q253 AND symb_decoder(16#37#)) OR
 					(reg_q253 AND symb_decoder(16#36#)) OR
 					(reg_q253 AND symb_decoder(16#34#));
reg_q253_init <= '0' ;
	p_reg_q253: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q253 <= reg_q253_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q253 <= reg_q253_init;
        else
          reg_q253 <= reg_q253_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1712_in <= (reg_q1710 AND symb_decoder(16#4f#)) OR
 					(reg_q1710 AND symb_decoder(16#6f#));
reg_q1712_init <= '0' ;
	p_reg_q1712: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1712 <= reg_q1712_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1712 <= reg_q1712_init;
        else
          reg_q1712 <= reg_q1712_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1714_in <= (reg_q1712 AND symb_decoder(16#72#)) OR
 					(reg_q1712 AND symb_decoder(16#52#));
reg_q1714_init <= '0' ;
	p_reg_q1714: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1714 <= reg_q1714_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1714 <= reg_q1714_init;
        else
          reg_q1714 <= reg_q1714_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q371_in <= (reg_q371 AND symb_decoder(16#09#)) OR
 					(reg_q371 AND symb_decoder(16#0c#)) OR
 					(reg_q371 AND symb_decoder(16#0a#)) OR
 					(reg_q371 AND symb_decoder(16#20#)) OR
 					(reg_q371 AND symb_decoder(16#0d#)) OR
 					(reg_q369 AND symb_decoder(16#20#)) OR
 					(reg_q369 AND symb_decoder(16#09#)) OR
 					(reg_q369 AND symb_decoder(16#0c#)) OR
 					(reg_q369 AND symb_decoder(16#0a#)) OR
 					(reg_q369 AND symb_decoder(16#0d#));
reg_q371_init <= '0' ;
	p_reg_q371: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q371 <= reg_q371_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q371 <= reg_q371_init;
        else
          reg_q371 <= reg_q371_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1756_in <= (reg_q1754 AND symb_decoder(16#0a#)) OR
 					(reg_q1754 AND symb_decoder(16#0d#)) OR
 					(reg_q1754 AND symb_decoder(16#20#)) OR
 					(reg_q1754 AND symb_decoder(16#0c#)) OR
 					(reg_q1754 AND symb_decoder(16#09#));
reg_q1756_init <= '0' ;
	p_reg_q1756: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1756 <= reg_q1756_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1756 <= reg_q1756_init;
        else
          reg_q1756 <= reg_q1756_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1758_in <= (reg_q1756 AND symb_decoder(16#0c#)) OR
 					(reg_q1756 AND symb_decoder(16#0d#)) OR
 					(reg_q1756 AND symb_decoder(16#0a#)) OR
 					(reg_q1756 AND symb_decoder(16#09#)) OR
 					(reg_q1756 AND symb_decoder(16#20#));
reg_q1758_init <= '0' ;
	p_reg_q1758: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1758 <= reg_q1758_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1758 <= reg_q1758_init;
        else
          reg_q1758 <= reg_q1758_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2468_in <= (reg_q2695 AND symb_decoder(16#2a#));
reg_q2468_init <= '0' ;
	p_reg_q2468: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2468 <= reg_q2468_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2468 <= reg_q2468_init;
        else
          reg_q2468 <= reg_q2468_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2470_in <= (reg_q2468 AND symb_decoder(16#50#));
reg_q2470_init <= '0' ;
	p_reg_q2470: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2470 <= reg_q2470_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2470 <= reg_q2470_init;
        else
          reg_q2470 <= reg_q2470_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1696_in <= (reg_q1694 AND symb_decoder(16#75#)) OR
 					(reg_q1694 AND symb_decoder(16#55#));
reg_q1696_init <= '0' ;
	p_reg_q1696: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1696 <= reg_q1696_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1696 <= reg_q1696_init;
        else
          reg_q1696 <= reg_q1696_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1698_in <= (reg_q1696 AND symb_decoder(16#61#)) OR
 					(reg_q1696 AND symb_decoder(16#41#));
reg_q1698_init <= '0' ;
	p_reg_q1698: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1698 <= reg_q1698_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1698 <= reg_q1698_init;
        else
          reg_q1698 <= reg_q1698_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q704_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q703 AND symb_decoder(16#0d#)) OR
 					(reg_q703 AND symb_decoder(16#0a#));
reg_q704_init <= '0' ;
	p_reg_q704: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q704 <= reg_q704_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q704 <= reg_q704_init;
        else
          reg_q704 <= reg_q704_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q901_in <= (reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q901 AND symb_decoder(16#36#)) OR
 					(reg_q901 AND symb_decoder(16#33#)) OR
 					(reg_q901 AND symb_decoder(16#34#)) OR
 					(reg_q901 AND symb_decoder(16#31#)) OR
 					(reg_q901 AND symb_decoder(16#38#)) OR
 					(reg_q901 AND symb_decoder(16#35#)) OR
 					(reg_q901 AND symb_decoder(16#30#)) OR
 					(reg_q901 AND symb_decoder(16#37#)) OR
 					(reg_q901 AND symb_decoder(16#32#)) OR
 					(reg_q901 AND symb_decoder(16#39#)) OR
 					(reg_q900 AND symb_decoder(16#35#)) OR
 					(reg_q900 AND symb_decoder(16#34#)) OR
 					(reg_q900 AND symb_decoder(16#31#)) OR
 					(reg_q900 AND symb_decoder(16#37#)) OR
 					(reg_q900 AND symb_decoder(16#38#)) OR
 					(reg_q900 AND symb_decoder(16#36#)) OR
 					(reg_q900 AND symb_decoder(16#33#)) OR
 					(reg_q900 AND symb_decoder(16#32#)) OR
 					(reg_q900 AND symb_decoder(16#30#)) OR
 					(reg_q900 AND symb_decoder(16#39#));
reg_q901_init <= '0' ;
	p_reg_q901: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q901 <= reg_q901_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q901 <= reg_q901_init;
        else
          reg_q901 <= reg_q901_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2624_in <= (reg_q2622 AND symb_decoder(16#54#)) OR
 					(reg_q2622 AND symb_decoder(16#74#));
reg_q2624_init <= '0' ;
	p_reg_q2624: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2624 <= reg_q2624_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2624 <= reg_q2624_init;
        else
          reg_q2624 <= reg_q2624_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q962_in <= (reg_q960 AND symb_decoder(16#2d#));
reg_q962_init <= '0' ;
	p_reg_q962: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q962 <= reg_q962_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q962 <= reg_q962_init;
        else
          reg_q962 <= reg_q962_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q964_in <= (reg_q962 AND symb_decoder(16#09#)) OR
 					(reg_q962 AND symb_decoder(16#20#)) OR
 					(reg_q962 AND symb_decoder(16#0d#)) OR
 					(reg_q962 AND symb_decoder(16#0c#)) OR
 					(reg_q962 AND symb_decoder(16#0a#)) OR
 					(reg_q964 AND symb_decoder(16#0a#)) OR
 					(reg_q964 AND symb_decoder(16#0c#)) OR
 					(reg_q964 AND symb_decoder(16#0d#)) OR
 					(reg_q964 AND symb_decoder(16#20#)) OR
 					(reg_q964 AND symb_decoder(16#09#));
reg_q964_init <= '0' ;
	p_reg_q964: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q964 <= reg_q964_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q964 <= reg_q964_init;
        else
          reg_q964 <= reg_q964_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q424_in <= (reg_q422 AND symb_decoder(16#45#)) OR
 					(reg_q422 AND symb_decoder(16#65#));
reg_q424_init <= '0' ;
	p_reg_q424: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q424 <= reg_q424_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q424 <= reg_q424_init;
        else
          reg_q424 <= reg_q424_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1822_in <= (reg_q1820 AND symb_decoder(16#2e#));
reg_q1822_init <= '0' ;
	p_reg_q1822: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1822 <= reg_q1822_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1822 <= reg_q1822_init;
        else
          reg_q1822 <= reg_q1822_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1824_in <= (reg_q1822 AND symb_decoder(16#34#)) OR
 					(reg_q1822 AND symb_decoder(16#37#)) OR
 					(reg_q1822 AND symb_decoder(16#35#)) OR
 					(reg_q1822 AND symb_decoder(16#36#)) OR
 					(reg_q1822 AND symb_decoder(16#39#)) OR
 					(reg_q1822 AND symb_decoder(16#30#)) OR
 					(reg_q1822 AND symb_decoder(16#32#)) OR
 					(reg_q1822 AND symb_decoder(16#38#)) OR
 					(reg_q1822 AND symb_decoder(16#31#)) OR
 					(reg_q1822 AND symb_decoder(16#33#)) OR
 					(reg_q1824 AND symb_decoder(16#39#)) OR
 					(reg_q1824 AND symb_decoder(16#34#)) OR
 					(reg_q1824 AND symb_decoder(16#30#)) OR
 					(reg_q1824 AND symb_decoder(16#33#)) OR
 					(reg_q1824 AND symb_decoder(16#38#)) OR
 					(reg_q1824 AND symb_decoder(16#31#)) OR
 					(reg_q1824 AND symb_decoder(16#35#)) OR
 					(reg_q1824 AND symb_decoder(16#36#)) OR
 					(reg_q1824 AND symb_decoder(16#32#)) OR
 					(reg_q1824 AND symb_decoder(16#37#));
reg_q1824_init <= '0' ;
	p_reg_q1824: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1824 <= reg_q1824_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1824 <= reg_q1824_init;
        else
          reg_q1824 <= reg_q1824_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1317_in <= (reg_q1315 AND symb_decoder(16#44#)) OR
 					(reg_q1315 AND symb_decoder(16#64#));
reg_q1317_init <= '0' ;
	p_reg_q1317: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1317 <= reg_q1317_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1317 <= reg_q1317_init;
        else
          reg_q1317 <= reg_q1317_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1319_in <= (reg_q1317 AND symb_decoder(16#0a#)) OR
 					(reg_q1317 AND symb_decoder(16#0d#)) OR
 					(reg_q1317 AND symb_decoder(16#09#)) OR
 					(reg_q1317 AND symb_decoder(16#20#)) OR
 					(reg_q1317 AND symb_decoder(16#0c#)) OR
 					(reg_q1319 AND symb_decoder(16#0c#)) OR
 					(reg_q1319 AND symb_decoder(16#0a#)) OR
 					(reg_q1319 AND symb_decoder(16#20#)) OR
 					(reg_q1319 AND symb_decoder(16#09#)) OR
 					(reg_q1319 AND symb_decoder(16#0d#));
reg_q1319_init <= '0' ;
	p_reg_q1319: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1319 <= reg_q1319_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1319 <= reg_q1319_init;
        else
          reg_q1319 <= reg_q1319_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2577_in <= (reg_q2575 AND symb_decoder(16#3a#));
reg_q2577_init <= '0' ;
	p_reg_q2577: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2577 <= reg_q2577_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2577 <= reg_q2577_init;
        else
          reg_q2577 <= reg_q2577_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q620_in <= (reg_q618 AND symb_decoder(16#53#)) OR
 					(reg_q618 AND symb_decoder(16#73#));
reg_q620_init <= '0' ;
	p_reg_q620: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q620 <= reg_q620_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q620 <= reg_q620_init;
        else
          reg_q620 <= reg_q620_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q692_in <= (reg_q690 AND symb_decoder(16#36#)) OR
 					(reg_q690 AND symb_decoder(16#34#)) OR
 					(reg_q690 AND symb_decoder(16#32#)) OR
 					(reg_q690 AND symb_decoder(16#37#)) OR
 					(reg_q690 AND symb_decoder(16#38#)) OR
 					(reg_q690 AND symb_decoder(16#31#)) OR
 					(reg_q690 AND symb_decoder(16#33#)) OR
 					(reg_q690 AND symb_decoder(16#35#)) OR
 					(reg_q690 AND symb_decoder(16#30#)) OR
 					(reg_q690 AND symb_decoder(16#39#)) OR
 					(reg_q692 AND symb_decoder(16#38#)) OR
 					(reg_q692 AND symb_decoder(16#39#)) OR
 					(reg_q692 AND symb_decoder(16#37#)) OR
 					(reg_q692 AND symb_decoder(16#30#)) OR
 					(reg_q692 AND symb_decoder(16#31#)) OR
 					(reg_q692 AND symb_decoder(16#36#)) OR
 					(reg_q692 AND symb_decoder(16#32#)) OR
 					(reg_q692 AND symb_decoder(16#33#)) OR
 					(reg_q692 AND symb_decoder(16#34#)) OR
 					(reg_q692 AND symb_decoder(16#35#));
reg_q692_init <= '0' ;
	p_reg_q692: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q692 <= reg_q692_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q692 <= reg_q692_init;
        else
          reg_q692 <= reg_q692_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q367_in <= (reg_q365 AND symb_decoder(16#2e#));
reg_q367_init <= '0' ;
	p_reg_q367: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q367 <= reg_q367_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q367 <= reg_q367_init;
        else
          reg_q367 <= reg_q367_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q369_in <= (reg_q367 AND symb_decoder(16#37#)) OR
 					(reg_q367 AND symb_decoder(16#33#)) OR
 					(reg_q367 AND symb_decoder(16#32#)) OR
 					(reg_q367 AND symb_decoder(16#30#)) OR
 					(reg_q367 AND symb_decoder(16#31#)) OR
 					(reg_q367 AND symb_decoder(16#38#)) OR
 					(reg_q367 AND symb_decoder(16#35#)) OR
 					(reg_q367 AND symb_decoder(16#39#)) OR
 					(reg_q367 AND symb_decoder(16#36#)) OR
 					(reg_q367 AND symb_decoder(16#34#)) OR
 					(reg_q369 AND symb_decoder(16#39#)) OR
 					(reg_q369 AND symb_decoder(16#31#)) OR
 					(reg_q369 AND symb_decoder(16#38#)) OR
 					(reg_q369 AND symb_decoder(16#37#)) OR
 					(reg_q369 AND symb_decoder(16#30#)) OR
 					(reg_q369 AND symb_decoder(16#34#)) OR
 					(reg_q369 AND symb_decoder(16#35#)) OR
 					(reg_q369 AND symb_decoder(16#33#)) OR
 					(reg_q369 AND symb_decoder(16#32#)) OR
 					(reg_q369 AND symb_decoder(16#36#));
reg_q369_init <= '0' ;
	p_reg_q369: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q369 <= reg_q369_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q369 <= reg_q369_init;
        else
          reg_q369 <= reg_q369_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2535_in <= (reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2534 AND symb_decoder(16#2f#));
reg_q2535_init <= '0' ;
	p_reg_q2535: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2535 <= reg_q2535_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2535 <= reg_q2535_init;
        else
          reg_q2535 <= reg_q2535_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1221_in <= (reg_q1219 AND symb_decoder(16#0a#)) OR
 					(reg_q1219 AND symb_decoder(16#0c#)) OR
 					(reg_q1219 AND symb_decoder(16#09#)) OR
 					(reg_q1219 AND symb_decoder(16#0d#)) OR
 					(reg_q1219 AND symb_decoder(16#20#)) OR
 					(reg_q1221 AND symb_decoder(16#20#)) OR
 					(reg_q1221 AND symb_decoder(16#0d#)) OR
 					(reg_q1221 AND symb_decoder(16#09#)) OR
 					(reg_q1221 AND symb_decoder(16#0c#)) OR
 					(reg_q1221 AND symb_decoder(16#0a#));
reg_q1221_init <= '0' ;
	p_reg_q1221: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1221 <= reg_q1221_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1221 <= reg_q1221_init;
        else
          reg_q1221 <= reg_q1221_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1108_in <= (reg_q1106 AND symb_decoder(16#37#)) OR
 					(reg_q1106 AND symb_decoder(16#30#)) OR
 					(reg_q1106 AND symb_decoder(16#36#)) OR
 					(reg_q1106 AND symb_decoder(16#32#)) OR
 					(reg_q1106 AND symb_decoder(16#39#)) OR
 					(reg_q1106 AND symb_decoder(16#31#)) OR
 					(reg_q1106 AND symb_decoder(16#34#)) OR
 					(reg_q1106 AND symb_decoder(16#35#)) OR
 					(reg_q1106 AND symb_decoder(16#38#)) OR
 					(reg_q1106 AND symb_decoder(16#33#)) OR
 					(reg_q1108 AND symb_decoder(16#38#)) OR
 					(reg_q1108 AND symb_decoder(16#34#)) OR
 					(reg_q1108 AND symb_decoder(16#30#)) OR
 					(reg_q1108 AND symb_decoder(16#31#)) OR
 					(reg_q1108 AND symb_decoder(16#37#)) OR
 					(reg_q1108 AND symb_decoder(16#36#)) OR
 					(reg_q1108 AND symb_decoder(16#35#)) OR
 					(reg_q1108 AND symb_decoder(16#39#)) OR
 					(reg_q1108 AND symb_decoder(16#33#)) OR
 					(reg_q1108 AND symb_decoder(16#32#));
reg_q1108_init <= '0' ;
	p_reg_q1108: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1108 <= reg_q1108_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1108 <= reg_q1108_init;
        else
          reg_q1108 <= reg_q1108_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q686_in <= (reg_q684 AND symb_decoder(16#20#)) OR
 					(reg_q684 AND symb_decoder(16#0d#)) OR
 					(reg_q684 AND symb_decoder(16#09#)) OR
 					(reg_q684 AND symb_decoder(16#0c#)) OR
 					(reg_q684 AND symb_decoder(16#0a#));
reg_q686_init <= '0' ;
	p_reg_q686: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q686 <= reg_q686_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q686 <= reg_q686_init;
        else
          reg_q686 <= reg_q686_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1580_in <= (reg_q1580 AND symb_decoder(16#34#)) OR
 					(reg_q1580 AND symb_decoder(16#32#)) OR
 					(reg_q1580 AND symb_decoder(16#39#)) OR
 					(reg_q1580 AND symb_decoder(16#37#)) OR
 					(reg_q1580 AND symb_decoder(16#38#)) OR
 					(reg_q1580 AND symb_decoder(16#36#)) OR
 					(reg_q1580 AND symb_decoder(16#33#)) OR
 					(reg_q1580 AND symb_decoder(16#30#)) OR
 					(reg_q1580 AND symb_decoder(16#31#)) OR
 					(reg_q1580 AND symb_decoder(16#35#)) OR
 					(reg_q1578 AND symb_decoder(16#39#)) OR
 					(reg_q1578 AND symb_decoder(16#37#)) OR
 					(reg_q1578 AND symb_decoder(16#32#)) OR
 					(reg_q1578 AND symb_decoder(16#31#)) OR
 					(reg_q1578 AND symb_decoder(16#38#)) OR
 					(reg_q1578 AND symb_decoder(16#35#)) OR
 					(reg_q1578 AND symb_decoder(16#36#)) OR
 					(reg_q1578 AND symb_decoder(16#34#)) OR
 					(reg_q1578 AND symb_decoder(16#33#)) OR
 					(reg_q1578 AND symb_decoder(16#30#));
reg_q1580_init <= '0' ;
	p_reg_q1580: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1580 <= reg_q1580_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1580 <= reg_q1580_init;
        else
          reg_q1580 <= reg_q1580_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q866_in <= (reg_q864 AND symb_decoder(16#6c#)) OR
 					(reg_q864 AND symb_decoder(16#4c#));
reg_q866_init <= '0' ;
	p_reg_q866: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q866 <= reg_q866_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q866 <= reg_q866_init;
        else
          reg_q866 <= reg_q866_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q868_in <= (reg_q866 AND symb_decoder(16#49#)) OR
 					(reg_q866 AND symb_decoder(16#69#));
reg_q868_init <= '0' ;
	p_reg_q868: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q868 <= reg_q868_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q868 <= reg_q868_init;
        else
          reg_q868 <= reg_q868_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1371_in <= (reg_q1369 AND symb_decoder(16#45#)) OR
 					(reg_q1369 AND symb_decoder(16#65#));
reg_q1371_init <= '0' ;
	p_reg_q1371: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1371 <= reg_q1371_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1371 <= reg_q1371_init;
        else
          reg_q1371 <= reg_q1371_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1373_in <= (reg_q1371 AND symb_decoder(16#0a#)) OR
 					(reg_q1371 AND symb_decoder(16#0d#)) OR
 					(reg_q1371 AND symb_decoder(16#0c#)) OR
 					(reg_q1371 AND symb_decoder(16#09#)) OR
 					(reg_q1371 AND symb_decoder(16#20#)) OR
 					(reg_q1373 AND symb_decoder(16#20#)) OR
 					(reg_q1373 AND symb_decoder(16#0a#)) OR
 					(reg_q1373 AND symb_decoder(16#09#)) OR
 					(reg_q1373 AND symb_decoder(16#0d#)) OR
 					(reg_q1373 AND symb_decoder(16#0c#));
reg_q1373_init <= '0' ;
	p_reg_q1373: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1373 <= reg_q1373_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1373 <= reg_q1373_init;
        else
          reg_q1373 <= reg_q1373_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1558_in <= (reg_q1558 AND symb_decoder(16#09#)) OR
 					(reg_q1558 AND symb_decoder(16#20#)) OR
 					(reg_q1558 AND symb_decoder(16#0d#)) OR
 					(reg_q1558 AND symb_decoder(16#0a#)) OR
 					(reg_q1558 AND symb_decoder(16#0c#)) OR
 					(reg_q1556 AND symb_decoder(16#0d#)) OR
 					(reg_q1556 AND symb_decoder(16#0a#)) OR
 					(reg_q1556 AND symb_decoder(16#0c#)) OR
 					(reg_q1556 AND symb_decoder(16#09#)) OR
 					(reg_q1556 AND symb_decoder(16#20#));
reg_q1558_init <= '0' ;
	p_reg_q1558: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1558 <= reg_q1558_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1558 <= reg_q1558_init;
        else
          reg_q1558 <= reg_q1558_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1045_in <= (reg_q1043 AND symb_decoder(16#65#)) OR
 					(reg_q1043 AND symb_decoder(16#45#));
reg_q1045_init <= '0' ;
	p_reg_q1045: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1045 <= reg_q1045_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1045 <= reg_q1045_init;
        else
          reg_q1045 <= reg_q1045_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1047_in <= (reg_q1045 AND symb_decoder(16#72#)) OR
 					(reg_q1045 AND symb_decoder(16#52#));
reg_q1047_init <= '0' ;
	p_reg_q1047: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1047 <= reg_q1047_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1047 <= reg_q1047_init;
        else
          reg_q1047 <= reg_q1047_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2599_in <= (reg_q2597 AND symb_decoder(16#74#)) OR
 					(reg_q2597 AND symb_decoder(16#54#));
reg_q2599_init <= '0' ;
	p_reg_q2599: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2599 <= reg_q2599_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2599 <= reg_q2599_init;
        else
          reg_q2599 <= reg_q2599_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2016_in <= (reg_q2014 AND symb_decoder(16#46#)) OR
 					(reg_q2014 AND symb_decoder(16#66#));
reg_q2016_init <= '0' ;
	p_reg_q2016: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2016 <= reg_q2016_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2016 <= reg_q2016_init;
        else
          reg_q2016 <= reg_q2016_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2018_in <= (reg_q2016 AND symb_decoder(16#65#)) OR
 					(reg_q2016 AND symb_decoder(16#45#));
reg_q2018_init <= '0' ;
	p_reg_q2018: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2018 <= reg_q2018_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2018 <= reg_q2018_init;
        else
          reg_q2018 <= reg_q2018_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1989_in <= (reg_q1989 AND symb_decoder(16#36#)) OR
 					(reg_q1989 AND symb_decoder(16#33#)) OR
 					(reg_q1989 AND symb_decoder(16#30#)) OR
 					(reg_q1989 AND symb_decoder(16#35#)) OR
 					(reg_q1989 AND symb_decoder(16#38#)) OR
 					(reg_q1989 AND symb_decoder(16#37#)) OR
 					(reg_q1989 AND symb_decoder(16#31#)) OR
 					(reg_q1989 AND symb_decoder(16#34#)) OR
 					(reg_q1989 AND symb_decoder(16#39#)) OR
 					(reg_q1989 AND symb_decoder(16#32#)) OR
 					(reg_q1987 AND symb_decoder(16#30#)) OR
 					(reg_q1987 AND symb_decoder(16#31#)) OR
 					(reg_q1987 AND symb_decoder(16#39#)) OR
 					(reg_q1987 AND symb_decoder(16#33#)) OR
 					(reg_q1987 AND symb_decoder(16#34#)) OR
 					(reg_q1987 AND symb_decoder(16#37#)) OR
 					(reg_q1987 AND symb_decoder(16#36#)) OR
 					(reg_q1987 AND symb_decoder(16#38#)) OR
 					(reg_q1987 AND symb_decoder(16#32#)) OR
 					(reg_q1987 AND symb_decoder(16#35#));
reg_q1989_init <= '0' ;
	p_reg_q1989: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1989 <= reg_q1989_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1989 <= reg_q1989_init;
        else
          reg_q1989 <= reg_q1989_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2543_in <= (reg_q2541 AND symb_decoder(16#2c#));
reg_q2543_init <= '0' ;
	p_reg_q2543: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2543 <= reg_q2543_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2543 <= reg_q2543_init;
        else
          reg_q2543 <= reg_q2543_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2545_in <= (reg_q2543 AND symb_decoder(16#52#)) OR
 					(reg_q2543 AND symb_decoder(16#72#));
reg_q2545_init <= '0' ;
	p_reg_q2545: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2545 <= reg_q2545_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2545 <= reg_q2545_init;
        else
          reg_q2545 <= reg_q2545_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1728_in <= (reg_q1726 AND symb_decoder(16#52#)) OR
 					(reg_q1726 AND symb_decoder(16#72#));
reg_q1728_init <= '0' ;
	p_reg_q1728: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1728 <= reg_q1728_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1728 <= reg_q1728_init;
        else
          reg_q1728 <= reg_q1728_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1730_in <= (reg_q1728 AND symb_decoder(16#0d#)) OR
 					(reg_q1728 AND symb_decoder(16#09#)) OR
 					(reg_q1728 AND symb_decoder(16#20#)) OR
 					(reg_q1728 AND symb_decoder(16#0a#)) OR
 					(reg_q1728 AND symb_decoder(16#0c#)) OR
 					(reg_q1730 AND symb_decoder(16#09#)) OR
 					(reg_q1730 AND symb_decoder(16#0d#)) OR
 					(reg_q1730 AND symb_decoder(16#0c#)) OR
 					(reg_q1730 AND symb_decoder(16#20#)) OR
 					(reg_q1730 AND symb_decoder(16#0a#));
reg_q1730_init <= '0' ;
	p_reg_q1730: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1730 <= reg_q1730_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1730 <= reg_q1730_init;
        else
          reg_q1730 <= reg_q1730_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q438_in <= (reg_q436 AND symb_decoder(16#72#)) OR
 					(reg_q436 AND symb_decoder(16#52#));
reg_q438_init <= '0' ;
	p_reg_q438: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q438 <= reg_q438_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q438 <= reg_q438_init;
        else
          reg_q438 <= reg_q438_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q440_in <= (reg_q438 AND symb_decoder(16#0d#)) OR
 					(reg_q438 AND symb_decoder(16#0a#)) OR
 					(reg_q438 AND symb_decoder(16#0c#)) OR
 					(reg_q438 AND symb_decoder(16#09#)) OR
 					(reg_q438 AND symb_decoder(16#20#)) OR
 					(reg_q440 AND symb_decoder(16#0a#)) OR
 					(reg_q440 AND symb_decoder(16#20#)) OR
 					(reg_q440 AND symb_decoder(16#09#)) OR
 					(reg_q440 AND symb_decoder(16#0d#)) OR
 					(reg_q440 AND symb_decoder(16#0c#));
reg_q440_init <= '0' ;
	p_reg_q440: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q440 <= reg_q440_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q440 <= reg_q440_init;
        else
          reg_q440 <= reg_q440_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q772_in <= (reg_q770 AND symb_decoder(16#72#)) OR
 					(reg_q770 AND symb_decoder(16#52#));
reg_q772_init <= '0' ;
	p_reg_q772: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q772 <= reg_q772_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q772 <= reg_q772_init;
        else
          reg_q772 <= reg_q772_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q774_in <= (reg_q772 AND symb_decoder(16#59#)) OR
 					(reg_q772 AND symb_decoder(16#79#));
reg_q774_init <= '0' ;
	p_reg_q774: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q774 <= reg_q774_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q774 <= reg_q774_init;
        else
          reg_q774 <= reg_q774_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2630_in <= (reg_q2628 AND symb_decoder(16#55#)) OR
 					(reg_q2628 AND symb_decoder(16#75#));
reg_q2630_init <= '0' ;
	p_reg_q2630: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2630 <= reg_q2630_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2630 <= reg_q2630_init;
        else
          reg_q2630 <= reg_q2630_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2632_in <= (reg_q2630 AND symb_decoder(16#73#)) OR
 					(reg_q2630 AND symb_decoder(16#53#));
reg_q2632_init <= '0' ;
	p_reg_q2632: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2632 <= reg_q2632_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2632 <= reg_q2632_init;
        else
          reg_q2632 <= reg_q2632_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q528_in <= (reg_q526 AND symb_decoder(16#2e#));
reg_q528_init <= '0' ;
	p_reg_q528: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q528 <= reg_q528_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q528 <= reg_q528_init;
        else
          reg_q528 <= reg_q528_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1963_in <= (reg_q1961 AND symb_decoder(16#53#)) OR
 					(reg_q1961 AND symb_decoder(16#73#));
reg_q1963_init <= '0' ;
	p_reg_q1963: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1963 <= reg_q1963_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1963 <= reg_q1963_init;
        else
          reg_q1963 <= reg_q1963_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1965_in <= (reg_q1963 AND symb_decoder(16#45#)) OR
 					(reg_q1963 AND symb_decoder(16#65#));
reg_q1965_init <= '0' ;
	p_reg_q1965: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1965 <= reg_q1965_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1965 <= reg_q1965_init;
        else
          reg_q1965 <= reg_q1965_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1264_in <= (reg_q1262 AND symb_decoder(16#45#)) OR
 					(reg_q1262 AND symb_decoder(16#65#));
reg_q1264_init <= '0' ;
	p_reg_q1264: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1264 <= reg_q1264_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1264 <= reg_q1264_init;
        else
          reg_q1264 <= reg_q1264_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1266_in <= (reg_q1264 AND symb_decoder(16#72#)) OR
 					(reg_q1264 AND symb_decoder(16#52#));
reg_q1266_init <= '0' ;
	p_reg_q1266: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1266 <= reg_q1266_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1266 <= reg_q1266_init;
        else
          reg_q1266 <= reg_q1266_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q255_in <= (reg_q253 AND symb_decoder(16#ff#));
reg_q255_init <= '0' ;
	p_reg_q255: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q255 <= reg_q255_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q255 <= reg_q255_init;
        else
          reg_q255 <= reg_q255_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q596_in <= (reg_q596 AND symb_decoder(16#0a#)) OR
 					(reg_q596 AND symb_decoder(16#20#)) OR
 					(reg_q596 AND symb_decoder(16#0c#)) OR
 					(reg_q596 AND symb_decoder(16#09#)) OR
 					(reg_q596 AND symb_decoder(16#0d#)) OR
 					(reg_q594 AND symb_decoder(16#0a#)) OR
 					(reg_q594 AND symb_decoder(16#0c#)) OR
 					(reg_q594 AND symb_decoder(16#0d#)) OR
 					(reg_q594 AND symb_decoder(16#09#)) OR
 					(reg_q594 AND symb_decoder(16#20#));
reg_q596_init <= '0' ;
	p_reg_q596: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q596 <= reg_q596_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q596 <= reg_q596_init;
        else
          reg_q596 <= reg_q596_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q245_in <= (reg_q245 AND symb_decoder(16#36#)) OR
 					(reg_q245 AND symb_decoder(16#31#)) OR
 					(reg_q245 AND symb_decoder(16#32#)) OR
 					(reg_q245 AND symb_decoder(16#35#)) OR
 					(reg_q245 AND symb_decoder(16#33#)) OR
 					(reg_q245 AND symb_decoder(16#38#)) OR
 					(reg_q245 AND symb_decoder(16#37#)) OR
 					(reg_q245 AND symb_decoder(16#30#)) OR
 					(reg_q245 AND symb_decoder(16#39#)) OR
 					(reg_q245 AND symb_decoder(16#34#)) OR
 					(reg_q243 AND symb_decoder(16#35#)) OR
 					(reg_q243 AND symb_decoder(16#39#)) OR
 					(reg_q243 AND symb_decoder(16#36#)) OR
 					(reg_q243 AND symb_decoder(16#38#)) OR
 					(reg_q243 AND symb_decoder(16#32#)) OR
 					(reg_q243 AND symb_decoder(16#30#)) OR
 					(reg_q243 AND symb_decoder(16#33#)) OR
 					(reg_q243 AND symb_decoder(16#34#)) OR
 					(reg_q243 AND symb_decoder(16#31#)) OR
 					(reg_q243 AND symb_decoder(16#37#));
reg_q245_init <= '0' ;
	p_reg_q245: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q245 <= reg_q245_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q245 <= reg_q245_init;
        else
          reg_q245 <= reg_q245_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2160_in <= (reg_q2158 AND symb_decoder(16#0a#)) OR
 					(reg_q2158 AND symb_decoder(16#09#)) OR
 					(reg_q2158 AND symb_decoder(16#0c#)) OR
 					(reg_q2158 AND symb_decoder(16#0d#)) OR
 					(reg_q2158 AND symb_decoder(16#20#)) OR
 					(reg_q2160 AND symb_decoder(16#0a#)) OR
 					(reg_q2160 AND symb_decoder(16#0c#)) OR
 					(reg_q2160 AND symb_decoder(16#09#)) OR
 					(reg_q2160 AND symb_decoder(16#20#)) OR
 					(reg_q2160 AND symb_decoder(16#0d#));
reg_q2160_init <= '0' ;
	p_reg_q2160: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2160 <= reg_q2160_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2160 <= reg_q2160_init;
        else
          reg_q2160 <= reg_q2160_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2573_in <= (reg_q2571 AND symb_decoder(16#45#)) OR
 					(reg_q2571 AND symb_decoder(16#65#));
reg_q2573_init <= '0' ;
	p_reg_q2573: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2573 <= reg_q2573_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2573 <= reg_q2573_init;
        else
          reg_q2573 <= reg_q2573_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1648_in <= (reg_q1646 AND symb_decoder(16#74#)) OR
 					(reg_q1646 AND symb_decoder(16#54#));
reg_q1648_init <= '0' ;
	p_reg_q1648: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1648 <= reg_q1648_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1648 <= reg_q1648_init;
        else
          reg_q1648 <= reg_q1648_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1650_in <= (reg_q1648 AND symb_decoder(16#62#)) OR
 					(reg_q1648 AND symb_decoder(16#42#));
reg_q1650_init <= '0' ;
	p_reg_q1650: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1650 <= reg_q1650_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1650 <= reg_q1650_init;
        else
          reg_q1650 <= reg_q1650_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2480_in <= (reg_q2478 AND symb_decoder(16#2a#));
reg_q2480_init <= '0' ;
	p_reg_q2480: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2480 <= reg_q2480_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2480 <= reg_q2480_init;
        else
          reg_q2480 <= reg_q2480_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2482_in <= (reg_q2480 AND symb_decoder(16#38#)) OR
 					(reg_q2480 AND symb_decoder(16#37#)) OR
 					(reg_q2480 AND symb_decoder(16#36#)) OR
 					(reg_q2480 AND symb_decoder(16#39#)) OR
 					(reg_q2480 AND symb_decoder(16#34#)) OR
 					(reg_q2480 AND symb_decoder(16#32#)) OR
 					(reg_q2480 AND symb_decoder(16#35#)) OR
 					(reg_q2480 AND symb_decoder(16#33#)) OR
 					(reg_q2480 AND symb_decoder(16#30#)) OR
 					(reg_q2480 AND symb_decoder(16#31#)) OR
 					(reg_q2482 AND symb_decoder(16#33#)) OR
 					(reg_q2482 AND symb_decoder(16#39#)) OR
 					(reg_q2482 AND symb_decoder(16#35#)) OR
 					(reg_q2482 AND symb_decoder(16#38#)) OR
 					(reg_q2482 AND symb_decoder(16#37#)) OR
 					(reg_q2482 AND symb_decoder(16#34#)) OR
 					(reg_q2482 AND symb_decoder(16#30#)) OR
 					(reg_q2482 AND symb_decoder(16#36#)) OR
 					(reg_q2482 AND symb_decoder(16#32#)) OR
 					(reg_q2482 AND symb_decoder(16#31#));
reg_q2482_init <= '0' ;
	p_reg_q2482: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2482 <= reg_q2482_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2482 <= reg_q2482_init;
        else
          reg_q2482 <= reg_q2482_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q107_in <= (reg_q105 AND symb_decoder(16#49#)) OR
 					(reg_q105 AND symb_decoder(16#69#));
reg_q107_init <= '0' ;
	p_reg_q107: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q107 <= reg_q107_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q107 <= reg_q107_init;
        else
          reg_q107 <= reg_q107_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q109_in <= (reg_q107 AND symb_decoder(16#78#)) OR
 					(reg_q107 AND symb_decoder(16#58#));
reg_q109_init <= '0' ;
	p_reg_q109: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q109 <= reg_q109_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q109 <= reg_q109_init;
        else
          reg_q109 <= reg_q109_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1213_in <= (reg_q1211 AND symb_decoder(16#69#)) OR
 					(reg_q1211 AND symb_decoder(16#49#));
reg_q1213_init <= '0' ;
	p_reg_q1213: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1213 <= reg_q1213_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1213 <= reg_q1213_init;
        else
          reg_q1213 <= reg_q1213_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1215_in <= (reg_q1213 AND symb_decoder(16#6d#)) OR
 					(reg_q1213 AND symb_decoder(16#4d#));
reg_q1215_init <= '0' ;
	p_reg_q1215: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1215 <= reg_q1215_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1215 <= reg_q1215_init;
        else
          reg_q1215 <= reg_q1215_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2355_in <= (reg_q2353 AND symb_decoder(16#61#)) OR
 					(reg_q2353 AND symb_decoder(16#41#));
reg_q2355_init <= '0' ;
	p_reg_q2355: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2355 <= reg_q2355_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2355 <= reg_q2355_init;
        else
          reg_q2355 <= reg_q2355_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2357_in <= (reg_q2355 AND symb_decoder(16#6e#)) OR
 					(reg_q2355 AND symb_decoder(16#4e#));
reg_q2357_init <= '0' ;
	p_reg_q2357: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2357 <= reg_q2357_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2357 <= reg_q2357_init;
        else
          reg_q2357 <= reg_q2357_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1609_in <= (reg_q1607 AND symb_decoder(16#43#)) OR
 					(reg_q1607 AND symb_decoder(16#63#));
reg_q1609_init <= '0' ;
	p_reg_q1609: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1609 <= reg_q1609_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1609 <= reg_q1609_init;
        else
          reg_q1609 <= reg_q1609_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1611_in <= (reg_q1609 AND symb_decoder(16#6b#)) OR
 					(reg_q1609 AND symb_decoder(16#4b#));
reg_q1611_init <= '0' ;
	p_reg_q1611: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1611 <= reg_q1611_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1611 <= reg_q1611_init;
        else
          reg_q1611 <= reg_q1611_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2092_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2091 AND symb_decoder(16#0a#)) OR
 					(reg_q2091 AND symb_decoder(16#0d#));
reg_q2092_init <= '0' ;
	p_reg_q2092: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2092 <= reg_q2092_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2092 <= reg_q2092_init;
        else
          reg_q2092 <= reg_q2092_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1613_in <= (reg_q1611 AND symb_decoder(16#0d#)) OR
 					(reg_q1611 AND symb_decoder(16#0c#)) OR
 					(reg_q1611 AND symb_decoder(16#09#)) OR
 					(reg_q1611 AND symb_decoder(16#0a#)) OR
 					(reg_q1611 AND symb_decoder(16#20#)) OR
 					(reg_q1613 AND symb_decoder(16#09#)) OR
 					(reg_q1613 AND symb_decoder(16#0d#)) OR
 					(reg_q1613 AND symb_decoder(16#0c#)) OR
 					(reg_q1613 AND symb_decoder(16#20#)) OR
 					(reg_q1613 AND symb_decoder(16#0a#));
reg_q1613_init <= '0' ;
	p_reg_q1613: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1613 <= reg_q1613_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1613 <= reg_q1613_init;
        else
          reg_q1613 <= reg_q1613_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2152_in <= (reg_q2150 AND symb_decoder(16#52#)) OR
 					(reg_q2150 AND symb_decoder(16#72#));
reg_q2152_init <= '0' ;
	p_reg_q2152: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2152 <= reg_q2152_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2152 <= reg_q2152_init;
        else
          reg_q2152 <= reg_q2152_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2154_in <= (reg_q2152 AND symb_decoder(16#65#)) OR
 					(reg_q2152 AND symb_decoder(16#45#));
reg_q2154_init <= '0' ;
	p_reg_q2154: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2154 <= reg_q2154_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2154 <= reg_q2154_init;
        else
          reg_q2154 <= reg_q2154_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1460_in <= (reg_q1458 AND symb_decoder(16#54#)) OR
 					(reg_q1458 AND symb_decoder(16#74#));
reg_q1460_init <= '0' ;
	p_reg_q1460: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1460 <= reg_q1460_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1460 <= reg_q1460_init;
        else
          reg_q1460 <= reg_q1460_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1339_in <= (reg_q1339 AND symb_decoder(16#36#)) OR
 					(reg_q1339 AND symb_decoder(16#35#)) OR
 					(reg_q1339 AND symb_decoder(16#39#)) OR
 					(reg_q1339 AND symb_decoder(16#30#)) OR
 					(reg_q1339 AND symb_decoder(16#38#)) OR
 					(reg_q1339 AND symb_decoder(16#34#)) OR
 					(reg_q1339 AND symb_decoder(16#31#)) OR
 					(reg_q1339 AND symb_decoder(16#32#)) OR
 					(reg_q1339 AND symb_decoder(16#33#)) OR
 					(reg_q1339 AND symb_decoder(16#37#)) OR
 					(reg_q1337 AND symb_decoder(16#35#)) OR
 					(reg_q1337 AND symb_decoder(16#36#)) OR
 					(reg_q1337 AND symb_decoder(16#31#)) OR
 					(reg_q1337 AND symb_decoder(16#39#)) OR
 					(reg_q1337 AND symb_decoder(16#32#)) OR
 					(reg_q1337 AND symb_decoder(16#30#)) OR
 					(reg_q1337 AND symb_decoder(16#38#)) OR
 					(reg_q1337 AND symb_decoder(16#37#)) OR
 					(reg_q1337 AND symb_decoder(16#33#)) OR
 					(reg_q1337 AND symb_decoder(16#34#));
reg_q1339_init <= '0' ;
	p_reg_q1339: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1339 <= reg_q1339_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1339 <= reg_q1339_init;
        else
          reg_q1339 <= reg_q1339_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2528_in <= (reg_q2526 AND symb_decoder(16#3b#));
reg_q2528_init <= '0' ;
	p_reg_q2528: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2528 <= reg_q2528_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2528 <= reg_q2528_init;
        else
          reg_q2528 <= reg_q2528_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q694_in <= (reg_q692 AND symb_decoder(16#2e#));
reg_q694_init <= '0' ;
	p_reg_q694: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q694 <= reg_q694_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q694 <= reg_q694_init;
        else
          reg_q694 <= reg_q694_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1578_in <= (reg_q1576 AND symb_decoder(16#2e#));
reg_q1578_init <= '0' ;
	p_reg_q1578: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1578 <= reg_q1578_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1578 <= reg_q1578_init;
        else
          reg_q1578 <= reg_q1578_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2520_in <= (reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2518 AND symb_decoder(16#2f#));
reg_q2520_init <= '0' ;
	p_reg_q2520: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2520 <= reg_q2520_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2520 <= reg_q2520_init;
        else
          reg_q2520 <= reg_q2520_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2042_in <= (reg_q2040 AND symb_decoder(16#66#)) OR
 					(reg_q2040 AND symb_decoder(16#46#));
reg_q2042_init <= '0' ;
	p_reg_q2042: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2042 <= reg_q2042_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2042 <= reg_q2042_init;
        else
          reg_q2042 <= reg_q2042_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2044_in <= (reg_q2042 AND symb_decoder(16#72#)) OR
 					(reg_q2042 AND symb_decoder(16#52#));
reg_q2044_init <= '0' ;
	p_reg_q2044: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2044 <= reg_q2044_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2044 <= reg_q2044_init;
        else
          reg_q2044 <= reg_q2044_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2524_in <= (reg_q2522 AND symb_decoder(16#52#)) OR
 					(reg_q2522 AND symb_decoder(16#72#));
reg_q2524_init <= '0' ;
	p_reg_q2524: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2524 <= reg_q2524_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2524 <= reg_q2524_init;
        else
          reg_q2524 <= reg_q2524_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2526_in <= (reg_q2524 AND symb_decoder(16#36#)) OR
 					(reg_q2524 AND symb_decoder(16#30#)) OR
 					(reg_q2524 AND symb_decoder(16#31#)) OR
 					(reg_q2524 AND symb_decoder(16#34#)) OR
 					(reg_q2524 AND symb_decoder(16#39#)) OR
 					(reg_q2524 AND symb_decoder(16#38#)) OR
 					(reg_q2524 AND symb_decoder(16#33#)) OR
 					(reg_q2524 AND symb_decoder(16#35#)) OR
 					(reg_q2524 AND symb_decoder(16#32#)) OR
 					(reg_q2524 AND symb_decoder(16#37#)) OR
 					(reg_q2526 AND symb_decoder(16#35#)) OR
 					(reg_q2526 AND symb_decoder(16#34#)) OR
 					(reg_q2526 AND symb_decoder(16#33#)) OR
 					(reg_q2526 AND symb_decoder(16#37#)) OR
 					(reg_q2526 AND symb_decoder(16#31#)) OR
 					(reg_q2526 AND symb_decoder(16#32#)) OR
 					(reg_q2526 AND symb_decoder(16#30#)) OR
 					(reg_q2526 AND symb_decoder(16#39#)) OR
 					(reg_q2526 AND symb_decoder(16#38#)) OR
 					(reg_q2526 AND symb_decoder(16#36#));
reg_q2526_init <= '0' ;
	p_reg_q2526: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2526 <= reg_q2526_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2526 <= reg_q2526_init;
        else
          reg_q2526 <= reg_q2526_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1272_in <= (reg_q1270 AND symb_decoder(16#72#)) OR
 					(reg_q1270 AND symb_decoder(16#52#));
reg_q1272_init <= '0' ;
	p_reg_q1272: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1272 <= reg_q1272_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1272 <= reg_q1272_init;
        else
          reg_q1272 <= reg_q1272_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1274_in <= (reg_q1272 AND symb_decoder(16#0a#)) OR
 					(reg_q1272 AND symb_decoder(16#09#)) OR
 					(reg_q1272 AND symb_decoder(16#0c#)) OR
 					(reg_q1272 AND symb_decoder(16#0d#)) OR
 					(reg_q1272 AND symb_decoder(16#20#)) OR
 					(reg_q1274 AND symb_decoder(16#09#)) OR
 					(reg_q1274 AND symb_decoder(16#0c#)) OR
 					(reg_q1274 AND symb_decoder(16#0a#)) OR
 					(reg_q1274 AND symb_decoder(16#20#)) OR
 					(reg_q1274 AND symb_decoder(16#0d#));
reg_q1274_init <= '0' ;
	p_reg_q1274: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1274 <= reg_q1274_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1274 <= reg_q1274_init;
        else
          reg_q1274 <= reg_q1274_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q111_in <= (reg_q109 AND symb_decoder(16#20#)) OR
 					(reg_q109 AND symb_decoder(16#0d#)) OR
 					(reg_q109 AND symb_decoder(16#0a#)) OR
 					(reg_q109 AND symb_decoder(16#0c#)) OR
 					(reg_q109 AND symb_decoder(16#09#)) OR
 					(reg_q111 AND symb_decoder(16#09#)) OR
 					(reg_q111 AND symb_decoder(16#0a#)) OR
 					(reg_q111 AND symb_decoder(16#0d#)) OR
 					(reg_q111 AND symb_decoder(16#20#)) OR
 					(reg_q111 AND symb_decoder(16#0c#));
reg_q111_init <= '0' ;
	p_reg_q111: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q111 <= reg_q111_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q111 <= reg_q111_init;
        else
          reg_q111 <= reg_q111_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q941_in <= (reg_q939 AND symb_decoder(16#2e#));
reg_q941_init <= '0' ;
	p_reg_q941: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q941 <= reg_q941_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q941 <= reg_q941_init;
        else
          reg_q941 <= reg_q941_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q943_in <= (reg_q941 AND symb_decoder(16#33#)) OR
 					(reg_q941 AND symb_decoder(16#37#)) OR
 					(reg_q941 AND symb_decoder(16#35#)) OR
 					(reg_q941 AND symb_decoder(16#30#)) OR
 					(reg_q941 AND symb_decoder(16#32#)) OR
 					(reg_q941 AND symb_decoder(16#34#)) OR
 					(reg_q941 AND symb_decoder(16#38#)) OR
 					(reg_q941 AND symb_decoder(16#36#)) OR
 					(reg_q941 AND symb_decoder(16#39#)) OR
 					(reg_q941 AND symb_decoder(16#31#)) OR
 					(reg_q943 AND symb_decoder(16#38#)) OR
 					(reg_q943 AND symb_decoder(16#35#)) OR
 					(reg_q943 AND symb_decoder(16#37#)) OR
 					(reg_q943 AND symb_decoder(16#32#)) OR
 					(reg_q943 AND symb_decoder(16#34#)) OR
 					(reg_q943 AND symb_decoder(16#31#)) OR
 					(reg_q943 AND symb_decoder(16#30#)) OR
 					(reg_q943 AND symb_decoder(16#39#)) OR
 					(reg_q943 AND symb_decoder(16#33#)) OR
 					(reg_q943 AND symb_decoder(16#36#));
reg_q943_init <= '0' ;
	p_reg_q943: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q943 <= reg_q943_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q943 <= reg_q943_init;
        else
          reg_q943 <= reg_q943_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q709_in <= (reg_q707 AND symb_decoder(16#0d#)) OR
 					(reg_q707 AND symb_decoder(16#0c#)) OR
 					(reg_q707 AND symb_decoder(16#0a#)) OR
 					(reg_q707 AND symb_decoder(16#20#)) OR
 					(reg_q707 AND symb_decoder(16#09#));
reg_q709_init <= '0' ;
	p_reg_q709: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q709 <= reg_q709_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q709 <= reg_q709_init;
        else
          reg_q709 <= reg_q709_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q711_in <= (reg_q709 AND symb_decoder(16#37#)) OR
 					(reg_q709 AND symb_decoder(16#30#)) OR
 					(reg_q709 AND symb_decoder(16#31#)) OR
 					(reg_q709 AND symb_decoder(16#39#)) OR
 					(reg_q709 AND symb_decoder(16#34#)) OR
 					(reg_q709 AND symb_decoder(16#36#)) OR
 					(reg_q709 AND symb_decoder(16#32#)) OR
 					(reg_q709 AND symb_decoder(16#35#)) OR
 					(reg_q709 AND symb_decoder(16#38#)) OR
 					(reg_q709 AND symb_decoder(16#33#)) OR
 					(reg_q711 AND symb_decoder(16#30#)) OR
 					(reg_q711 AND symb_decoder(16#39#)) OR
 					(reg_q711 AND symb_decoder(16#31#)) OR
 					(reg_q711 AND symb_decoder(16#33#)) OR
 					(reg_q711 AND symb_decoder(16#37#)) OR
 					(reg_q711 AND symb_decoder(16#34#)) OR
 					(reg_q711 AND symb_decoder(16#32#)) OR
 					(reg_q711 AND symb_decoder(16#35#)) OR
 					(reg_q711 AND symb_decoder(16#36#)) OR
 					(reg_q711 AND symb_decoder(16#38#));
reg_q711_init <= '0' ;
	p_reg_q711: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q711 <= reg_q711_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q711 <= reg_q711_init;
        else
          reg_q711 <= reg_q711_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1226_in <= (reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1225 AND symb_decoder(16#67#)) OR
 					(reg_q1225 AND symb_decoder(16#47#));
reg_q1226_init <= '0' ;
	p_reg_q1226: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1226 <= reg_q1226_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1226 <= reg_q1226_init;
        else
          reg_q1226 <= reg_q1226_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1228_in <= (reg_q1226 AND symb_decoder(16#61#)) OR
 					(reg_q1226 AND symb_decoder(16#41#));
reg_q1228_init <= '0' ;
	p_reg_q1228: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1228 <= reg_q1228_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1228 <= reg_q1228_init;
        else
          reg_q1228 <= reg_q1228_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q101_in <= (reg_q99 AND symb_decoder(16#6f#)) OR
 					(reg_q99 AND symb_decoder(16#4f#));
reg_q101_init <= '0' ;
	p_reg_q101: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q101 <= reg_q101_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q101 <= reg_q101_init;
        else
          reg_q101 <= reg_q101_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q103_in <= (reg_q101 AND symb_decoder(16#70#)) OR
 					(reg_q101 AND symb_decoder(16#50#));
reg_q103_init <= '0' ;
	p_reg_q103: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q103 <= reg_q103_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q103 <= reg_q103_init;
        else
          reg_q103 <= reg_q103_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q237_in <= (reg_q237 AND symb_decoder(16#38#)) OR
 					(reg_q237 AND symb_decoder(16#35#)) OR
 					(reg_q237 AND symb_decoder(16#36#)) OR
 					(reg_q237 AND symb_decoder(16#37#)) OR
 					(reg_q237 AND symb_decoder(16#30#)) OR
 					(reg_q237 AND symb_decoder(16#39#)) OR
 					(reg_q237 AND symb_decoder(16#34#)) OR
 					(reg_q237 AND symb_decoder(16#31#)) OR
 					(reg_q237 AND symb_decoder(16#33#)) OR
 					(reg_q237 AND symb_decoder(16#32#)) OR
 					(reg_q235 AND symb_decoder(16#31#)) OR
 					(reg_q235 AND symb_decoder(16#36#)) OR
 					(reg_q235 AND symb_decoder(16#35#)) OR
 					(reg_q235 AND symb_decoder(16#37#)) OR
 					(reg_q235 AND symb_decoder(16#30#)) OR
 					(reg_q235 AND symb_decoder(16#38#)) OR
 					(reg_q235 AND symb_decoder(16#39#)) OR
 					(reg_q235 AND symb_decoder(16#32#)) OR
 					(reg_q235 AND symb_decoder(16#33#)) OR
 					(reg_q235 AND symb_decoder(16#34#));
reg_q237_init <= '0' ;
	p_reg_q237: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q237 <= reg_q237_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q237 <= reg_q237_init;
        else
          reg_q237 <= reg_q237_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q226_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q225 AND symb_decoder(16#0a#)) OR
 					(reg_q225 AND symb_decoder(16#0d#));
reg_q226_init <= '0' ;
	p_reg_q226: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q226 <= reg_q226_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q226 <= reg_q226_init;
        else
          reg_q226 <= reg_q226_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q937_in <= (reg_q933 AND symb_decoder(16#00#)) OR
 					(reg_q955 AND symb_decoder(16#00#));
reg_q937_init <= '0' ;
	p_reg_q937: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q937 <= reg_q937_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q937 <= reg_q937_init;
        else
          reg_q937 <= reg_q937_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q939_in <= (reg_q937 AND symb_decoder(16#36#)) OR
 					(reg_q937 AND symb_decoder(16#35#)) OR
 					(reg_q937 AND symb_decoder(16#31#)) OR
 					(reg_q937 AND symb_decoder(16#33#)) OR
 					(reg_q937 AND symb_decoder(16#34#)) OR
 					(reg_q937 AND symb_decoder(16#30#)) OR
 					(reg_q937 AND symb_decoder(16#39#)) OR
 					(reg_q937 AND symb_decoder(16#38#)) OR
 					(reg_q937 AND symb_decoder(16#32#)) OR
 					(reg_q937 AND symb_decoder(16#37#)) OR
 					(reg_q939 AND symb_decoder(16#31#)) OR
 					(reg_q939 AND symb_decoder(16#37#)) OR
 					(reg_q939 AND symb_decoder(16#35#)) OR
 					(reg_q939 AND symb_decoder(16#30#)) OR
 					(reg_q939 AND symb_decoder(16#34#)) OR
 					(reg_q939 AND symb_decoder(16#32#)) OR
 					(reg_q939 AND symb_decoder(16#38#)) OR
 					(reg_q939 AND symb_decoder(16#33#)) OR
 					(reg_q939 AND symb_decoder(16#36#)) OR
 					(reg_q939 AND symb_decoder(16#39#));
reg_q939_init <= '0' ;
	p_reg_q939: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q939 <= reg_q939_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q939 <= reg_q939_init;
        else
          reg_q939 <= reg_q939_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q321_in <= (reg_q319 AND symb_decoder(16#00#));
reg_q321_init <= '0' ;
	p_reg_q321: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q321 <= reg_q321_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q321 <= reg_q321_init;
        else
          reg_q321 <= reg_q321_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q323_in <= (reg_q321 AND symb_decoder(16#00#));
reg_q323_init <= '0' ;
	p_reg_q323: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q323 <= reg_q323_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q323 <= reg_q323_init;
        else
          reg_q323 <= reg_q323_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2253_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2252 AND symb_decoder(16#0a#)) OR
 					(reg_q2252 AND symb_decoder(16#0d#));
reg_q2253_init <= '0' ;
	p_reg_q2253: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2253 <= reg_q2253_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2253 <= reg_q2253_init;
        else
          reg_q2253 <= reg_q2253_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2178_in <= (reg_q2176 AND symb_decoder(16#49#)) OR
 					(reg_q2176 AND symb_decoder(16#69#));
reg_q2178_init <= '0' ;
	p_reg_q2178: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2178 <= reg_q2178_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2178 <= reg_q2178_init;
        else
          reg_q2178 <= reg_q2178_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2180_in <= (reg_q2178 AND symb_decoder(16#63#)) OR
 					(reg_q2178 AND symb_decoder(16#43#));
reg_q2180_init <= '0' ;
	p_reg_q2180: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2180 <= reg_q2180_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2180 <= reg_q2180_init;
        else
          reg_q2180 <= reg_q2180_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2565_in <= (reg_q2565 AND symb_decoder(16#09#)) OR
 					(reg_q2565 AND symb_decoder(16#0c#)) OR
 					(reg_q2565 AND symb_decoder(16#20#)) OR
 					(reg_q2565 AND symb_decoder(16#0d#)) OR
 					(reg_q2565 AND symb_decoder(16#0a#)) OR
 					(reg_q2563 AND symb_decoder(16#0d#)) OR
 					(reg_q2563 AND symb_decoder(16#20#)) OR
 					(reg_q2563 AND symb_decoder(16#09#)) OR
 					(reg_q2563 AND symb_decoder(16#0c#)) OR
 					(reg_q2563 AND symb_decoder(16#0a#));
reg_q2565_init <= '0' ;
	p_reg_q2565: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2565 <= reg_q2565_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2565 <= reg_q2565_init;
        else
          reg_q2565 <= reg_q2565_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1443_in <= (reg_q1441 AND symb_decoder(16#73#)) OR
 					(reg_q1441 AND symb_decoder(16#53#));
reg_q1443_init <= '0' ;
	p_reg_q1443: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1443 <= reg_q1443_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1443 <= reg_q1443_init;
        else
          reg_q1443 <= reg_q1443_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1445_in <= (reg_q1443 AND symb_decoder(16#54#)) OR
 					(reg_q1443 AND symb_decoder(16#74#));
reg_q1445_init <= '0' ;
	p_reg_q1445: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1445 <= reg_q1445_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1445 <= reg_q1445_init;
        else
          reg_q1445 <= reg_q1445_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2148_in <= (reg_q2148 AND symb_decoder(16#0a#)) OR
 					(reg_q2148 AND symb_decoder(16#20#)) OR
 					(reg_q2148 AND symb_decoder(16#0c#)) OR
 					(reg_q2148 AND symb_decoder(16#09#)) OR
 					(reg_q2148 AND symb_decoder(16#0d#)) OR
 					(reg_q2146 AND symb_decoder(16#0a#)) OR
 					(reg_q2146 AND symb_decoder(16#09#)) OR
 					(reg_q2146 AND symb_decoder(16#0d#)) OR
 					(reg_q2146 AND symb_decoder(16#20#)) OR
 					(reg_q2146 AND symb_decoder(16#0c#));
reg_q2148_init <= '0' ;
	p_reg_q2148: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2148 <= reg_q2148_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2148 <= reg_q2148_init;
        else
          reg_q2148 <= reg_q2148_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q590_in <= (reg_q588 AND symb_decoder(16#74#)) OR
 					(reg_q588 AND symb_decoder(16#54#));
reg_q590_init <= '0' ;
	p_reg_q590: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q590 <= reg_q590_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q590 <= reg_q590_init;
        else
          reg_q590 <= reg_q590_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q592_in <= (reg_q590 AND symb_decoder(16#69#)) OR
 					(reg_q590 AND symb_decoder(16#49#));
reg_q592_init <= '0' ;
	p_reg_q592: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q592 <= reg_q592_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q592 <= reg_q592_init;
        else
          reg_q592 <= reg_q592_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q949_in <= (reg_q947 AND symb_decoder(16#2e#));
reg_q949_init <= '0' ;
	p_reg_q949: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q949 <= reg_q949_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q949 <= reg_q949_init;
        else
          reg_q949 <= reg_q949_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q951_in <= (reg_q949 AND symb_decoder(16#35#)) OR
 					(reg_q949 AND symb_decoder(16#36#)) OR
 					(reg_q949 AND symb_decoder(16#37#)) OR
 					(reg_q949 AND symb_decoder(16#34#)) OR
 					(reg_q949 AND symb_decoder(16#30#)) OR
 					(reg_q949 AND symb_decoder(16#32#)) OR
 					(reg_q949 AND symb_decoder(16#31#)) OR
 					(reg_q949 AND symb_decoder(16#33#)) OR
 					(reg_q949 AND symb_decoder(16#39#)) OR
 					(reg_q949 AND symb_decoder(16#38#)) OR
 					(reg_q951 AND symb_decoder(16#31#)) OR
 					(reg_q951 AND symb_decoder(16#38#)) OR
 					(reg_q951 AND symb_decoder(16#37#)) OR
 					(reg_q951 AND symb_decoder(16#39#)) OR
 					(reg_q951 AND symb_decoder(16#35#)) OR
 					(reg_q951 AND symb_decoder(16#36#)) OR
 					(reg_q951 AND symb_decoder(16#30#)) OR
 					(reg_q951 AND symb_decoder(16#33#)) OR
 					(reg_q951 AND symb_decoder(16#32#)) OR
 					(reg_q951 AND symb_decoder(16#34#));
reg_q951_init <= '0' ;
	p_reg_q951: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q951 <= reg_q951_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q951 <= reg_q951_init;
        else
          reg_q951 <= reg_q951_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1660_in <= (reg_q1660 AND symb_decoder(16#0a#)) OR
 					(reg_q1660 AND symb_decoder(16#0c#)) OR
 					(reg_q1660 AND symb_decoder(16#09#)) OR
 					(reg_q1660 AND symb_decoder(16#0d#)) OR
 					(reg_q1660 AND symb_decoder(16#20#)) OR
 					(reg_q1658 AND symb_decoder(16#20#)) OR
 					(reg_q1658 AND symb_decoder(16#09#)) OR
 					(reg_q1658 AND symb_decoder(16#0a#)) OR
 					(reg_q1658 AND symb_decoder(16#0d#)) OR
 					(reg_q1658 AND symb_decoder(16#0c#));
reg_q1660_init <= '0' ;
	p_reg_q1660: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1660 <= reg_q1660_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1660 <= reg_q1660_init;
        else
          reg_q1660 <= reg_q1660_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1113_in <= (reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q1112 AND symb_decoder(16#66#)) OR
 					(reg_q1112 AND symb_decoder(16#46#));
reg_q1113_init <= '0' ;
	p_reg_q1113: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1113 <= reg_q1113_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1113 <= reg_q1113_init;
        else
          reg_q1113 <= reg_q1113_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q974_in <= (reg_q972 AND symb_decoder(16#6f#)) OR
 					(reg_q972 AND symb_decoder(16#4f#));
reg_q974_init <= '0' ;
	p_reg_q974: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q974 <= reg_q974_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q974 <= reg_q974_init;
        else
          reg_q974 <= reg_q974_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q976_in <= (reg_q974 AND symb_decoder(16#4d#)) OR
 					(reg_q974 AND symb_decoder(16#6d#));
reg_q976_init <= '0' ;
	p_reg_q976: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q976 <= reg_q976_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q976 <= reg_q976_init;
        else
          reg_q976 <= reg_q976_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q84_in <= (reg_q82 AND symb_decoder(16#52#)) OR
 					(reg_q82 AND symb_decoder(16#72#));
reg_q84_init <= '0' ;
	p_reg_q84: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q84 <= reg_q84_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q84 <= reg_q84_init;
        else
          reg_q84 <= reg_q84_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1902_in <= (reg_q1900 AND symb_decoder(16#54#)) OR
 					(reg_q1900 AND symb_decoder(16#74#));
reg_q1902_init <= '0' ;
	p_reg_q1902: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1902 <= reg_q1902_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1902 <= reg_q1902_init;
        else
          reg_q1902 <= reg_q1902_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1904_in <= (reg_q1902 AND symb_decoder(16#0d#)) OR
 					(reg_q1902 AND symb_decoder(16#0a#)) OR
 					(reg_q1902 AND symb_decoder(16#09#)) OR
 					(reg_q1902 AND symb_decoder(16#0c#)) OR
 					(reg_q1902 AND symb_decoder(16#20#)) OR
 					(reg_q1904 AND symb_decoder(16#0a#)) OR
 					(reg_q1904 AND symb_decoder(16#0d#)) OR
 					(reg_q1904 AND symb_decoder(16#09#)) OR
 					(reg_q1904 AND symb_decoder(16#20#)) OR
 					(reg_q1904 AND symb_decoder(16#0c#));
reg_q1904_init <= '0' ;
	p_reg_q1904: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1904 <= reg_q1904_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1904 <= reg_q1904_init;
        else
          reg_q1904 <= reg_q1904_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2613_in <= (reg_q2613 AND symb_decoder(16#09#)) OR
 					(reg_q2613 AND symb_decoder(16#0d#)) OR
 					(reg_q2613 AND symb_decoder(16#20#)) OR
 					(reg_q2613 AND symb_decoder(16#0c#)) OR
 					(reg_q2613 AND symb_decoder(16#0a#)) OR
 					(reg_q2611 AND symb_decoder(16#0a#)) OR
 					(reg_q2611 AND symb_decoder(16#0c#)) OR
 					(reg_q2611 AND symb_decoder(16#0d#)) OR
 					(reg_q2611 AND symb_decoder(16#20#)) OR
 					(reg_q2611 AND symb_decoder(16#09#));
reg_q2613_init <= '0' ;
	p_reg_q2613: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2613 <= reg_q2613_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2613 <= reg_q2613_init;
        else
          reg_q2613 <= reg_q2613_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q532_in <= (reg_q530 AND symb_decoder(16#2e#));
reg_q532_init <= '0' ;
	p_reg_q532: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q532 <= reg_q532_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q532 <= reg_q532_init;
        else
          reg_q532 <= reg_q532_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q534_in <= (reg_q532 AND symb_decoder(16#39#)) OR
 					(reg_q532 AND symb_decoder(16#37#)) OR
 					(reg_q532 AND symb_decoder(16#35#)) OR
 					(reg_q532 AND symb_decoder(16#33#)) OR
 					(reg_q532 AND symb_decoder(16#30#)) OR
 					(reg_q532 AND symb_decoder(16#38#)) OR
 					(reg_q532 AND symb_decoder(16#31#)) OR
 					(reg_q532 AND symb_decoder(16#32#)) OR
 					(reg_q532 AND symb_decoder(16#34#)) OR
 					(reg_q532 AND symb_decoder(16#36#)) OR
 					(reg_q534 AND symb_decoder(16#36#)) OR
 					(reg_q534 AND symb_decoder(16#38#)) OR
 					(reg_q534 AND symb_decoder(16#33#)) OR
 					(reg_q534 AND symb_decoder(16#34#)) OR
 					(reg_q534 AND symb_decoder(16#32#)) OR
 					(reg_q534 AND symb_decoder(16#35#)) OR
 					(reg_q534 AND symb_decoder(16#37#)) OR
 					(reg_q534 AND symb_decoder(16#31#)) OR
 					(reg_q534 AND symb_decoder(16#30#)) OR
 					(reg_q534 AND symb_decoder(16#39#));
reg_q534_init <= '0' ;
	p_reg_q534: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q534 <= reg_q534_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q534 <= reg_q534_init;
        else
          reg_q534 <= reg_q534_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1916_in <= (reg_q1914 AND symb_decoder(16#45#)) OR
 					(reg_q1914 AND symb_decoder(16#65#));
reg_q1916_init <= '0' ;
	p_reg_q1916: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1916 <= reg_q1916_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1916 <= reg_q1916_init;
        else
          reg_q1916 <= reg_q1916_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1498_in <= (reg_q1496 AND symb_decoder(16#56#)) OR
 					(reg_q1496 AND symb_decoder(16#76#));
reg_q1498_init <= '0' ;
	p_reg_q1498: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1498 <= reg_q1498_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1498 <= reg_q1498_init;
        else
          reg_q1498 <= reg_q1498_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1500_in <= (reg_q1498 AND symb_decoder(16#65#)) OR
 					(reg_q1498 AND symb_decoder(16#45#));
reg_q1500_init <= '0' ;
	p_reg_q1500: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1500 <= reg_q1500_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1500 <= reg_q1500_init;
        else
          reg_q1500 <= reg_q1500_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q684_in <= (reg_q682 AND symb_decoder(16#31#));
reg_q684_init <= '0' ;
	p_reg_q684: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q684 <= reg_q684_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q684 <= reg_q684_init;
        else
          reg_q684 <= reg_q684_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2506_in <= (reg_q2504 AND symb_decoder(16#4f#));
reg_q2506_init <= '0' ;
	p_reg_q2506: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2506 <= reg_q2506_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2506 <= reg_q2506_init;
        else
          reg_q2506 <= reg_q2506_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2508_in <= (reg_q2506 AND symb_decoder(16#52#));
reg_q2508_init <= '0' ;
	p_reg_q2508: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2508 <= reg_q2508_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2508 <= reg_q2508_init;
        else
          reg_q2508 <= reg_q2508_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1894_in <= (reg_q1892 AND symb_decoder(16#6f#)) OR
 					(reg_q1892 AND symb_decoder(16#4f#));
reg_q1894_init <= '0' ;
	p_reg_q1894: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1894 <= reg_q1894_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1894 <= reg_q1894_init;
        else
          reg_q1894 <= reg_q1894_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1896_in <= (reg_q1894 AND symb_decoder(16#77#)) OR
 					(reg_q1894 AND symb_decoder(16#57#));
reg_q1896_init <= '0' ;
	p_reg_q1896: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1896 <= reg_q1896_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1896 <= reg_q1896_init;
        else
          reg_q1896 <= reg_q1896_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q304_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q303 AND symb_decoder(16#0a#)) OR
 					(reg_q303 AND symb_decoder(16#0d#));
reg_q304_init <= '0' ;
	p_reg_q304: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q304 <= reg_q304_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q304 <= reg_q304_init;
        else
          reg_q304 <= reg_q304_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q462_in <= (reg_q460 AND symb_decoder(16#3d#));
reg_q462_init <= '0' ;
	p_reg_q462: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q462 <= reg_q462_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q462 <= reg_q462_init;
        else
          reg_q462 <= reg_q462_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q464_in <= (reg_q462 AND symb_decoder(16#46#)) OR
 					(reg_q462 AND symb_decoder(16#66#));
reg_q464_init <= '0' ;
	p_reg_q464: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q464 <= reg_q464_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q464 <= reg_q464_init;
        else
          reg_q464 <= reg_q464_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2646_in <= (reg_q2644 AND symb_decoder(16#52#)) OR
 					(reg_q2644 AND symb_decoder(16#72#));
reg_q2646_init <= '0' ;
	p_reg_q2646: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2646 <= reg_q2646_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2646 <= reg_q2646_init;
        else
          reg_q2646 <= reg_q2646_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2648_in <= (reg_q2646 AND symb_decoder(16#20#)) OR
 					(reg_q2646 AND symb_decoder(16#0c#)) OR
 					(reg_q2646 AND symb_decoder(16#0a#)) OR
 					(reg_q2646 AND symb_decoder(16#0d#)) OR
 					(reg_q2646 AND symb_decoder(16#09#));
reg_q2648_init <= '0' ;
	p_reg_q2648: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2648 <= reg_q2648_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2648 <= reg_q2648_init;
        else
          reg_q2648 <= reg_q2648_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1149_in <= (reg_q1147 AND symb_decoder(16#0d#));
reg_q1149_init <= '0' ;
	p_reg_q1149: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1149 <= reg_q1149_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1149 <= reg_q1149_init;
        else
          reg_q1149 <= reg_q1149_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2658_in <= (reg_q2656 AND symb_decoder(16#59#)) OR
 					(reg_q2656 AND symb_decoder(16#79#));
reg_q2658_init <= '0' ;
	p_reg_q2658: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2658 <= reg_q2658_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2658 <= reg_q2658_init;
        else
          reg_q2658 <= reg_q2658_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2660_in <= (reg_q2658 AND symb_decoder(16#4c#)) OR
 					(reg_q2658 AND symb_decoder(16#6c#));
reg_q2660_init <= '0' ;
	p_reg_q2660: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2660 <= reg_q2660_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2660 <= reg_q2660_init;
        else
          reg_q2660 <= reg_q2660_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1076_in <= (reg_q1074 AND symb_decoder(16#72#)) OR
 					(reg_q1074 AND symb_decoder(16#52#));
reg_q1076_init <= '0' ;
	p_reg_q1076: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1076 <= reg_q1076_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1076 <= reg_q1076_init;
        else
          reg_q1076 <= reg_q1076_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1078_in <= (reg_q1076 AND symb_decoder(16#56#)) OR
 					(reg_q1076 AND symb_decoder(16#76#));
reg_q1078_init <= '0' ;
	p_reg_q1078: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1078 <= reg_q1078_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1078 <= reg_q1078_init;
        else
          reg_q1078 <= reg_q1078_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q658_in <= (reg_q656 AND symb_decoder(16#25#));
reg_q658_init <= '0' ;
	p_reg_q658: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q658 <= reg_q658_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q658 <= reg_q658_init;
        else
          reg_q658 <= reg_q658_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q660_in <= (reg_q658 AND symb_decoder(16#32#));
reg_q660_init <= '0' ;
	p_reg_q660: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q660 <= reg_q660_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q660 <= reg_q660_init;
        else
          reg_q660 <= reg_q660_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q418_in <= (reg_q416 AND symb_decoder(16#4c#)) OR
 					(reg_q416 AND symb_decoder(16#6c#));
reg_q418_init <= '0' ;
	p_reg_q418: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q418 <= reg_q418_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q418 <= reg_q418_init;
        else
          reg_q418 <= reg_q418_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q420_in <= (reg_q418 AND symb_decoder(16#61#)) OR
 					(reg_q418 AND symb_decoder(16#41#));
reg_q420_init <= '0' ;
	p_reg_q420: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q420 <= reg_q420_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q420 <= reg_q420_init;
        else
          reg_q420 <= reg_q420_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1086_in <= (reg_q1086 AND symb_decoder(16#35#)) OR
 					(reg_q1086 AND symb_decoder(16#39#)) OR
 					(reg_q1086 AND symb_decoder(16#31#)) OR
 					(reg_q1086 AND symb_decoder(16#33#)) OR
 					(reg_q1086 AND symb_decoder(16#30#)) OR
 					(reg_q1086 AND symb_decoder(16#37#)) OR
 					(reg_q1086 AND symb_decoder(16#36#)) OR
 					(reg_q1086 AND symb_decoder(16#38#)) OR
 					(reg_q1086 AND symb_decoder(16#32#)) OR
 					(reg_q1086 AND symb_decoder(16#34#)) OR
 					(reg_q1084 AND symb_decoder(16#35#)) OR
 					(reg_q1084 AND symb_decoder(16#30#)) OR
 					(reg_q1084 AND symb_decoder(16#34#)) OR
 					(reg_q1084 AND symb_decoder(16#36#)) OR
 					(reg_q1084 AND symb_decoder(16#38#)) OR
 					(reg_q1084 AND symb_decoder(16#37#)) OR
 					(reg_q1084 AND symb_decoder(16#32#)) OR
 					(reg_q1084 AND symb_decoder(16#33#)) OR
 					(reg_q1084 AND symb_decoder(16#39#)) OR
 					(reg_q1084 AND symb_decoder(16#31#));
reg_q1086_init <= '0' ;
	p_reg_q1086: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1086 <= reg_q1086_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1086 <= reg_q1086_init;
        else
          reg_q1086 <= reg_q1086_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q726_in <= (reg_q724 AND symb_decoder(16#54#)) OR
 					(reg_q724 AND symb_decoder(16#74#));
reg_q726_init <= '0' ;
	p_reg_q726: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q726 <= reg_q726_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q726 <= reg_q726_init;
        else
          reg_q726 <= reg_q726_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q728_in <= (reg_q726 AND symb_decoder(16#69#)) OR
 					(reg_q726 AND symb_decoder(16#49#));
reg_q728_init <= '0' ;
	p_reg_q728: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q728 <= reg_q728_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q728 <= reg_q728_init;
        else
          reg_q728 <= reg_q728_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q795_in <= (reg_q813 AND symb_decoder(16#5e#)) OR
 					(reg_q791 AND symb_decoder(16#5e#));
reg_q795_init <= '0' ;
	p_reg_q795: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q795 <= reg_q795_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q795 <= reg_q795_init;
        else
          reg_q795 <= reg_q795_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q978_in <= (reg_q976 AND symb_decoder(16#65#)) OR
 					(reg_q976 AND symb_decoder(16#45#));
reg_q978_init <= '0' ;
	p_reg_q978: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q978 <= reg_q978_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q978 <= reg_q978_init;
        else
          reg_q978 <= reg_q978_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1778_in <= (reg_q1776 AND symb_decoder(16#0c#)) OR
 					(reg_q1776 AND symb_decoder(16#09#)) OR
 					(reg_q1776 AND symb_decoder(16#0d#)) OR
 					(reg_q1776 AND symb_decoder(16#20#)) OR
 					(reg_q1776 AND symb_decoder(16#0a#));
reg_q1778_init <= '0' ;
	p_reg_q1778: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1778 <= reg_q1778_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1778 <= reg_q1778_init;
        else
          reg_q1778 <= reg_q1778_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1780_in <= (reg_q1778 AND symb_decoder(16#0d#)) OR
 					(reg_q1778 AND symb_decoder(16#09#)) OR
 					(reg_q1778 AND symb_decoder(16#20#)) OR
 					(reg_q1778 AND symb_decoder(16#0c#)) OR
 					(reg_q1778 AND symb_decoder(16#0a#));
reg_q1780_init <= '0' ;
	p_reg_q1780: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1780 <= reg_q1780_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1780 <= reg_q1780_init;
        else
          reg_q1780 <= reg_q1780_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q47_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q46 AND symb_decoder(16#0d#)) OR
 					(reg_q46 AND symb_decoder(16#0a#));
reg_q47_init <= '0' ;
	p_reg_q47: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q47 <= reg_q47_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q47 <= reg_q47_init;
        else
          reg_q47 <= reg_q47_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q48_in <= (reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q47 AND symb_decoder(16#30#));
reg_q48_init <= '0' ;
	p_reg_q48: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q48 <= reg_q48_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q48 <= reg_q48_init;
        else
          reg_q48 <= reg_q48_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q707_in <= (reg_q705 AND symb_decoder(16#32#));
reg_q707_init <= '0' ;
	p_reg_q707: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q707 <= reg_q707_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q707 <= reg_q707_init;
        else
          reg_q707 <= reg_q707_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1199_in <= (reg_q1197 AND symb_decoder(16#74#)) OR
 					(reg_q1197 AND symb_decoder(16#54#));
reg_q1199_init <= '0' ;
	p_reg_q1199: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1199 <= reg_q1199_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1199 <= reg_q1199_init;
        else
          reg_q1199 <= reg_q1199_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1201_in <= (reg_q1199 AND symb_decoder(16#70#)) OR
 					(reg_q1199 AND symb_decoder(16#50#));
reg_q1201_init <= '0' ;
	p_reg_q1201: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1201 <= reg_q1201_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1201 <= reg_q1201_init;
        else
          reg_q1201 <= reg_q1201_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2304_in <= (reg_q2302 AND symb_decoder(16#4f#)) OR
 					(reg_q2302 AND symb_decoder(16#6f#));
reg_q2304_init <= '0' ;
	p_reg_q2304: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2304 <= reg_q2304_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2304 <= reg_q2304_init;
        else
          reg_q2304 <= reg_q2304_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2306_in <= (reg_q2304 AND symb_decoder(16#6e#)) OR
 					(reg_q2304 AND symb_decoder(16#4e#));
reg_q2306_init <= '0' ;
	p_reg_q2306: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2306 <= reg_q2306_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2306 <= reg_q2306_init;
        else
          reg_q2306 <= reg_q2306_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q448_in <= (reg_q448 AND symb_decoder(16#0c#)) OR
 					(reg_q448 AND symb_decoder(16#20#)) OR
 					(reg_q448 AND symb_decoder(16#0d#)) OR
 					(reg_q448 AND symb_decoder(16#0a#)) OR
 					(reg_q448 AND symb_decoder(16#09#)) OR
 					(reg_q446 AND symb_decoder(16#0c#)) OR
 					(reg_q446 AND symb_decoder(16#20#)) OR
 					(reg_q446 AND symb_decoder(16#0a#)) OR
 					(reg_q446 AND symb_decoder(16#09#)) OR
 					(reg_q446 AND symb_decoder(16#0d#));
reg_q448_init <= '0' ;
	p_reg_q448: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q448 <= reg_q448_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q448 <= reg_q448_init;
        else
          reg_q448 <= reg_q448_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1453_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1452 AND symb_decoder(16#0d#)) OR
 					(reg_q1452 AND symb_decoder(16#0a#));
reg_q1453_init <= '0' ;
	p_reg_q1453: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1453 <= reg_q1453_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1453 <= reg_q1453_init;
        else
          reg_q1453 <= reg_q1453_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1363_in <= (reg_q1361 AND symb_decoder(16#30#));
reg_q1363_init <= '0' ;
	p_reg_q1363: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1363 <= reg_q1363_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1363 <= reg_q1363_init;
        else
          reg_q1363 <= reg_q1363_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1365_in <= (reg_q1363 AND symb_decoder(16#32#));
reg_q1365_init <= '0' ;
	p_reg_q1365: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1365 <= reg_q1365_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1365 <= reg_q1365_init;
        else
          reg_q1365 <= reg_q1365_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1631_in <= (reg_q1629 AND symb_decoder(16#43#)) OR
 					(reg_q1629 AND symb_decoder(16#63#));
reg_q1631_init <= '0' ;
	p_reg_q1631: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1631 <= reg_q1631_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1631 <= reg_q1631_init;
        else
          reg_q1631 <= reg_q1631_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1633_in <= (reg_q1631 AND symb_decoder(16#54#)) OR
 					(reg_q1631 AND symb_decoder(16#74#));
reg_q1633_init <= '0' ;
	p_reg_q1633: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1633 <= reg_q1633_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1633 <= reg_q1633_init;
        else
          reg_q1633 <= reg_q1633_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1790_in <= (reg_q1788 AND symb_decoder(16#64#)) OR
 					(reg_q1788 AND symb_decoder(16#44#));
reg_q1790_init <= '0' ;
	p_reg_q1790: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1790 <= reg_q1790_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1790 <= reg_q1790_init;
        else
          reg_q1790 <= reg_q1790_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1792_in <= (reg_q1790 AND symb_decoder(16#69#)) OR
 					(reg_q1790 AND symb_decoder(16#49#));
reg_q1792_init <= '0' ;
	p_reg_q1792: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1792 <= reg_q1792_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1792 <= reg_q1792_init;
        else
          reg_q1792 <= reg_q1792_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q836_in <= (reg_q836 AND symb_decoder(16#33#)) OR
 					(reg_q836 AND symb_decoder(16#31#)) OR
 					(reg_q836 AND symb_decoder(16#38#)) OR
 					(reg_q836 AND symb_decoder(16#34#)) OR
 					(reg_q836 AND symb_decoder(16#35#)) OR
 					(reg_q836 AND symb_decoder(16#37#)) OR
 					(reg_q836 AND symb_decoder(16#32#)) OR
 					(reg_q836 AND symb_decoder(16#30#)) OR
 					(reg_q836 AND symb_decoder(16#39#)) OR
 					(reg_q836 AND symb_decoder(16#36#)) OR
 					(reg_q834 AND symb_decoder(16#31#)) OR
 					(reg_q834 AND symb_decoder(16#32#)) OR
 					(reg_q834 AND symb_decoder(16#38#)) OR
 					(reg_q834 AND symb_decoder(16#34#)) OR
 					(reg_q834 AND symb_decoder(16#33#)) OR
 					(reg_q834 AND symb_decoder(16#36#)) OR
 					(reg_q834 AND symb_decoder(16#30#)) OR
 					(reg_q834 AND symb_decoder(16#37#)) OR
 					(reg_q834 AND symb_decoder(16#39#)) OR
 					(reg_q834 AND symb_decoder(16#35#));
reg_q836_init <= '0' ;
	p_reg_q836: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q836 <= reg_q836_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q836 <= reg_q836_init;
        else
          reg_q836 <= reg_q836_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1539_in <= (reg_q1537 AND symb_decoder(16#2e#));
reg_q1539_init <= '0' ;
	p_reg_q1539: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1539 <= reg_q1539_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1539 <= reg_q1539_init;
        else
          reg_q1539 <= reg_q1539_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q510_in <= (reg_q508 AND symb_decoder(16#32#));
reg_q510_init <= '0' ;
	p_reg_q510: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q510 <= reg_q510_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q510 <= reg_q510_init;
        else
          reg_q510 <= reg_q510_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q512_in <= (reg_q510 AND symb_decoder(16#30#));
reg_q512_init <= '0' ;
	p_reg_q512: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q512 <= reg_q512_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q512 <= reg_q512_init;
        else
          reg_q512 <= reg_q512_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1284_in <= (reg_q1282 AND symb_decoder(16#69#)) OR
 					(reg_q1282 AND symb_decoder(16#49#));
reg_q1284_init <= '0' ;
	p_reg_q1284: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1284 <= reg_q1284_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1284 <= reg_q1284_init;
        else
          reg_q1284 <= reg_q1284_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1286_in <= (reg_q1284 AND symb_decoder(16#4e#)) OR
 					(reg_q1284 AND symb_decoder(16#6e#));
reg_q1286_init <= '0' ;
	p_reg_q1286: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1286 <= reg_q1286_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1286 <= reg_q1286_init;
        else
          reg_q1286 <= reg_q1286_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1256_in <= (reg_q1256 AND symb_decoder(16#30#)) OR
 					(reg_q1256 AND symb_decoder(16#32#)) OR
 					(reg_q1256 AND symb_decoder(16#38#)) OR
 					(reg_q1256 AND symb_decoder(16#33#)) OR
 					(reg_q1256 AND symb_decoder(16#34#)) OR
 					(reg_q1256 AND symb_decoder(16#36#)) OR
 					(reg_q1256 AND symb_decoder(16#31#)) OR
 					(reg_q1256 AND symb_decoder(16#39#)) OR
 					(reg_q1256 AND symb_decoder(16#35#)) OR
 					(reg_q1256 AND symb_decoder(16#37#)) OR
 					(reg_q1254 AND symb_decoder(16#31#)) OR
 					(reg_q1254 AND symb_decoder(16#37#)) OR
 					(reg_q1254 AND symb_decoder(16#32#)) OR
 					(reg_q1254 AND symb_decoder(16#34#)) OR
 					(reg_q1254 AND symb_decoder(16#35#)) OR
 					(reg_q1254 AND symb_decoder(16#36#)) OR
 					(reg_q1254 AND symb_decoder(16#38#)) OR
 					(reg_q1254 AND symb_decoder(16#33#)) OR
 					(reg_q1254 AND symb_decoder(16#30#)) OR
 					(reg_q1254 AND symb_decoder(16#39#));
reg_q1256_init <= '0' ;
	p_reg_q1256: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1256 <= reg_q1256_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1256 <= reg_q1256_init;
        else
          reg_q1256 <= reg_q1256_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1258_in <= (reg_q1256 AND symb_decoder(16#2c#));
reg_q1258_init <= '0' ;
	p_reg_q1258: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1258 <= reg_q1258_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1258 <= reg_q1258_init;
        else
          reg_q1258 <= reg_q1258_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q113_in <= (reg_q111 AND symb_decoder(16#70#)) OR
 					(reg_q111 AND symb_decoder(16#50#));
reg_q113_init <= '0' ;
	p_reg_q113: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q113 <= reg_q113_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q113 <= reg_q113_init;
        else
          reg_q113 <= reg_q113_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1987_in <= (reg_q1985 AND symb_decoder(16#2e#));
reg_q1987_init <= '0' ;
	p_reg_q1987: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1987 <= reg_q1987_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1987 <= reg_q1987_init;
        else
          reg_q1987 <= reg_q1987_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q298_in <= (reg_q296 AND symb_decoder(16#4d#)) OR
 					(reg_q296 AND symb_decoder(16#6d#));
reg_q298_init <= '0' ;
	p_reg_q298: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q298 <= reg_q298_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q298 <= reg_q298_init;
        else
          reg_q298 <= reg_q298_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q300_in <= (reg_q298 AND symb_decoder(16#45#)) OR
 					(reg_q298 AND symb_decoder(16#65#));
reg_q300_init <= '0' ;
	p_reg_q300: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q300 <= reg_q300_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q300 <= reg_q300_init;
        else
          reg_q300 <= reg_q300_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1025_in <= (reg_q1023 AND symb_decoder(16#52#)) OR
 					(reg_q1023 AND symb_decoder(16#72#));
reg_q1025_init <= '0' ;
	p_reg_q1025: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1025 <= reg_q1025_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1025 <= reg_q1025_init;
        else
          reg_q1025 <= reg_q1025_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1027_in <= (reg_q1025 AND symb_decoder(16#0d#)) OR
 					(reg_q1025 AND symb_decoder(16#0a#)) OR
 					(reg_q1025 AND symb_decoder(16#0c#)) OR
 					(reg_q1025 AND symb_decoder(16#09#)) OR
 					(reg_q1025 AND symb_decoder(16#20#)) OR
 					(reg_q1027 AND symb_decoder(16#20#)) OR
 					(reg_q1027 AND symb_decoder(16#09#)) OR
 					(reg_q1027 AND symb_decoder(16#0d#)) OR
 					(reg_q1027 AND symb_decoder(16#0a#)) OR
 					(reg_q1027 AND symb_decoder(16#0c#));
reg_q1027_init <= '0' ;
	p_reg_q1027: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1027 <= reg_q1027_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1027 <= reg_q1027_init;
        else
          reg_q1027 <= reg_q1027_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q179_in <= (reg_q178 AND symb_decoder(16#0d#)) OR
 					(reg_q178 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#));
reg_q179_init <= '0' ;
	p_reg_q179: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q179 <= reg_q179_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q179 <= reg_q179_init;
        else
          reg_q179 <= reg_q179_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1621_in <= (reg_q1619 AND symb_decoder(16#41#)) OR
 					(reg_q1619 AND symb_decoder(16#61#));
reg_q1621_init <= '0' ;
	p_reg_q1621: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1621 <= reg_q1621_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1621 <= reg_q1621_init;
        else
          reg_q1621 <= reg_q1621_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1623_in <= (reg_q1621 AND symb_decoder(16#4b#)) OR
 					(reg_q1621 AND symb_decoder(16#6b#));
reg_q1623_init <= '0' ;
	p_reg_q1623: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1623 <= reg_q1623_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1623 <= reg_q1623_init;
        else
          reg_q1623 <= reg_q1623_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q766_in <= (reg_q764 AND symb_decoder(16#63#)) OR
 					(reg_q764 AND symb_decoder(16#43#));
reg_q766_init <= '0' ;
	p_reg_q766: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q766 <= reg_q766_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q766 <= reg_q766_init;
        else
          reg_q766 <= reg_q766_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q768_in <= (reg_q766 AND symb_decoder(16#74#)) OR
 					(reg_q766 AND symb_decoder(16#54#));
reg_q768_init <= '0' ;
	p_reg_q768: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q768 <= reg_q768_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q768 <= reg_q768_init;
        else
          reg_q768 <= reg_q768_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1752_in <= (reg_q1750 AND symb_decoder(16#20#)) OR
 					(reg_q1750 AND symb_decoder(16#09#)) OR
 					(reg_q1750 AND symb_decoder(16#0d#)) OR
 					(reg_q1750 AND symb_decoder(16#0a#)) OR
 					(reg_q1750 AND symb_decoder(16#0c#));
reg_q1752_init <= '0' ;
	p_reg_q1752: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1752 <= reg_q1752_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1752 <= reg_q1752_init;
        else
          reg_q1752 <= reg_q1752_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1754_in <= (reg_q1752 AND symb_decoder(16#09#)) OR
 					(reg_q1752 AND symb_decoder(16#0a#)) OR
 					(reg_q1752 AND symb_decoder(16#20#)) OR
 					(reg_q1752 AND symb_decoder(16#0d#)) OR
 					(reg_q1752 AND symb_decoder(16#0c#));
reg_q1754_init <= '0' ;
	p_reg_q1754: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1754 <= reg_q1754_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1754 <= reg_q1754_init;
        else
          reg_q1754 <= reg_q1754_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1072_in <= (reg_q1070 AND symb_decoder(16#53#)) OR
 					(reg_q1070 AND symb_decoder(16#73#));
reg_q1072_init <= '0' ;
	p_reg_q1072: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1072 <= reg_q1072_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1072 <= reg_q1072_init;
        else
          reg_q1072 <= reg_q1072_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2324_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2323 AND symb_decoder(16#0a#)) OR
 					(reg_q2323 AND symb_decoder(16#0d#));
reg_q2324_init <= '0' ;
	p_reg_q2324: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2324 <= reg_q2324_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2324 <= reg_q2324_init;
        else
          reg_q2324 <= reg_q2324_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1850_in <= (reg_q1848 AND symb_decoder(16#73#)) OR
 					(reg_q1848 AND symb_decoder(16#53#));
reg_q1850_init <= '0' ;
	p_reg_q1850: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1850 <= reg_q1850_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1850 <= reg_q1850_init;
        else
          reg_q1850 <= reg_q1850_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1852_in <= (reg_q1850 AND symb_decoder(16#65#)) OR
 					(reg_q1850 AND symb_decoder(16#45#));
reg_q1852_init <= '0' ;
	p_reg_q1852: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1852 <= reg_q1852_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1852 <= reg_q1852_init;
        else
          reg_q1852 <= reg_q1852_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q137_in <= (reg_q135 AND symb_decoder(16#4e#)) OR
 					(reg_q135 AND symb_decoder(16#6e#));
reg_q137_init <= '0' ;
	p_reg_q137: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q137 <= reg_q137_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q137 <= reg_q137_init;
        else
          reg_q137 <= reg_q137_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q139_in <= (reg_q137 AND symb_decoder(16#45#)) OR
 					(reg_q137 AND symb_decoder(16#65#));
reg_q139_init <= '0' ;
	p_reg_q139: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q139 <= reg_q139_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q139 <= reg_q139_init;
        else
          reg_q139 <= reg_q139_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2278_in <= (reg_q2278 AND symb_decoder(16#09#)) OR
 					(reg_q2278 AND symb_decoder(16#20#)) OR
 					(reg_q2278 AND symb_decoder(16#0c#)) OR
 					(reg_q2278 AND symb_decoder(16#0a#)) OR
 					(reg_q2278 AND symb_decoder(16#0d#)) OR
 					(reg_q2276 AND symb_decoder(16#20#)) OR
 					(reg_q2276 AND symb_decoder(16#0a#)) OR
 					(reg_q2276 AND symb_decoder(16#0d#)) OR
 					(reg_q2276 AND symb_decoder(16#0c#)) OR
 					(reg_q2276 AND symb_decoder(16#09#));
reg_q2278_init <= '0' ;
	p_reg_q2278: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2278 <= reg_q2278_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2278 <= reg_q2278_init;
        else
          reg_q2278 <= reg_q2278_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q286_in <= (reg_q284 AND symb_decoder(16#20#));
reg_q286_init <= '0' ;
	p_reg_q286: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q286 <= reg_q286_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q286 <= reg_q286_init;
        else
          reg_q286 <= reg_q286_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q288_in <= (reg_q286 AND symb_decoder(16#57#)) OR
 					(reg_q286 AND symb_decoder(16#77#));
reg_q288_init <= '0' ;
	p_reg_q288: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q288 <= reg_q288_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q288 <= reg_q288_init;
        else
          reg_q288 <= reg_q288_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q614_in <= (reg_q612 AND symb_decoder(16#45#)) OR
 					(reg_q612 AND symb_decoder(16#65#));
reg_q614_init <= '0' ;
	p_reg_q614: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q614 <= reg_q614_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q614 <= reg_q614_init;
        else
          reg_q614 <= reg_q614_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q887_in <= (reg_q887 AND symb_decoder(16#20#)) OR
 					(reg_q887 AND symb_decoder(16#0d#)) OR
 					(reg_q887 AND symb_decoder(16#0c#)) OR
 					(reg_q887 AND symb_decoder(16#09#)) OR
 					(reg_q887 AND symb_decoder(16#0a#)) OR
 					(reg_q884 AND symb_decoder(16#20#)) OR
 					(reg_q884 AND symb_decoder(16#0c#)) OR
 					(reg_q884 AND symb_decoder(16#0d#)) OR
 					(reg_q884 AND symb_decoder(16#0a#)) OR
 					(reg_q884 AND symb_decoder(16#09#));
reg_q887_init <= '0' ;
	p_reg_q887: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q887 <= reg_q887_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q887 <= reg_q887_init;
        else
          reg_q887 <= reg_q887_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q231_in <= (reg_q229 AND symb_decoder(16#36#));
reg_q231_init <= '0' ;
	p_reg_q231: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q231 <= reg_q231_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q231 <= reg_q231_init;
        else
          reg_q231 <= reg_q231_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2429_in <= (reg_q2427 AND symb_decoder(16#43#)) OR
 					(reg_q2427 AND symb_decoder(16#63#));
reg_q2429_init <= '0' ;
	p_reg_q2429: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2429 <= reg_q2429_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2429 <= reg_q2429_init;
        else
          reg_q2429 <= reg_q2429_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2431_in <= (reg_q2429 AND symb_decoder(16#4f#)) OR
 					(reg_q2429 AND symb_decoder(16#6f#));
reg_q2431_init <= '0' ;
	p_reg_q2431: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2431 <= reg_q2431_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2431 <= reg_q2431_init;
        else
          reg_q2431 <= reg_q2431_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1545_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1544 AND symb_decoder(16#0a#)) OR
 					(reg_q1544 AND symb_decoder(16#0d#));
reg_q1545_init <= '0' ;
	p_reg_q1545: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1545 <= reg_q1545_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1545 <= reg_q1545_init;
        else
          reg_q1545 <= reg_q1545_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1546_in <= (reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q1545 AND symb_decoder(16#6e#)) OR
 					(reg_q1545 AND symb_decoder(16#4e#));
reg_q1546_init <= '0' ;
	p_reg_q1546: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1546 <= reg_q1546_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1546 <= reg_q1546_init;
        else
          reg_q1546 <= reg_q1546_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1806_in <= (reg_q1804 AND symb_decoder(16#45#)) OR
 					(reg_q1804 AND symb_decoder(16#65#));
reg_q1806_init <= '0' ;
	p_reg_q1806: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1806 <= reg_q1806_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1806 <= reg_q1806_init;
        else
          reg_q1806 <= reg_q1806_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1808_in <= (reg_q1806 AND symb_decoder(16#52#)) OR
 					(reg_q1806 AND symb_decoder(16#72#));
reg_q1808_init <= '0' ;
	p_reg_q1808: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1808 <= reg_q1808_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1808 <= reg_q1808_init;
        else
          reg_q1808 <= reg_q1808_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2202_in <= (reg_q2200 AND symb_decoder(16#6d#)) OR
 					(reg_q2200 AND symb_decoder(16#4d#));
reg_q2202_init <= '0' ;
	p_reg_q2202: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2202 <= reg_q2202_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2202 <= reg_q2202_init;
        else
          reg_q2202 <= reg_q2202_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2204_in <= (reg_q2202 AND symb_decoder(16#6f#)) OR
 					(reg_q2202 AND symb_decoder(16#4f#));
reg_q2204_init <= '0' ;
	p_reg_q2204: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2204 <= reg_q2204_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2204 <= reg_q2204_init;
        else
          reg_q2204 <= reg_q2204_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1554_in <= (reg_q1552 AND symb_decoder(16#70#)) OR
 					(reg_q1552 AND symb_decoder(16#50#));
reg_q1554_init <= '0' ;
	p_reg_q1554: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1554 <= reg_q1554_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1554 <= reg_q1554_init;
        else
          reg_q1554 <= reg_q1554_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1556_in <= (reg_q1554 AND symb_decoder(16#79#)) OR
 					(reg_q1554 AND symb_decoder(16#59#));
reg_q1556_init <= '0' ;
	p_reg_q1556: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1556 <= reg_q1556_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1556 <= reg_q1556_init;
        else
          reg_q1556 <= reg_q1556_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1882_in <= (reg_q1882 AND symb_decoder(16#34#)) OR
 					(reg_q1882 AND symb_decoder(16#39#)) OR
 					(reg_q1882 AND symb_decoder(16#32#)) OR
 					(reg_q1882 AND symb_decoder(16#33#)) OR
 					(reg_q1882 AND symb_decoder(16#38#)) OR
 					(reg_q1882 AND symb_decoder(16#30#)) OR
 					(reg_q1882 AND symb_decoder(16#37#)) OR
 					(reg_q1882 AND symb_decoder(16#31#)) OR
 					(reg_q1882 AND symb_decoder(16#35#)) OR
 					(reg_q1882 AND symb_decoder(16#36#)) OR
 					(reg_q1880 AND symb_decoder(16#31#)) OR
 					(reg_q1880 AND symb_decoder(16#32#)) OR
 					(reg_q1880 AND symb_decoder(16#35#)) OR
 					(reg_q1880 AND symb_decoder(16#36#)) OR
 					(reg_q1880 AND symb_decoder(16#30#)) OR
 					(reg_q1880 AND symb_decoder(16#39#)) OR
 					(reg_q1880 AND symb_decoder(16#34#)) OR
 					(reg_q1880 AND symb_decoder(16#37#)) OR
 					(reg_q1880 AND symb_decoder(16#33#)) OR
 					(reg_q1880 AND symb_decoder(16#38#));
reg_q1882_init <= '0' ;
	p_reg_q1882: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1882 <= reg_q1882_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1882 <= reg_q1882_init;
        else
          reg_q1882 <= reg_q1882_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1165_in <= (reg_q1163 AND symb_decoder(16#4e#)) OR
 					(reg_q1163 AND symb_decoder(16#6e#));
reg_q1165_init <= '0' ;
	p_reg_q1165: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1165 <= reg_q1165_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1165 <= reg_q1165_init;
        else
          reg_q1165 <= reg_q1165_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1167_in <= (reg_q1165 AND symb_decoder(16#6e#)) OR
 					(reg_q1165 AND symb_decoder(16#4e#));
reg_q1167_init <= '0' ;
	p_reg_q1167: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1167 <= reg_q1167_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1167 <= reg_q1167_init;
        else
          reg_q1167 <= reg_q1167_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1846_in <= (reg_q1844 AND symb_decoder(16#52#)) OR
 					(reg_q1844 AND symb_decoder(16#72#));
reg_q1846_init <= '0' ;
	p_reg_q1846: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1846 <= reg_q1846_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1846 <= reg_q1846_init;
        else
          reg_q1846 <= reg_q1846_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q884_in <= (reg_q882 AND symb_decoder(16#3a#));
reg_q884_init <= '0' ;
	p_reg_q884: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q884 <= reg_q884_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q884 <= reg_q884_init;
        else
          reg_q884 <= reg_q884_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2537_in <= (reg_q2535 AND symb_decoder(16#6e#)) OR
 					(reg_q2535 AND symb_decoder(16#4e#));
reg_q2537_init <= '0' ;
	p_reg_q2537: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2537 <= reg_q2537_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2537 <= reg_q2537_init;
        else
          reg_q2537 <= reg_q2537_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q149_in <= (reg_q149 AND symb_decoder(16#20#)) OR
 					(reg_q149 AND symb_decoder(16#0c#)) OR
 					(reg_q149 AND symb_decoder(16#09#)) OR
 					(reg_q149 AND symb_decoder(16#0d#)) OR
 					(reg_q149 AND symb_decoder(16#0a#)) OR
 					(reg_q147 AND symb_decoder(16#20#)) OR
 					(reg_q147 AND symb_decoder(16#0c#)) OR
 					(reg_q147 AND symb_decoder(16#0d#)) OR
 					(reg_q147 AND symb_decoder(16#0a#)) OR
 					(reg_q147 AND symb_decoder(16#09#));
reg_q149_init <= '0' ;
	p_reg_q149: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q149 <= reg_q149_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q149 <= reg_q149_init;
        else
          reg_q149 <= reg_q149_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q151_in <= (reg_q149 AND symb_decoder(16#53#)) OR
 					(reg_q149 AND symb_decoder(16#73#));
reg_q151_init <= '0' ;
	p_reg_q151: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q151 <= reg_q151_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q151 <= reg_q151_init;
        else
          reg_q151 <= reg_q151_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1173_in <= (reg_q1171 AND symb_decoder(16#54#)) OR
 					(reg_q1171 AND symb_decoder(16#74#));
reg_q1173_init <= '0' ;
	p_reg_q1173: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1173 <= reg_q1173_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1173 <= reg_q1173_init;
        else
          reg_q1173 <= reg_q1173_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1175_in <= (reg_q1173 AND symb_decoder(16#69#)) OR
 					(reg_q1173 AND symb_decoder(16#49#));
reg_q1175_init <= '0' ;
	p_reg_q1175: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1175 <= reg_q1175_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1175 <= reg_q1175_init;
        else
          reg_q1175 <= reg_q1175_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2351_in <= (reg_q2351 AND symb_decoder(16#20#)) OR
 					(reg_q2351 AND symb_decoder(16#0c#)) OR
 					(reg_q2351 AND symb_decoder(16#09#)) OR
 					(reg_q2351 AND symb_decoder(16#0d#)) OR
 					(reg_q2351 AND symb_decoder(16#0a#)) OR
 					(reg_q2349 AND symb_decoder(16#20#)) OR
 					(reg_q2349 AND symb_decoder(16#0d#)) OR
 					(reg_q2349 AND symb_decoder(16#09#)) OR
 					(reg_q2349 AND symb_decoder(16#0a#)) OR
 					(reg_q2349 AND symb_decoder(16#0c#));
reg_q2351_init <= '0' ;
	p_reg_q2351: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2351 <= reg_q2351_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2351 <= reg_q2351_init;
        else
          reg_q2351 <= reg_q2351_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2553_in <= (reg_q2551 AND symb_decoder(16#53#)) OR
 					(reg_q2551 AND symb_decoder(16#73#));
reg_q2553_init <= '0' ;
	p_reg_q2553: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2553 <= reg_q2553_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2553 <= reg_q2553_init;
        else
          reg_q2553 <= reg_q2553_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2555_in <= (reg_q2553 AND symb_decoder(16#74#)) OR
 					(reg_q2553 AND symb_decoder(16#54#));
reg_q2555_init <= '0' ;
	p_reg_q2555: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2555 <= reg_q2555_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2555 <= reg_q2555_init;
        else
          reg_q2555 <= reg_q2555_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q20_in <= (reg_q18 AND symb_decoder(16#53#)) OR
 					(reg_q18 AND symb_decoder(16#73#));
reg_q20_init <= '0' ;
	p_reg_q20: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q20 <= reg_q20_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q20 <= reg_q20_init;
        else
          reg_q20 <= reg_q20_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2245_in <= (reg_q2243 AND symb_decoder(16#30#)) OR
 					(reg_q2243 AND symb_decoder(16#38#)) OR
 					(reg_q2243 AND symb_decoder(16#32#)) OR
 					(reg_q2243 AND symb_decoder(16#39#)) OR
 					(reg_q2243 AND symb_decoder(16#35#)) OR
 					(reg_q2243 AND symb_decoder(16#33#)) OR
 					(reg_q2243 AND symb_decoder(16#36#)) OR
 					(reg_q2243 AND symb_decoder(16#37#)) OR
 					(reg_q2243 AND symb_decoder(16#31#)) OR
 					(reg_q2243 AND symb_decoder(16#34#)) OR
 					(reg_q2245 AND symb_decoder(16#31#)) OR
 					(reg_q2245 AND symb_decoder(16#35#)) OR
 					(reg_q2245 AND symb_decoder(16#33#)) OR
 					(reg_q2245 AND symb_decoder(16#38#)) OR
 					(reg_q2245 AND symb_decoder(16#39#)) OR
 					(reg_q2245 AND symb_decoder(16#36#)) OR
 					(reg_q2245 AND symb_decoder(16#30#)) OR
 					(reg_q2245 AND symb_decoder(16#37#)) OR
 					(reg_q2245 AND symb_decoder(16#32#)) OR
 					(reg_q2245 AND symb_decoder(16#34#));
reg_q2245_init <= '0' ;
	p_reg_q2245: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2245 <= reg_q2245_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2245 <= reg_q2245_init;
        else
          reg_q2245 <= reg_q2245_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1041_in <= (reg_q1039 AND symb_decoder(16#52#)) OR
 					(reg_q1039 AND symb_decoder(16#72#));
reg_q1041_init <= '0' ;
	p_reg_q1041: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1041 <= reg_q1041_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1041 <= reg_q1041_init;
        else
          reg_q1041 <= reg_q1041_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1043_in <= (reg_q1041 AND symb_decoder(16#76#)) OR
 					(reg_q1041 AND symb_decoder(16#56#));
reg_q1043_init <= '0' ;
	p_reg_q1043: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1043 <= reg_q1043_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1043 <= reg_q1043_init;
        else
          reg_q1043 <= reg_q1043_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1981_in <= (reg_q1981 AND symb_decoder(16#32#)) OR
 					(reg_q1981 AND symb_decoder(16#34#)) OR
 					(reg_q1981 AND symb_decoder(16#30#)) OR
 					(reg_q1981 AND symb_decoder(16#33#)) OR
 					(reg_q1981 AND symb_decoder(16#36#)) OR
 					(reg_q1981 AND symb_decoder(16#31#)) OR
 					(reg_q1981 AND symb_decoder(16#35#)) OR
 					(reg_q1981 AND symb_decoder(16#37#)) OR
 					(reg_q1981 AND symb_decoder(16#39#)) OR
 					(reg_q1981 AND symb_decoder(16#38#)) OR
 					(reg_q1979 AND symb_decoder(16#31#)) OR
 					(reg_q1979 AND symb_decoder(16#30#)) OR
 					(reg_q1979 AND symb_decoder(16#34#)) OR
 					(reg_q1979 AND symb_decoder(16#32#)) OR
 					(reg_q1979 AND symb_decoder(16#36#)) OR
 					(reg_q1979 AND symb_decoder(16#37#)) OR
 					(reg_q1979 AND symb_decoder(16#33#)) OR
 					(reg_q1979 AND symb_decoder(16#38#)) OR
 					(reg_q1979 AND symb_decoder(16#35#)) OR
 					(reg_q1979 AND symb_decoder(16#39#));
reg_q1981_init <= '0' ;
	p_reg_q1981: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1981 <= reg_q1981_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1981 <= reg_q1981_init;
        else
          reg_q1981 <= reg_q1981_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2276_in <= (reg_q2274 AND symb_decoder(16#4f#)) OR
 					(reg_q2274 AND symb_decoder(16#6f#));
reg_q2276_init <= '0' ;
	p_reg_q2276: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2276 <= reg_q2276_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2276 <= reg_q2276_init;
        else
          reg_q2276 <= reg_q2276_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1288_in <= (reg_q1286 AND symb_decoder(16#65#)) OR
 					(reg_q1286 AND symb_decoder(16#45#));
reg_q1288_init <= '0' ;
	p_reg_q1288: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1288 <= reg_q1288_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1288 <= reg_q1288_init;
        else
          reg_q1288 <= reg_q1288_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q602_in <= (reg_q600 AND symb_decoder(16#4f#)) OR
 					(reg_q600 AND symb_decoder(16#6f#));
reg_q602_init <= '0' ;
	p_reg_q602: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q602 <= reg_q602_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q602 <= reg_q602_init;
        else
          reg_q602 <= reg_q602_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q604_in <= (reg_q602 AND symb_decoder(16#0d#)) OR
 					(reg_q602 AND symb_decoder(16#0a#)) OR
 					(reg_q602 AND symb_decoder(16#20#)) OR
 					(reg_q602 AND symb_decoder(16#09#)) OR
 					(reg_q602 AND symb_decoder(16#0c#)) OR
 					(reg_q604 AND symb_decoder(16#0a#)) OR
 					(reg_q604 AND symb_decoder(16#20#)) OR
 					(reg_q604 AND symb_decoder(16#09#)) OR
 					(reg_q604 AND symb_decoder(16#0d#)) OR
 					(reg_q604 AND symb_decoder(16#0c#));
reg_q604_init <= '0' ;
	p_reg_q604: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q604 <= reg_q604_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q604 <= reg_q604_init;
        else
          reg_q604 <= reg_q604_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2034_in <= (reg_q2032 AND symb_decoder(16#69#)) OR
 					(reg_q2032 AND symb_decoder(16#49#));
reg_q2034_init <= '0' ;
	p_reg_q2034: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2034 <= reg_q2034_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2034 <= reg_q2034_init;
        else
          reg_q2034 <= reg_q2034_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1006_in <= (reg_q1004 AND symb_decoder(16#29#));
reg_q1006_init <= '0' ;
	p_reg_q1006: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1006 <= reg_q1006_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1006 <= reg_q1006_init;
        else
          reg_q1006 <= reg_q1006_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1008_in <= (reg_q1006 AND symb_decoder(16#0d#));
reg_q1008_init <= '0' ;
	p_reg_q1008: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1008 <= reg_q1008_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1008 <= reg_q1008_init;
        else
          reg_q1008 <= reg_q1008_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q266_in <= (reg_q264 AND symb_decoder(16#2d#));
reg_q266_init <= '0' ;
	p_reg_q266: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q266 <= reg_q266_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q266 <= reg_q266_init;
        else
          reg_q266 <= reg_q266_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q268_in <= (reg_q266 AND symb_decoder(16#33#));
reg_q268_init <= '0' ;
	p_reg_q268: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q268 <= reg_q268_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q268 <= reg_q268_init;
        else
          reg_q268 <= reg_q268_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2333_in <= (reg_q2331 AND symb_decoder(16#6c#)) OR
 					(reg_q2331 AND symb_decoder(16#4c#));
reg_q2333_init <= '0' ;
	p_reg_q2333: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2333 <= reg_q2333_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2333 <= reg_q2333_init;
        else
          reg_q2333 <= reg_q2333_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2335_in <= (reg_q2333 AND symb_decoder(16#66#)) OR
 					(reg_q2333 AND symb_decoder(16#46#));
reg_q2335_init <= '0' ;
	p_reg_q2335: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2335 <= reg_q2335_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2335 <= reg_q2335_init;
        else
          reg_q2335 <= reg_q2335_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1211_in <= (reg_q1209 AND symb_decoder(16#54#)) OR
 					(reg_q1209 AND symb_decoder(16#74#));
reg_q1211_init <= '0' ;
	p_reg_q1211: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1211 <= reg_q1211_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1211 <= reg_q1211_init;
        else
          reg_q1211 <= reg_q1211_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1197_in <= (reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q1195 AND symb_decoder(16#66#)) OR
 					(reg_q1195 AND symb_decoder(16#46#));
reg_q1197_init <= '0' ;
	p_reg_q1197: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1197 <= reg_q1197_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1197 <= reg_q1197_init;
        else
          reg_q1197 <= reg_q1197_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1242_in <= (reg_q1240 AND symb_decoder(16#68#)) OR
 					(reg_q1240 AND symb_decoder(16#48#));
reg_q1242_init <= '0' ;
	p_reg_q1242: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1242 <= reg_q1242_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1242 <= reg_q1242_init;
        else
          reg_q1242 <= reg_q1242_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1244_in <= (reg_q1242 AND symb_decoder(16#45#)) OR
 					(reg_q1242 AND symb_decoder(16#65#));
reg_q1244_init <= '0' ;
	p_reg_q1244: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1244 <= reg_q1244_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1244 <= reg_q1244_init;
        else
          reg_q1244 <= reg_q1244_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q198_in <= (reg_q196 AND symb_decoder(16#4e#)) OR
 					(reg_q196 AND symb_decoder(16#6e#));
reg_q198_init <= '0' ;
	p_reg_q198: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q198 <= reg_q198_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q198 <= reg_q198_init;
        else
          reg_q198 <= reg_q198_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q200_in <= (reg_q198 AND symb_decoder(16#54#)) OR
 					(reg_q198 AND symb_decoder(16#74#));
reg_q200_init <= '0' ;
	p_reg_q200: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q200 <= reg_q200_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q200 <= reg_q200_init;
        else
          reg_q200 <= reg_q200_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2487_in <= (reg_q2485 AND symb_decoder(16#50#));
reg_q2487_init <= '0' ;
	p_reg_q2487: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2487 <= reg_q2487_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2487 <= reg_q2487_init;
        else
          reg_q2487 <= reg_q2487_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2489_in <= (reg_q2487 AND symb_decoder(16#4f#));
reg_q2489_init <= '0' ;
	p_reg_q2489: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2489 <= reg_q2489_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2489 <= reg_q2489_init;
        else
          reg_q2489 <= reg_q2489_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2268_in <= (reg_q2266 AND symb_decoder(16#78#)) OR
 					(reg_q2266 AND symb_decoder(16#58#));
reg_q2268_init <= '0' ;
	p_reg_q2268: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2268 <= reg_q2268_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2268 <= reg_q2268_init;
        else
          reg_q2268 <= reg_q2268_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2270_in <= (reg_q2268 AND symb_decoder(16#0c#)) OR
 					(reg_q2268 AND symb_decoder(16#09#)) OR
 					(reg_q2268 AND symb_decoder(16#20#)) OR
 					(reg_q2268 AND symb_decoder(16#0d#)) OR
 					(reg_q2268 AND symb_decoder(16#0a#)) OR
 					(reg_q2270 AND symb_decoder(16#20#)) OR
 					(reg_q2270 AND symb_decoder(16#0c#)) OR
 					(reg_q2270 AND symb_decoder(16#0a#)) OR
 					(reg_q2270 AND symb_decoder(16#0d#)) OR
 					(reg_q2270 AND symb_decoder(16#09#));
reg_q2270_init <= '0' ;
	p_reg_q2270: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2270 <= reg_q2270_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2270 <= reg_q2270_init;
        else
          reg_q2270 <= reg_q2270_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q243_in <= (reg_q241 AND symb_decoder(16#ff#));
reg_q243_init <= '0' ;
	p_reg_q243: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q243 <= reg_q243_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q243 <= reg_q243_init;
        else
          reg_q243 <= reg_q243_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1056_in <= (reg_q1054 AND symb_decoder(16#50#)) OR
 					(reg_q1054 AND symb_decoder(16#70#));
reg_q1056_init <= '0' ;
	p_reg_q1056: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1056 <= reg_q1056_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1056 <= reg_q1056_init;
        else
          reg_q1056 <= reg_q1056_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1058_in <= (reg_q1056 AND symb_decoder(16#6c#)) OR
 					(reg_q1056 AND symb_decoder(16#4c#));
reg_q1058_init <= '0' ;
	p_reg_q1058: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1058 <= reg_q1058_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1058 <= reg_q1058_init;
        else
          reg_q1058 <= reg_q1058_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1115_in <= (reg_q1113 AND symb_decoder(16#6f#)) OR
 					(reg_q1113 AND symb_decoder(16#4f#));
reg_q1115_init <= '0' ;
	p_reg_q1115: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1115 <= reg_q1115_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1115 <= reg_q1115_init;
        else
          reg_q1115 <= reg_q1115_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1117_in <= (reg_q1115 AND symb_decoder(16#52#)) OR
 					(reg_q1115 AND symb_decoder(16#72#));
reg_q1117_init <= '0' ;
	p_reg_q1117: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1117 <= reg_q1117_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1117 <= reg_q1117_init;
        else
          reg_q1117 <= reg_q1117_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1135_in <= (reg_q1133 AND symb_decoder(16#59#)) OR
 					(reg_q1133 AND symb_decoder(16#79#));
reg_q1135_init <= '0' ;
	p_reg_q1135: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1135 <= reg_q1135_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1135 <= reg_q1135_init;
        else
          reg_q1135 <= reg_q1135_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q864_in <= (reg_q864 AND symb_decoder(16#09#)) OR
 					(reg_q864 AND symb_decoder(16#0c#)) OR
 					(reg_q864 AND symb_decoder(16#20#)) OR
 					(reg_q864 AND symb_decoder(16#0d#)) OR
 					(reg_q864 AND symb_decoder(16#0a#)) OR
 					(reg_q862 AND symb_decoder(16#0c#)) OR
 					(reg_q862 AND symb_decoder(16#0d#)) OR
 					(reg_q862 AND symb_decoder(16#20#)) OR
 					(reg_q862 AND symb_decoder(16#09#)) OR
 					(reg_q862 AND symb_decoder(16#0a#));
reg_q864_init <= '0' ;
	p_reg_q864: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q864 <= reg_q864_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q864 <= reg_q864_init;
        else
          reg_q864 <= reg_q864_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2048_in <= (reg_q2046 AND symb_decoder(16#4d#)) OR
 					(reg_q2046 AND symb_decoder(16#6d#));
reg_q2048_init <= '0' ;
	p_reg_q2048: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2048 <= reg_q2048_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2048 <= reg_q2048_init;
        else
          reg_q2048 <= reg_q2048_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2050_in <= (reg_q2048 AND symb_decoder(16#3a#));
reg_q2050_init <= '0' ;
	p_reg_q2050: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2050 <= reg_q2050_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2050 <= reg_q2050_init;
        else
          reg_q2050 <= reg_q2050_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2113_in <= (reg_q2111 AND symb_decoder(16#79#)) OR
 					(reg_q2111 AND symb_decoder(16#59#));
reg_q2113_init <= '0' ;
	p_reg_q2113: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2113 <= reg_q2113_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2113 <= reg_q2113_init;
        else
          reg_q2113 <= reg_q2113_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2115_in <= (reg_q2113 AND symb_decoder(16#61#)) OR
 					(reg_q2113 AND symb_decoder(16#41#));
reg_q2115_init <= '0' ;
	p_reg_q2115: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2115 <= reg_q2115_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2115 <= reg_q2115_init;
        else
          reg_q2115 <= reg_q2115_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2095_in <= (reg_q2093 AND symb_decoder(16#61#)) OR
 					(reg_q2093 AND symb_decoder(16#41#));
reg_q2095_init <= '0' ;
	p_reg_q2095: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2095 <= reg_q2095_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2095 <= reg_q2095_init;
        else
          reg_q2095 <= reg_q2095_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2097_in <= (reg_q2095 AND symb_decoder(16#49#)) OR
 					(reg_q2095 AND symb_decoder(16#69#));
reg_q2097_init <= '0' ;
	p_reg_q2097: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2097 <= reg_q2097_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2097 <= reg_q2097_init;
        else
          reg_q2097 <= reg_q2097_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q145_in <= (reg_q143 AND symb_decoder(16#65#)) OR
 					(reg_q143 AND symb_decoder(16#45#));
reg_q145_init <= '0' ;
	p_reg_q145: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q145 <= reg_q145_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q145 <= reg_q145_init;
        else
          reg_q145 <= reg_q145_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q147_in <= (reg_q145 AND symb_decoder(16#64#)) OR
 					(reg_q145 AND symb_decoder(16#44#));
reg_q147_init <= '0' ;
	p_reg_q147: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q147 <= reg_q147_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q147 <= reg_q147_init;
        else
          reg_q147 <= reg_q147_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q900_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q899 AND symb_decoder(16#0a#)) OR
 					(reg_q899 AND symb_decoder(16#0d#));
reg_q900_init <= '0' ;
	p_reg_q900: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q900 <= reg_q900_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q900 <= reg_q900_init;
        else
          reg_q900 <= reg_q900_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2233_in <= (reg_q2231 AND symb_decoder(16#45#)) OR
 					(reg_q2231 AND symb_decoder(16#65#));
reg_q2233_init <= '0' ;
	p_reg_q2233: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2233 <= reg_q2233_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2233 <= reg_q2233_init;
        else
          reg_q2233 <= reg_q2233_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2235_in <= (reg_q2233 AND symb_decoder(16#52#)) OR
 					(reg_q2233 AND symb_decoder(16#72#));
reg_q2235_init <= '0' ;
	p_reg_q2235: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2235 <= reg_q2235_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2235 <= reg_q2235_init;
        else
          reg_q2235 <= reg_q2235_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1104_in <= (reg_q1102 AND symb_decoder(16#54#)) OR
 					(reg_q1102 AND symb_decoder(16#74#));
reg_q1104_init <= '0' ;
	p_reg_q1104: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1104 <= reg_q1104_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1104 <= reg_q1104_init;
        else
          reg_q1104 <= reg_q1104_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1482_in <= (reg_q1482 AND symb_decoder(16#09#)) OR
 					(reg_q1482 AND symb_decoder(16#0c#)) OR
 					(reg_q1482 AND symb_decoder(16#0d#)) OR
 					(reg_q1482 AND symb_decoder(16#20#)) OR
 					(reg_q1482 AND symb_decoder(16#0a#)) OR
 					(reg_q1480 AND symb_decoder(16#09#)) OR
 					(reg_q1480 AND symb_decoder(16#20#)) OR
 					(reg_q1480 AND symb_decoder(16#0c#)) OR
 					(reg_q1480 AND symb_decoder(16#0a#)) OR
 					(reg_q1480 AND symb_decoder(16#0d#));
reg_q1482_init <= '0' ;
	p_reg_q1482: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1482 <= reg_q1482_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1482 <= reg_q1482_init;
        else
          reg_q1482 <= reg_q1482_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q715_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q714 AND symb_decoder(16#0d#)) OR
 					(reg_q714 AND symb_decoder(16#0a#));
reg_q715_init <= '0' ;
	p_reg_q715: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q715 <= reg_q715_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q715 <= reg_q715_init;
        else
          reg_q715 <= reg_q715_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q716_in <= (reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q715 AND symb_decoder(16#44#)) OR
 					(reg_q715 AND symb_decoder(16#64#));
reg_q716_init <= '0' ;
	p_reg_q716: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q716 <= reg_q716_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q716 <= reg_q716_init;
        else
          reg_q716 <= reg_q716_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q514_in <= (reg_q512 AND symb_decoder(16#5b#));
reg_q514_init <= '0' ;
	p_reg_q514: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q514 <= reg_q514_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q514 <= reg_q514_init;
        else
          reg_q514 <= reg_q514_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q516_in <= (reg_q514 AND symb_decoder(16#69#)) OR
 					(reg_q514 AND symb_decoder(16#49#));
reg_q516_init <= '0' ;
	p_reg_q516: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q516 <= reg_q516_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q516 <= reg_q516_init;
        else
          reg_q516 <= reg_q516_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q24_in <= (reg_q22 AND symb_decoder(16#65#)) OR
 					(reg_q22 AND symb_decoder(16#45#));
reg_q24_init <= '0' ;
	p_reg_q24: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q24 <= reg_q24_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q24 <= reg_q24_init;
        else
          reg_q24 <= reg_q24_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q26_in <= (reg_q24 AND symb_decoder(16#58#)) OR
 					(reg_q24 AND symb_decoder(16#78#));
reg_q26_init <= '0' ;
	p_reg_q26: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q26 <= reg_q26_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q26 <= reg_q26_init;
        else
          reg_q26 <= reg_q26_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q454_in <= (reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q452 AND symb_decoder(16#42#)) OR
 					(reg_q452 AND symb_decoder(16#62#));
reg_q454_init <= '0' ;
	p_reg_q454: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q454 <= reg_q454_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q454 <= reg_q454_init;
        else
          reg_q454 <= reg_q454_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q752_in <= (reg_q750 AND symb_decoder(16#6f#)) OR
 					(reg_q750 AND symb_decoder(16#4f#));
reg_q752_init <= '0' ;
	p_reg_q752: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q752 <= reg_q752_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q752 <= reg_q752_init;
        else
          reg_q752 <= reg_q752_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q754_in <= (reg_q752 AND symb_decoder(16#46#)) OR
 					(reg_q752 AND symb_decoder(16#66#));
reg_q754_init <= '0' ;
	p_reg_q754: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q754 <= reg_q754_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q754 <= reg_q754_init;
        else
          reg_q754 <= reg_q754_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1720_in <= (reg_q1720 AND symb_decoder(16#20#)) OR
 					(reg_q1720 AND symb_decoder(16#0a#)) OR
 					(reg_q1720 AND symb_decoder(16#09#)) OR
 					(reg_q1720 AND symb_decoder(16#0d#)) OR
 					(reg_q1720 AND symb_decoder(16#0c#)) OR
 					(reg_q1718 AND symb_decoder(16#20#)) OR
 					(reg_q1718 AND symb_decoder(16#09#)) OR
 					(reg_q1718 AND symb_decoder(16#0d#)) OR
 					(reg_q1718 AND symb_decoder(16#0c#)) OR
 					(reg_q1718 AND symb_decoder(16#0a#));
reg_q1720_init <= '0' ;
	p_reg_q1720: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1720 <= reg_q1720_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1720 <= reg_q1720_init;
        else
          reg_q1720 <= reg_q1720_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1886_in <= (reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q1884 AND symb_decoder(16#53#)) OR
 					(reg_q1884 AND symb_decoder(16#73#));
reg_q1886_init <= '0' ;
	p_reg_q1886: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1886 <= reg_q1886_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1886 <= reg_q1886_init;
        else
          reg_q1886 <= reg_q1886_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2164_in <= (reg_q2162 AND symb_decoder(16#61#)) OR
 					(reg_q2162 AND symb_decoder(16#41#));
reg_q2164_init <= '0' ;
	p_reg_q2164: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2164 <= reg_q2164_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2164 <= reg_q2164_init;
        else
          reg_q2164 <= reg_q2164_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2166_in <= (reg_q2164 AND symb_decoder(16#45#)) OR
 					(reg_q2164 AND symb_decoder(16#65#));
reg_q2166_init <= '0' ;
	p_reg_q2166: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2166 <= reg_q2166_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2166 <= reg_q2166_init;
        else
          reg_q2166 <= reg_q2166_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1435_in <= (reg_q1433 AND symb_decoder(16#67#)) OR
 					(reg_q1433 AND symb_decoder(16#47#));
reg_q1435_init <= '0' ;
	p_reg_q1435: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1435 <= reg_q1435_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1435 <= reg_q1435_init;
        else
          reg_q1435 <= reg_q1435_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1437_in <= (reg_q1435 AND symb_decoder(16#0a#)) OR
 					(reg_q1435 AND symb_decoder(16#09#)) OR
 					(reg_q1435 AND symb_decoder(16#0c#)) OR
 					(reg_q1435 AND symb_decoder(16#20#)) OR
 					(reg_q1435 AND symb_decoder(16#0d#)) OR
 					(reg_q1437 AND symb_decoder(16#0d#)) OR
 					(reg_q1437 AND symb_decoder(16#0a#)) OR
 					(reg_q1437 AND symb_decoder(16#20#)) OR
 					(reg_q1437 AND symb_decoder(16#0c#)) OR
 					(reg_q1437 AND symb_decoder(16#09#));
reg_q1437_init <= '0' ;
	p_reg_q1437: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1437 <= reg_q1437_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1437 <= reg_q1437_init;
        else
          reg_q1437 <= reg_q1437_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1810_in <= (reg_q1808 AND symb_decoder(16#76#)) OR
 					(reg_q1808 AND symb_decoder(16#56#));
reg_q1810_init <= '0' ;
	p_reg_q1810: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1810 <= reg_q1810_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1810 <= reg_q1810_init;
        else
          reg_q1810 <= reg_q1810_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1254_in <= (reg_q1252 AND symb_decoder(16#2e#));
reg_q1254_init <= '0' ;
	p_reg_q1254: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1254 <= reg_q1254_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1254 <= reg_q1254_init;
        else
          reg_q1254 <= reg_q1254_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1652_in <= (reg_q1650 AND symb_decoder(16#0d#)) OR
 					(reg_q1650 AND symb_decoder(16#0c#)) OR
 					(reg_q1650 AND symb_decoder(16#20#)) OR
 					(reg_q1650 AND symb_decoder(16#09#)) OR
 					(reg_q1650 AND symb_decoder(16#0a#)) OR
 					(reg_q1652 AND symb_decoder(16#0a#)) OR
 					(reg_q1652 AND symb_decoder(16#0c#)) OR
 					(reg_q1652 AND symb_decoder(16#0d#)) OR
 					(reg_q1652 AND symb_decoder(16#20#)) OR
 					(reg_q1652 AND symb_decoder(16#09#));
reg_q1652_init <= '0' ;
	p_reg_q1652: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1652 <= reg_q1652_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1652 <= reg_q1652_init;
        else
          reg_q1652 <= reg_q1652_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1654_in <= (reg_q1652 AND symb_decoder(16#36#));
reg_q1654_init <= '0' ;
	p_reg_q1654: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1654 <= reg_q1654_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1654 <= reg_q1654_init;
        else
          reg_q1654 <= reg_q1654_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1327_in <= (reg_q1325 AND symb_decoder(16#76#)) OR
 					(reg_q1325 AND symb_decoder(16#56#));
reg_q1327_init <= '0' ;
	p_reg_q1327: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1327 <= reg_q1327_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1327 <= reg_q1327_init;
        else
          reg_q1327 <= reg_q1327_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1329_in <= (reg_q1327 AND symb_decoder(16#45#)) OR
 					(reg_q1327 AND symb_decoder(16#65#));
reg_q1329_init <= '0' ;
	p_reg_q1329: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1329 <= reg_q1329_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1329 <= reg_q1329_init;
        else
          reg_q1329 <= reg_q1329_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2070_in <= (reg_q2068 AND symb_decoder(16#54#));
reg_q2070_init <= '0' ;
	p_reg_q2070: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2070 <= reg_q2070_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2070 <= reg_q2070_init;
        else
          reg_q2070 <= reg_q2070_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1125_in <= (reg_q1125 AND symb_decoder(16#0c#)) OR
 					(reg_q1125 AND symb_decoder(16#0d#)) OR
 					(reg_q1125 AND symb_decoder(16#09#)) OR
 					(reg_q1125 AND symb_decoder(16#0a#)) OR
 					(reg_q1125 AND symb_decoder(16#20#)) OR
 					(reg_q1123 AND symb_decoder(16#09#)) OR
 					(reg_q1123 AND symb_decoder(16#0d#)) OR
 					(reg_q1123 AND symb_decoder(16#0c#)) OR
 					(reg_q1123 AND symb_decoder(16#0a#)) OR
 					(reg_q1123 AND symb_decoder(16#20#));
reg_q1125_init <= '0' ;
	p_reg_q1125: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1125 <= reg_q1125_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1125 <= reg_q1125_init;
        else
          reg_q1125 <= reg_q1125_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2409_in <= (reg_q2407 AND symb_decoder(16#52#)) OR
 					(reg_q2407 AND symb_decoder(16#72#));
reg_q2409_init <= '0' ;
	p_reg_q2409: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2409 <= reg_q2409_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2409 <= reg_q2409_init;
        else
          reg_q2409 <= reg_q2409_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q986_in <= (reg_q986 AND symb_decoder(16#0c#)) OR
 					(reg_q986 AND symb_decoder(16#0d#)) OR
 					(reg_q986 AND symb_decoder(16#09#)) OR
 					(reg_q986 AND symb_decoder(16#20#)) OR
 					(reg_q986 AND symb_decoder(16#0a#)) OR
 					(reg_q984 AND symb_decoder(16#0c#)) OR
 					(reg_q984 AND symb_decoder(16#0d#)) OR
 					(reg_q984 AND symb_decoder(16#0a#)) OR
 					(reg_q984 AND symb_decoder(16#09#)) OR
 					(reg_q984 AND symb_decoder(16#20#));
reg_q986_init <= '0' ;
	p_reg_q986: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q986 <= reg_q986_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q986 <= reg_q986_init;
        else
          reg_q986 <= reg_q986_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1794_in <= (reg_q1792 AND symb_decoder(16#6d#)) OR
 					(reg_q1792 AND symb_decoder(16#4d#));
reg_q1794_init <= '0' ;
	p_reg_q1794: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1794 <= reg_q1794_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1794 <= reg_q1794_init;
        else
          reg_q1794 <= reg_q1794_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1796_in <= (reg_q1794 AND symb_decoder(16#62#)) OR
 					(reg_q1794 AND symb_decoder(16#42#));
reg_q1796_init <= '0' ;
	p_reg_q1796: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1796 <= reg_q1796_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1796 <= reg_q1796_init;
        else
          reg_q1796 <= reg_q1796_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q385_in <= (reg_q383 AND symb_decoder(16#6e#)) OR
 					(reg_q383 AND symb_decoder(16#4e#));
reg_q385_init <= '0' ;
	p_reg_q385: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q385 <= reg_q385_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q385 <= reg_q385_init;
        else
          reg_q385 <= reg_q385_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q387_in <= (reg_q385 AND symb_decoder(16#73#)) OR
 					(reg_q385 AND symb_decoder(16#53#));
reg_q387_init <= '0' ;
	p_reg_q387: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q387 <= reg_q387_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q387 <= reg_q387_init;
        else
          reg_q387 <= reg_q387_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1490_in <= (reg_q1490 AND symb_decoder(16#0d#)) OR
 					(reg_q1490 AND symb_decoder(16#09#)) OR
 					(reg_q1490 AND symb_decoder(16#20#)) OR
 					(reg_q1490 AND symb_decoder(16#0a#)) OR
 					(reg_q1490 AND symb_decoder(16#0c#)) OR
 					(reg_q1488 AND symb_decoder(16#20#)) OR
 					(reg_q1488 AND symb_decoder(16#09#)) OR
 					(reg_q1488 AND symb_decoder(16#0a#)) OR
 					(reg_q1488 AND symb_decoder(16#0d#)) OR
 					(reg_q1488 AND symb_decoder(16#0c#));
reg_q1490_init <= '0' ;
	p_reg_q1490: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1490 <= reg_q1490_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1490 <= reg_q1490_init;
        else
          reg_q1490 <= reg_q1490_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1922_in <= (reg_q1920 AND symb_decoder(16#65#)) OR
 					(reg_q1920 AND symb_decoder(16#45#));
reg_q1922_init <= '0' ;
	p_reg_q1922: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1922 <= reg_q1922_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1922 <= reg_q1922_init;
        else
          reg_q1922 <= reg_q1922_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1924_in <= (reg_q1922 AND symb_decoder(16#42#)) OR
 					(reg_q1922 AND symb_decoder(16#62#));
reg_q1924_init <= '0' ;
	p_reg_q1924: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1924 <= reg_q1924_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1924 <= reg_q1924_init;
        else
          reg_q1924 <= reg_q1924_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q862_in <= (reg_q860 AND symb_decoder(16#65#)) OR
 					(reg_q860 AND symb_decoder(16#45#));
reg_q862_init <= '0' ;
	p_reg_q862: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q862 <= reg_q862_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q862 <= reg_q862_init;
        else
          reg_q862 <= reg_q862_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2258_in <= (reg_q2256 AND symb_decoder(16#21#));
reg_q2258_init <= '0' ;
	p_reg_q2258: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2258 <= reg_q2258_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2258 <= reg_q2258_init;
        else
          reg_q2258 <= reg_q2258_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1433_in <= (reg_q1431 AND symb_decoder(16#4e#)) OR
 					(reg_q1431 AND symb_decoder(16#6e#));
reg_q1433_init <= '0' ;
	p_reg_q1433: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1433 <= reg_q1433_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1433 <= reg_q1433_init;
        else
          reg_q1433 <= reg_q1433_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1920_in <= (reg_q1918 AND symb_decoder(16#77#)) OR
 					(reg_q1918 AND symb_decoder(16#57#));
reg_q1920_init <= '0' ;
	p_reg_q1920: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1920 <= reg_q1920_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1920 <= reg_q1920_init;
        else
          reg_q1920 <= reg_q1920_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2341_in <= (reg_q2339 AND symb_decoder(16#65#)) OR
 					(reg_q2339 AND symb_decoder(16#45#));
reg_q2341_init <= '0' ;
	p_reg_q2341: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2341 <= reg_q2341_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2341 <= reg_q2341_init;
        else
          reg_q2341 <= reg_q2341_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2343_in <= (reg_q2341 AND symb_decoder(16#6d#)) OR
 					(reg_q2341 AND symb_decoder(16#4d#));
reg_q2343_init <= '0' ;
	p_reg_q2343: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2343 <= reg_q2343_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2343 <= reg_q2343_init;
        else
          reg_q2343 <= reg_q2343_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1309_in <= (reg_q1307 AND symb_decoder(16#52#)) OR
 					(reg_q1307 AND symb_decoder(16#72#));
reg_q1309_init <= '0' ;
	p_reg_q1309: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1309 <= reg_q1309_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1309 <= reg_q1309_init;
        else
          reg_q1309 <= reg_q1309_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1311_in <= (reg_q1309 AND symb_decoder(16#49#)) OR
 					(reg_q1309 AND symb_decoder(16#69#));
reg_q1311_init <= '0' ;
	p_reg_q1311: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1311 <= reg_q1311_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1311 <= reg_q1311_init;
        else
          reg_q1311 <= reg_q1311_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2286_in <= (reg_q2286 AND symb_decoder(16#33#)) OR
 					(reg_q2286 AND symb_decoder(16#37#)) OR
 					(reg_q2286 AND symb_decoder(16#35#)) OR
 					(reg_q2286 AND symb_decoder(16#38#)) OR
 					(reg_q2286 AND symb_decoder(16#31#)) OR
 					(reg_q2286 AND symb_decoder(16#32#)) OR
 					(reg_q2286 AND symb_decoder(16#30#)) OR
 					(reg_q2286 AND symb_decoder(16#39#)) OR
 					(reg_q2286 AND symb_decoder(16#36#)) OR
 					(reg_q2286 AND symb_decoder(16#34#)) OR
 					(reg_q2284 AND symb_decoder(16#38#)) OR
 					(reg_q2284 AND symb_decoder(16#39#)) OR
 					(reg_q2284 AND symb_decoder(16#32#)) OR
 					(reg_q2284 AND symb_decoder(16#37#)) OR
 					(reg_q2284 AND symb_decoder(16#31#)) OR
 					(reg_q2284 AND symb_decoder(16#36#)) OR
 					(reg_q2284 AND symb_decoder(16#33#)) OR
 					(reg_q2284 AND symb_decoder(16#30#)) OR
 					(reg_q2284 AND symb_decoder(16#34#)) OR
 					(reg_q2284 AND symb_decoder(16#35#));
reg_q2286_init <= '0' ;
	p_reg_q2286: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2286 <= reg_q2286_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2286 <= reg_q2286_init;
        else
          reg_q2286 <= reg_q2286_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q325_in <= (reg_q323 AND symb_decoder(16#00#));
reg_q325_init <= '0' ;
	p_reg_q325: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q325 <= reg_q325_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q325 <= reg_q325_init;
        else
          reg_q325 <= reg_q325_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q327_in <= (reg_q325 AND symb_decoder(16#00#));
reg_q327_init <= '0' ;
	p_reg_q327: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q327 <= reg_q327_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q327 <= reg_q327_init;
        else
          reg_q327 <= reg_q327_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2247_in <= (reg_q2245 AND symb_decoder(16#2e#));
reg_q2247_init <= '0' ;
	p_reg_q2247: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2247 <= reg_q2247_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2247 <= reg_q2247_init;
        else
          reg_q2247 <= reg_q2247_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1193_in <= (reg_q1191 AND symb_decoder(16#65#)) OR
 					(reg_q1191 AND symb_decoder(16#45#));
reg_q1193_init <= '0' ;
	p_reg_q1193: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1193 <= reg_q1193_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1193 <= reg_q1193_init;
        else
          reg_q1193 <= reg_q1193_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q450_in <= (reg_q448 AND symb_decoder(16#35#)) OR
 					(reg_q448 AND symb_decoder(16#33#)) OR
 					(reg_q448 AND symb_decoder(16#37#)) OR
 					(reg_q448 AND symb_decoder(16#31#)) OR
 					(reg_q448 AND symb_decoder(16#32#)) OR
 					(reg_q448 AND symb_decoder(16#39#)) OR
 					(reg_q448 AND symb_decoder(16#38#)) OR
 					(reg_q448 AND symb_decoder(16#34#)) OR
 					(reg_q448 AND symb_decoder(16#30#)) OR
 					(reg_q448 AND symb_decoder(16#36#)) OR
 					(reg_q450 AND symb_decoder(16#36#)) OR
 					(reg_q450 AND symb_decoder(16#30#)) OR
 					(reg_q450 AND symb_decoder(16#35#)) OR
 					(reg_q450 AND symb_decoder(16#38#)) OR
 					(reg_q450 AND symb_decoder(16#39#)) OR
 					(reg_q450 AND symb_decoder(16#32#)) OR
 					(reg_q450 AND symb_decoder(16#31#)) OR
 					(reg_q450 AND symb_decoder(16#37#)) OR
 					(reg_q450 AND symb_decoder(16#34#)) OR
 					(reg_q450 AND symb_decoder(16#33#));
reg_q450_init <= '0' ;
	p_reg_q450: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q450 <= reg_q450_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q450 <= reg_q450_init;
        else
          reg_q450 <= reg_q450_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q911_in <= (reg_q909 AND symb_decoder(16#53#)) OR
 					(reg_q909 AND symb_decoder(16#73#));
reg_q911_init <= '0' ;
	p_reg_q911: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q911 <= reg_q911_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q911 <= reg_q911_init;
        else
          reg_q911 <= reg_q911_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q980_in <= (reg_q978 AND symb_decoder(16#20#)) OR
 					(reg_q978 AND symb_decoder(16#0a#)) OR
 					(reg_q978 AND symb_decoder(16#0d#)) OR
 					(reg_q978 AND symb_decoder(16#0c#)) OR
 					(reg_q978 AND symb_decoder(16#09#)) OR
 					(reg_q980 AND symb_decoder(16#09#)) OR
 					(reg_q980 AND symb_decoder(16#20#)) OR
 					(reg_q980 AND symb_decoder(16#0d#)) OR
 					(reg_q980 AND symb_decoder(16#0a#)) OR
 					(reg_q980 AND symb_decoder(16#0c#));
reg_q980_init <= '0' ;
	p_reg_q980: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q980 <= reg_q980_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q980 <= reg_q980_init;
        else
          reg_q980 <= reg_q980_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1268_in <= (reg_q1266 AND symb_decoder(16#76#)) OR
 					(reg_q1266 AND symb_decoder(16#56#));
reg_q1268_init <= '0' ;
	p_reg_q1268: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1268 <= reg_q1268_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1268 <= reg_q1268_init;
        else
          reg_q1268 <= reg_q1268_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1270_in <= (reg_q1268 AND symb_decoder(16#65#)) OR
 					(reg_q1268 AND symb_decoder(16#45#));
reg_q1270_init <= '0' ;
	p_reg_q1270: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1270 <= reg_q1270_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1270 <= reg_q1270_init;
        else
          reg_q1270 <= reg_q1270_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q305_in <= (reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q304 AND symb_decoder(16#61#)) OR
 					(reg_q304 AND symb_decoder(16#41#));
reg_q305_init <= '0' ;
	p_reg_q305: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q305 <= reg_q305_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q305 <= reg_q305_init;
        else
          reg_q305 <= reg_q305_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q988_in <= (reg_q986 AND symb_decoder(16#65#)) OR
 					(reg_q986 AND symb_decoder(16#45#));
reg_q988_init <= '0' ;
	p_reg_q988: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q988 <= reg_q988_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q988 <= reg_q988_init;
        else
          reg_q988 <= reg_q988_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q990_in <= (reg_q988 AND symb_decoder(16#76#)) OR
 					(reg_q988 AND symb_decoder(16#56#));
reg_q990_init <= '0' ;
	p_reg_q990: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q990 <= reg_q990_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q990 <= reg_q990_init;
        else
          reg_q990 <= reg_q990_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1750_in <= (reg_q1748 AND symb_decoder(16#0d#)) OR
 					(reg_q1748 AND symb_decoder(16#20#)) OR
 					(reg_q1748 AND symb_decoder(16#0c#)) OR
 					(reg_q1748 AND symb_decoder(16#0a#)) OR
 					(reg_q1748 AND symb_decoder(16#09#));
reg_q1750_init <= '0' ;
	p_reg_q1750: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1750 <= reg_q1750_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1750 <= reg_q1750_init;
        else
          reg_q1750 <= reg_q1750_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1419_in <= (reg_q1417 AND symb_decoder(16#4f#)) OR
 					(reg_q1417 AND symb_decoder(16#6f#));
reg_q1419_init <= '0' ;
	p_reg_q1419: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1419 <= reg_q1419_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1419 <= reg_q1419_init;
        else
          reg_q1419 <= reg_q1419_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1854_in <= (reg_q1852 AND symb_decoder(16#72#)) OR
 					(reg_q1852 AND symb_decoder(16#52#));
reg_q1854_init <= '0' ;
	p_reg_q1854: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1854 <= reg_q1854_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1854 <= reg_q1854_init;
        else
          reg_q1854 <= reg_q1854_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q88_in <= (reg_q86 AND symb_decoder(16#3f#));
reg_q88_init <= '0' ;
	p_reg_q88: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q88 <= reg_q88_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q88 <= reg_q88_init;
        else
          reg_q88 <= reg_q88_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1800_in <= (reg_q1798 AND symb_decoder(16#53#)) OR
 					(reg_q1798 AND symb_decoder(16#73#));
reg_q1800_init <= '0' ;
	p_reg_q1800: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1800 <= reg_q1800_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1800 <= reg_q1800_init;
        else
          reg_q1800 <= reg_q1800_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1802_in <= (reg_q1800 AND symb_decoder(16#20#)) OR
 					(reg_q1800 AND symb_decoder(16#0a#)) OR
 					(reg_q1800 AND symb_decoder(16#09#)) OR
 					(reg_q1800 AND symb_decoder(16#0c#)) OR
 					(reg_q1800 AND symb_decoder(16#0d#)) OR
 					(reg_q1802 AND symb_decoder(16#09#)) OR
 					(reg_q1802 AND symb_decoder(16#0a#)) OR
 					(reg_q1802 AND symb_decoder(16#20#)) OR
 					(reg_q1802 AND symb_decoder(16#0c#)) OR
 					(reg_q1802 AND symb_decoder(16#0d#));
reg_q1802_init <= '0' ;
	p_reg_q1802: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1802 <= reg_q1802_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1802 <= reg_q1802_init;
        else
          reg_q1802 <= reg_q1802_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2002_in <= (reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2001 AND symb_decoder(16#54#)) OR
 					(reg_q2001 AND symb_decoder(16#74#));
reg_q2002_init <= '0' ;
	p_reg_q2002: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2002 <= reg_q2002_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2002 <= reg_q2002_init;
        else
          reg_q2002 <= reg_q2002_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2296_in <= (reg_q2294 AND symb_decoder(16#76#)) OR
 					(reg_q2294 AND symb_decoder(16#56#));
reg_q2296_init <= '0' ;
	p_reg_q2296: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2296 <= reg_q2296_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2296 <= reg_q2296_init;
        else
          reg_q2296 <= reg_q2296_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2298_in <= (reg_q2296 AND symb_decoder(16#65#)) OR
 					(reg_q2296 AND symb_decoder(16#45#));
reg_q2298_init <= '0' ;
	p_reg_q2298: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2298 <= reg_q2298_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2298 <= reg_q2298_init;
        else
          reg_q2298 <= reg_q2298_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q966_in <= (reg_q964 AND symb_decoder(16#57#)) OR
 					(reg_q964 AND symb_decoder(16#77#));
reg_q966_init <= '0' ;
	p_reg_q966: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q966 <= reg_q966_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q966 <= reg_q966_init;
        else
          reg_q966 <= reg_q966_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2652_in <= (reg_q2650 AND symb_decoder(16#0a#)) OR
 					(reg_q2650 AND symb_decoder(16#09#)) OR
 					(reg_q2650 AND symb_decoder(16#0c#)) OR
 					(reg_q2650 AND symb_decoder(16#0d#)) OR
 					(reg_q2650 AND symb_decoder(16#20#));
reg_q2652_init <= '0' ;
	p_reg_q2652: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2652 <= reg_q2652_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2652 <= reg_q2652_init;
        else
          reg_q2652 <= reg_q2652_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2654_in <= (reg_q2652 AND symb_decoder(16#6b#)) OR
 					(reg_q2652 AND symb_decoder(16#4b#));
reg_q2654_init <= '0' ;
	p_reg_q2654: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2654 <= reg_q2654_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2654 <= reg_q2654_init;
        else
          reg_q2654 <= reg_q2654_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1938_in <= (reg_q1938 AND symb_decoder(16#20#)) OR
 					(reg_q1938 AND symb_decoder(16#09#)) OR
 					(reg_q1938 AND symb_decoder(16#0a#)) OR
 					(reg_q1938 AND symb_decoder(16#0c#)) OR
 					(reg_q1938 AND symb_decoder(16#0d#)) OR
 					(reg_q1936 AND symb_decoder(16#0a#)) OR
 					(reg_q1936 AND symb_decoder(16#0d#)) OR
 					(reg_q1936 AND symb_decoder(16#0c#)) OR
 					(reg_q1936 AND symb_decoder(16#09#)) OR
 					(reg_q1936 AND symb_decoder(16#20#));
reg_q1938_init <= '0' ;
	p_reg_q1938: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1938 <= reg_q1938_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1938 <= reg_q1938_init;
        else
          reg_q1938 <= reg_q1938_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1102_in <= (reg_q1100 AND symb_decoder(16#52#)) OR
 					(reg_q1100 AND symb_decoder(16#72#));
reg_q1102_init <= '0' ;
	p_reg_q1102: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1102 <= reg_q1102_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1102 <= reg_q1102_init;
        else
          reg_q1102 <= reg_q1102_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1766_in <= (reg_q1764 AND symb_decoder(16#09#)) OR
 					(reg_q1764 AND symb_decoder(16#0c#)) OR
 					(reg_q1764 AND symb_decoder(16#0d#)) OR
 					(reg_q1764 AND symb_decoder(16#0a#)) OR
 					(reg_q1764 AND symb_decoder(16#20#));
reg_q1766_init <= '0' ;
	p_reg_q1766: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1766 <= reg_q1766_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1766 <= reg_q1766_init;
        else
          reg_q1766 <= reg_q1766_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1407_in <= (reg_q1405 AND symb_decoder(16#70#)) OR
 					(reg_q1405 AND symb_decoder(16#50#));
reg_q1407_init <= '0' ;
	p_reg_q1407: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1407 <= reg_q1407_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1407 <= reg_q1407_init;
        else
          reg_q1407 <= reg_q1407_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1409_in <= (reg_q1407 AND symb_decoder(16#41#)) OR
 					(reg_q1407 AND symb_decoder(16#61#));
reg_q1409_init <= '0' ;
	p_reg_q1409: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1409 <= reg_q1409_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1409 <= reg_q1409_init;
        else
          reg_q1409 <= reg_q1409_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q235_in <= (reg_q233 AND symb_decoder(16#ff#));
reg_q235_init <= '0' ;
	p_reg_q235: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q235 <= reg_q235_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q235 <= reg_q235_init;
        else
          reg_q235 <= reg_q235_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1381_in <= (reg_q1379 AND symb_decoder(16#65#)) OR
 					(reg_q1379 AND symb_decoder(16#45#));
reg_q1381_init <= '0' ;
	p_reg_q1381: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1381 <= reg_q1381_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1381 <= reg_q1381_init;
        else
          reg_q1381 <= reg_q1381_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1383_in <= (reg_q1381 AND symb_decoder(16#0c#)) OR
 					(reg_q1381 AND symb_decoder(16#0a#)) OR
 					(reg_q1381 AND symb_decoder(16#09#)) OR
 					(reg_q1381 AND symb_decoder(16#0d#)) OR
 					(reg_q1381 AND symb_decoder(16#20#)) OR
 					(reg_q1383 AND symb_decoder(16#20#)) OR
 					(reg_q1383 AND symb_decoder(16#0d#)) OR
 					(reg_q1383 AND symb_decoder(16#0c#)) OR
 					(reg_q1383 AND symb_decoder(16#09#)) OR
 					(reg_q1383 AND symb_decoder(16#0a#));
reg_q1383_init <= '0' ;
	p_reg_q1383: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1383 <= reg_q1383_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1383 <= reg_q1383_init;
        else
          reg_q1383 <= reg_q1383_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2642_in <= (reg_q2640 AND symb_decoder(16#76#)) OR
 					(reg_q2640 AND symb_decoder(16#56#));
reg_q2642_init <= '0' ;
	p_reg_q2642: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2642 <= reg_q2642_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2642 <= reg_q2642_init;
        else
          reg_q2642 <= reg_q2642_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2644_in <= (reg_q2642 AND symb_decoder(16#65#)) OR
 					(reg_q2642 AND symb_decoder(16#45#));
reg_q2644_init <= '0' ;
	p_reg_q2644: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2644 <= reg_q2644_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2644 <= reg_q2644_init;
        else
          reg_q2644 <= reg_q2644_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q740_in <= (reg_q738 AND symb_decoder(16#6e#)) OR
 					(reg_q738 AND symb_decoder(16#4e#));
reg_q740_init <= '0' ;
	p_reg_q740: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q740 <= reg_q740_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q740 <= reg_q740_init;
        else
          reg_q740 <= reg_q740_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1369_in <= (reg_q1367 AND symb_decoder(16#58#)) OR
 					(reg_q1367 AND symb_decoder(16#78#));
reg_q1369_init <= '0' ;
	p_reg_q1369: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1369 <= reg_q1369_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1369 <= reg_q1369_init;
        else
          reg_q1369 <= reg_q1369_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2399_in <= (reg_q2397 AND symb_decoder(16#50#)) OR
 					(reg_q2397 AND symb_decoder(16#70#));
reg_q2399_init <= '0' ;
	p_reg_q2399: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2399 <= reg_q2399_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2399 <= reg_q2399_init;
        else
          reg_q2399 <= reg_q2399_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2401_in <= (reg_q2399 AND symb_decoder(16#72#)) OR
 					(reg_q2399 AND symb_decoder(16#52#));
reg_q2401_init <= '0' ;
	p_reg_q2401: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2401 <= reg_q2401_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2401 <= reg_q2401_init;
        else
          reg_q2401 <= reg_q2401_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q92_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q91 AND symb_decoder(16#0a#)) OR
 					(reg_q91 AND symb_decoder(16#0d#));
reg_q92_init <= '0' ;
	p_reg_q92: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q92 <= reg_q92_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q92 <= reg_q92_init;
        else
          reg_q92 <= reg_q92_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q960_in <= (reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q960 AND symb_decoder(16#34#)) OR
 					(reg_q960 AND symb_decoder(16#32#)) OR
 					(reg_q960 AND symb_decoder(16#30#)) OR
 					(reg_q960 AND symb_decoder(16#38#)) OR
 					(reg_q960 AND symb_decoder(16#35#)) OR
 					(reg_q960 AND symb_decoder(16#39#)) OR
 					(reg_q960 AND symb_decoder(16#31#)) OR
 					(reg_q960 AND symb_decoder(16#33#)) OR
 					(reg_q960 AND symb_decoder(16#37#)) OR
 					(reg_q960 AND symb_decoder(16#36#)) OR
 					(reg_q959 AND symb_decoder(16#32#)) OR
 					(reg_q959 AND symb_decoder(16#30#)) OR
 					(reg_q959 AND symb_decoder(16#38#)) OR
 					(reg_q959 AND symb_decoder(16#33#)) OR
 					(reg_q959 AND symb_decoder(16#35#)) OR
 					(reg_q959 AND symb_decoder(16#34#)) OR
 					(reg_q959 AND symb_decoder(16#31#)) OR
 					(reg_q959 AND symb_decoder(16#39#)) OR
 					(reg_q959 AND symb_decoder(16#37#)) OR
 					(reg_q959 AND symb_decoder(16#36#));
reg_q960_init <= '0' ;
	p_reg_q960: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q960 <= reg_q960_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q960 <= reg_q960_init;
        else
          reg_q960 <= reg_q960_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q204_in <= (reg_q202 AND symb_decoder(16#56#)) OR
 					(reg_q202 AND symb_decoder(16#76#));
reg_q204_init <= '0' ;
	p_reg_q204: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q204 <= reg_q204_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q204 <= reg_q204_init;
        else
          reg_q204 <= reg_q204_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q206_in <= (reg_q204 AND symb_decoder(16#52#)) OR
 					(reg_q204 AND symb_decoder(16#72#));
reg_q206_init <= '0' ;
	p_reg_q206: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q206 <= reg_q206_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q206 <= reg_q206_init;
        else
          reg_q206 <= reg_q206_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1566_in <= (reg_q1564 AND symb_decoder(16#53#)) OR
 					(reg_q1564 AND symb_decoder(16#73#));
reg_q1566_init <= '0' ;
	p_reg_q1566: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1566 <= reg_q1566_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1566 <= reg_q1566_init;
        else
          reg_q1566 <= reg_q1566_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1568_in <= (reg_q1566 AND symb_decoder(16#49#)) OR
 					(reg_q1566 AND symb_decoder(16#69#));
reg_q1568_init <= '0' ;
	p_reg_q1568: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1568 <= reg_q1568_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1568 <= reg_q1568_init;
        else
          reg_q1568 <= reg_q1568_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2502_in <= (reg_q2695 AND symb_decoder(16#2a#));
reg_q2502_init <= '0' ;
	p_reg_q2502: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2502 <= reg_q2502_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2502 <= reg_q2502_init;
        else
          reg_q2502 <= reg_q2502_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2262_in <= (reg_q2260 AND symb_decoder(16#70#)) OR
 					(reg_q2260 AND symb_decoder(16#50#));
reg_q2262_init <= '0' ;
	p_reg_q2262: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2262 <= reg_q2262_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2262 <= reg_q2262_init;
        else
          reg_q2262 <= reg_q2262_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2264_in <= (reg_q2262 AND symb_decoder(16#74#)) OR
 					(reg_q2262 AND symb_decoder(16#54#));
reg_q2264_init <= '0' ;
	p_reg_q2264: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2264 <= reg_q2264_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2264 <= reg_q2264_init;
        else
          reg_q2264 <= reg_q2264_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q430_in <= (reg_q428 AND symb_decoder(16#55#)) OR
 					(reg_q428 AND symb_decoder(16#75#));
reg_q430_init <= '0' ;
	p_reg_q430: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q430 <= reg_q430_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q430 <= reg_q430_init;
        else
          reg_q430 <= reg_q430_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q432_in <= (reg_q430 AND symb_decoder(16#6e#)) OR
 					(reg_q430 AND symb_decoder(16#4e#));
reg_q432_init <= '0' ;
	p_reg_q432: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q432 <= reg_q432_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q432 <= reg_q432_init;
        else
          reg_q432 <= reg_q432_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2427_in <= (reg_q2427 AND symb_decoder(16#20#)) OR
 					(reg_q2427 AND symb_decoder(16#0a#)) OR
 					(reg_q2427 AND symb_decoder(16#0d#)) OR
 					(reg_q2427 AND symb_decoder(16#0c#)) OR
 					(reg_q2427 AND symb_decoder(16#09#)) OR
 					(reg_q2425 AND symb_decoder(16#0d#)) OR
 					(reg_q2425 AND symb_decoder(16#0a#)) OR
 					(reg_q2425 AND symb_decoder(16#20#)) OR
 					(reg_q2425 AND symb_decoder(16#0c#)) OR
 					(reg_q2425 AND symb_decoder(16#09#));
reg_q2427_init <= '0' ;
	p_reg_q2427: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2427 <= reg_q2427_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2427 <= reg_q2427_init;
        else
          reg_q2427 <= reg_q2427_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2371_in <= (reg_q2369 AND symb_decoder(16#76#)) OR
 					(reg_q2369 AND symb_decoder(16#56#));
reg_q2371_init <= '0' ;
	p_reg_q2371: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2371 <= reg_q2371_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2371 <= reg_q2371_init;
        else
          reg_q2371 <= reg_q2371_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1645_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1644 AND symb_decoder(16#0d#)) OR
 					(reg_q1644 AND symb_decoder(16#0a#));
reg_q1645_init <= '0' ;
	p_reg_q1645: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1645 <= reg_q1645_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1645 <= reg_q1645_init;
        else
          reg_q1645 <= reg_q1645_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1646_in <= (reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q1645 AND symb_decoder(16#72#)) OR
 					(reg_q1645 AND symb_decoder(16#52#));
reg_q1646_init <= '0' ;
	p_reg_q1646: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1646 <= reg_q1646_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1646 <= reg_q1646_init;
        else
          reg_q1646 <= reg_q1646_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2290_in <= (reg_q2288 AND symb_decoder(16#73#)) OR
 					(reg_q2288 AND symb_decoder(16#53#));
reg_q2290_init <= '0' ;
	p_reg_q2290: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2290 <= reg_q2290_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2290 <= reg_q2290_init;
        else
          reg_q2290 <= reg_q2290_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2292_in <= (reg_q2290 AND symb_decoder(16#45#)) OR
 					(reg_q2290 AND symb_decoder(16#65#));
reg_q2292_init <= '0' ;
	p_reg_q2292: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2292 <= reg_q2292_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2292 <= reg_q2292_init;
        else
          reg_q2292 <= reg_q2292_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2046_in <= (reg_q2044 AND symb_decoder(16#4f#)) OR
 					(reg_q2044 AND symb_decoder(16#6f#));
reg_q2046_init <= '0' ;
	p_reg_q2046: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2046 <= reg_q2046_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2046 <= reg_q2046_init;
        else
          reg_q2046 <= reg_q2046_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2064_in <= (reg_q2062 AND symb_decoder(16#32#));
reg_q2064_init <= '0' ;
	p_reg_q2064: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2064 <= reg_q2064_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2064 <= reg_q2064_init;
        else
          reg_q2064 <= reg_q2064_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1427_in <= (reg_q1425 AND symb_decoder(16#61#)) OR
 					(reg_q1425 AND symb_decoder(16#41#));
reg_q1427_init <= '0' ;
	p_reg_q1427: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1427 <= reg_q1427_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1427 <= reg_q1427_init;
        else
          reg_q1427 <= reg_q1427_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1429_in <= (reg_q1427 AND symb_decoder(16#74#)) OR
 					(reg_q1427 AND symb_decoder(16#54#));
reg_q1429_init <= '0' ;
	p_reg_q1429: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1429 <= reg_q1429_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1429 <= reg_q1429_init;
        else
          reg_q1429 <= reg_q1429_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2038_in <= (reg_q2036 AND symb_decoder(16#45#)) OR
 					(reg_q2036 AND symb_decoder(16#65#));
reg_q2038_init <= '0' ;
	p_reg_q2038: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2038 <= reg_q2038_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2038 <= reg_q2038_init;
        else
          reg_q2038 <= reg_q2038_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2040_in <= (reg_q2038 AND symb_decoder(16#0c#)) OR
 					(reg_q2038 AND symb_decoder(16#09#)) OR
 					(reg_q2038 AND symb_decoder(16#0a#)) OR
 					(reg_q2038 AND symb_decoder(16#0d#)) OR
 					(reg_q2038 AND symb_decoder(16#20#)) OR
 					(reg_q2040 AND symb_decoder(16#0a#)) OR
 					(reg_q2040 AND symb_decoder(16#09#)) OR
 					(reg_q2040 AND symb_decoder(16#0c#)) OR
 					(reg_q2040 AND symb_decoder(16#20#)) OR
 					(reg_q2040 AND symb_decoder(16#0d#));
reg_q2040_init <= '0' ;
	p_reg_q2040: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2040 <= reg_q2040_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2040 <= reg_q2040_init;
        else
          reg_q2040 <= reg_q2040_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2379_in <= (reg_q2377 AND symb_decoder(16#0d#));
reg_q2379_init <= '0' ;
	p_reg_q2379: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2379 <= reg_q2379_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2379 <= reg_q2379_init;
        else
          reg_q2379 <= reg_q2379_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q99_in <= (reg_q97 AND symb_decoder(16#ac#));
reg_q99_init <= '0' ;
	p_reg_q99: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q99 <= reg_q99_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q99 <= reg_q99_init;
        else
          reg_q99 <= reg_q99_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1880_in <= (reg_q1880 AND symb_decoder(16#0d#)) OR
 					(reg_q1880 AND symb_decoder(16#09#)) OR
 					(reg_q1880 AND symb_decoder(16#0a#)) OR
 					(reg_q1880 AND symb_decoder(16#0c#)) OR
 					(reg_q1880 AND symb_decoder(16#20#)) OR
 					(reg_q1878 AND symb_decoder(16#0c#)) OR
 					(reg_q1878 AND symb_decoder(16#09#)) OR
 					(reg_q1878 AND symb_decoder(16#20#)) OR
 					(reg_q1878 AND symb_decoder(16#0a#)) OR
 					(reg_q1878 AND symb_decoder(16#0d#));
reg_q1880_init <= '0' ;
	p_reg_q1880: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1880 <= reg_q1880_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1880 <= reg_q1880_init;
        else
          reg_q1880 <= reg_q1880_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1171_in <= (reg_q1169 AND symb_decoder(16#63#)) OR
 					(reg_q1169 AND symb_decoder(16#43#));
reg_q1171_init <= '0' ;
	p_reg_q1171: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1171 <= reg_q1171_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1171 <= reg_q1171_init;
        else
          reg_q1171 <= reg_q1171_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q870_in <= (reg_q868 AND symb_decoder(16#53#)) OR
 					(reg_q868 AND symb_decoder(16#73#));
reg_q870_init <= '0' ;
	p_reg_q870: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q870 <= reg_q870_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q870 <= reg_q870_init;
        else
          reg_q870 <= reg_q870_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q872_in <= (reg_q870 AND symb_decoder(16#54#)) OR
 					(reg_q870 AND symb_decoder(16#74#));
reg_q872_init <= '0' ;
	p_reg_q872: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q872 <= reg_q872_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q872 <= reg_q872_init;
        else
          reg_q872 <= reg_q872_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1064_in <= (reg_q1062 AND symb_decoder(16#74#)) OR
 					(reg_q1062 AND symb_decoder(16#54#));
reg_q1064_init <= '0' ;
	p_reg_q1064: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1064 <= reg_q1064_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1064 <= reg_q1064_init;
        else
          reg_q1064 <= reg_q1064_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2353_in <= (reg_q2351 AND symb_decoder(16#4d#)) OR
 					(reg_q2351 AND symb_decoder(16#6d#));
reg_q2353_init <= '0' ;
	p_reg_q2353: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2353 <= reg_q2353_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2353 <= reg_q2353_init;
        else
          reg_q2353 <= reg_q2353_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1718_in <= (reg_q1716 AND symb_decoder(16#2e#));
reg_q1718_init <= '0' ;
	p_reg_q1718: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1718 <= reg_q1718_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1718 <= reg_q1718_init;
        else
          reg_q1718 <= reg_q1718_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1828_in <= (reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q1826 AND symb_decoder(16#73#)) OR
 					(reg_q1826 AND symb_decoder(16#53#));
reg_q1828_init <= '0' ;
	p_reg_q1828: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1828 <= reg_q1828_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1828 <= reg_q1828_init;
        else
          reg_q1828 <= reg_q1828_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q70_in <= (reg_q68 AND symb_decoder(16#52#)) OR
 					(reg_q68 AND symb_decoder(16#72#));
reg_q70_init <= '0' ;
	p_reg_q70: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q70 <= reg_q70_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q70 <= reg_q70_init;
        else
          reg_q70 <= reg_q70_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q72_in <= (reg_q70 AND symb_decoder(16#09#)) OR
 					(reg_q70 AND symb_decoder(16#0a#)) OR
 					(reg_q70 AND symb_decoder(16#0d#)) OR
 					(reg_q70 AND symb_decoder(16#20#)) OR
 					(reg_q70 AND symb_decoder(16#0c#)) OR
 					(reg_q72 AND symb_decoder(16#09#)) OR
 					(reg_q72 AND symb_decoder(16#0c#)) OR
 					(reg_q72 AND symb_decoder(16#20#)) OR
 					(reg_q72 AND symb_decoder(16#0a#)) OR
 					(reg_q72 AND symb_decoder(16#0d#));
reg_q72_init <= '0' ;
	p_reg_q72: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q72 <= reg_q72_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q72 <= reg_q72_init;
        else
          reg_q72 <= reg_q72_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2119_in <= (reg_q2117 AND symb_decoder(16#45#)) OR
 					(reg_q2117 AND symb_decoder(16#65#));
reg_q2119_init <= '0' ;
	p_reg_q2119: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2119 <= reg_q2119_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2119 <= reg_q2119_init;
        else
          reg_q2119 <= reg_q2119_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2121_in <= (reg_q2119 AND symb_decoder(16#72#)) OR
 					(reg_q2119 AND symb_decoder(16#52#));
reg_q2121_init <= '0' ;
	p_reg_q2121: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2121 <= reg_q2121_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2121 <= reg_q2121_init;
        else
          reg_q2121 <= reg_q2121_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1343_in <= (reg_q1341 AND symb_decoder(16#2e#));
reg_q1343_init <= '0' ;
	p_reg_q1343: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1343 <= reg_q1343_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1343 <= reg_q1343_init;
        else
          reg_q1343 <= reg_q1343_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1112_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1111 AND symb_decoder(16#0a#)) OR
 					(reg_q1111 AND symb_decoder(16#0d#));
reg_q1112_init <= '0' ;
	p_reg_q1112: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1112 <= reg_q1112_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1112 <= reg_q1112_init;
        else
          reg_q1112 <= reg_q1112_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2227_in <= (reg_q2225 AND symb_decoder(16#68#)) OR
 					(reg_q2225 AND symb_decoder(16#48#));
reg_q2227_init <= '0' ;
	p_reg_q2227: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2227 <= reg_q2227_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2227 <= reg_q2227_init;
        else
          reg_q2227 <= reg_q2227_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1037_in <= (reg_q1035 AND symb_decoder(16#53#)) OR
 					(reg_q1035 AND symb_decoder(16#73#));
reg_q1037_init <= '0' ;
	p_reg_q1037: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1037 <= reg_q1037_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1037 <= reg_q1037_init;
        else
          reg_q1037 <= reg_q1037_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1039_in <= (reg_q1037 AND symb_decoder(16#45#)) OR
 					(reg_q1037 AND symb_decoder(16#65#));
reg_q1039_init <= '0' ;
	p_reg_q1039: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1039 <= reg_q1039_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1039 <= reg_q1039_init;
        else
          reg_q1039 <= reg_q1039_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1161_in <= (reg_q1159 AND symb_decoder(16#63#)) OR
 					(reg_q1159 AND symb_decoder(16#43#));
reg_q1161_init <= '0' ;
	p_reg_q1161: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1161 <= reg_q1161_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1161 <= reg_q1161_init;
        else
          reg_q1161 <= reg_q1161_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1163_in <= (reg_q1161 AND symb_decoder(16#6f#)) OR
 					(reg_q1161 AND symb_decoder(16#4f#));
reg_q1163_init <= '0' ;
	p_reg_q1163: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1163 <= reg_q1163_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1163 <= reg_q1163_init;
        else
          reg_q1163 <= reg_q1163_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1399_in <= (reg_q1397 AND symb_decoder(16#79#)) OR
 					(reg_q1397 AND symb_decoder(16#59#));
reg_q1399_init <= '0' ;
	p_reg_q1399: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1399 <= reg_q1399_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1399 <= reg_q1399_init;
        else
          reg_q1399 <= reg_q1399_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1401_in <= (reg_q1399 AND symb_decoder(16#62#)) OR
 					(reg_q1399 AND symb_decoder(16#42#));
reg_q1401_init <= '0' ;
	p_reg_q1401: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1401 <= reg_q1401_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1401 <= reg_q1401_init;
        else
          reg_q1401 <= reg_q1401_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1582_in <= (reg_q1580 AND symb_decoder(16#0d#));
reg_q1582_init <= '0' ;
	p_reg_q1582: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1582 <= reg_q1582_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1582 <= reg_q1582_init;
        else
          reg_q1582 <= reg_q1582_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1584_in <= (reg_q1582 AND symb_decoder(16#0a#));
reg_q1584_init <= '0' ;
	p_reg_q1584: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1584 <= reg_q1584_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1584 <= reg_q1584_init;
        else
          reg_q1584 <= reg_q1584_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q12_in <= (reg_q10 AND symb_decoder(16#4c#)) OR
 					(reg_q10 AND symb_decoder(16#6c#));
reg_q12_init <= '0' ;
	p_reg_q12: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q12 <= reg_q12_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q12 <= reg_q12_init;
        else
          reg_q12 <= reg_q12_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q143_in <= (reg_q141 AND symb_decoder(16#54#)) OR
 					(reg_q141 AND symb_decoder(16#74#));
reg_q143_init <= '0' ;
	p_reg_q143: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q143 <= reg_q143_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q143 <= reg_q143_init;
        else
          reg_q143 <= reg_q143_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1504_in <= (reg_q1504 AND symb_decoder(16#0d#)) OR
 					(reg_q1504 AND symb_decoder(16#0a#)) OR
 					(reg_q1504 AND symb_decoder(16#0c#)) OR
 					(reg_q1504 AND symb_decoder(16#09#)) OR
 					(reg_q1504 AND symb_decoder(16#20#)) OR
 					(reg_q1502 AND symb_decoder(16#0a#)) OR
 					(reg_q1502 AND symb_decoder(16#20#)) OR
 					(reg_q1502 AND symb_decoder(16#0c#)) OR
 					(reg_q1502 AND symb_decoder(16#0d#)) OR
 					(reg_q1502 AND symb_decoder(16#09#));
reg_q1504_init <= '0' ;
	p_reg_q1504: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1504 <= reg_q1504_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1504 <= reg_q1504_init;
        else
          reg_q1504 <= reg_q1504_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1506_in <= (reg_q1504 AND symb_decoder(16#76#)) OR
 					(reg_q1504 AND symb_decoder(16#56#));
reg_q1506_init <= '0' ;
	p_reg_q1506: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1506 <= reg_q1506_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1506 <= reg_q1506_init;
        else
          reg_q1506 <= reg_q1506_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q208_in <= (reg_q206 AND symb_decoder(16#5e#));
reg_q208_init <= '0' ;
	p_reg_q208: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q208 <= reg_q208_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q208 <= reg_q208_init;
        else
          reg_q208 <= reg_q208_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q210_in <= (reg_q208 AND symb_decoder(16#5e#));
reg_q210_init <= '0' ;
	p_reg_q210: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q210 <= reg_q210_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q210 <= reg_q210_init;
        else
          reg_q210 <= reg_q210_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2170_in <= (reg_q2168 AND symb_decoder(16#4f#)) OR
 					(reg_q2168 AND symb_decoder(16#6f#));
reg_q2170_init <= '0' ;
	p_reg_q2170: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2170 <= reg_q2170_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2170 <= reg_q2170_init;
        else
          reg_q2170 <= reg_q2170_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1844_in <= (reg_q1842 AND symb_decoder(16#65#)) OR
 					(reg_q1842 AND symb_decoder(16#45#));
reg_q1844_init <= '0' ;
	p_reg_q1844: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1844 <= reg_q1844_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1844 <= reg_q1844_init;
        else
          reg_q1844 <= reg_q1844_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q357_in <= (reg_q355 AND symb_decoder(16#76#)) OR
 					(reg_q355 AND symb_decoder(16#56#));
reg_q357_init <= '0' ;
	p_reg_q357: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q357 <= reg_q357_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q357 <= reg_q357_init;
        else
          reg_q357 <= reg_q357_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q359_in <= (reg_q357 AND symb_decoder(16#65#)) OR
 					(reg_q357 AND symb_decoder(16#45#));
reg_q359_init <= '0' ;
	p_reg_q359: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q359 <= reg_q359_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q359 <= reg_q359_init;
        else
          reg_q359 <= reg_q359_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q669_in <= (reg_q667 AND symb_decoder(16#4f#)) OR
 					(reg_q667 AND symb_decoder(16#6f#));
reg_q669_init <= '0' ;
	p_reg_q669: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q669 <= reg_q669_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q669 <= reg_q669_init;
        else
          reg_q669 <= reg_q669_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1942_in <= (reg_q1940 AND symb_decoder(16#50#)) OR
 					(reg_q1940 AND symb_decoder(16#70#));
reg_q1942_init <= '0' ;
	p_reg_q1942: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1942 <= reg_q1942_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1942 <= reg_q1942_init;
        else
          reg_q1942 <= reg_q1942_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1944_in <= (reg_q1942 AND symb_decoder(16#59#)) OR
 					(reg_q1942 AND symb_decoder(16#79#));
reg_q1944_init <= '0' ;
	p_reg_q1944: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1944 <= reg_q1944_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1944 <= reg_q1944_init;
        else
          reg_q1944 <= reg_q1944_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1029_in <= (reg_q1027 AND symb_decoder(16#53#)) OR
 					(reg_q1027 AND symb_decoder(16#73#));
reg_q1029_init <= '0' ;
	p_reg_q1029: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1029 <= reg_q1029_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1029 <= reg_q1029_init;
        else
          reg_q1029 <= reg_q1029_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1031_in <= (reg_q1029 AND symb_decoder(16#69#)) OR
 					(reg_q1029 AND symb_decoder(16#49#));
reg_q1031_init <= '0' ;
	p_reg_q1031: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1031 <= reg_q1031_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1031 <= reg_q1031_init;
        else
          reg_q1031 <= reg_q1031_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1361_in <= (reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q1359 AND symb_decoder(16#48#)) OR
 					(reg_q1359 AND symb_decoder(16#68#));
reg_q1361_init <= '0' ;
	p_reg_q1361: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1361 <= reg_q1361_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1361 <= reg_q1361_init;
        else
          reg_q1361 <= reg_q1361_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q383_in <= (reg_q381 AND symb_decoder(16#55#)) OR
 					(reg_q381 AND symb_decoder(16#75#));
reg_q383_init <= '0' ;
	p_reg_q383: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q383 <= reg_q383_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q383 <= reg_q383_init;
        else
          reg_q383 <= reg_q383_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q642_in <= (reg_q640 AND symb_decoder(16#6e#)) OR
 					(reg_q640 AND symb_decoder(16#4e#));
reg_q642_init <= '0' ;
	p_reg_q642: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q642 <= reg_q642_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q642 <= reg_q642_init;
        else
          reg_q642 <= reg_q642_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1604_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1603 AND symb_decoder(16#0d#)) OR
 					(reg_q1603 AND symb_decoder(16#0a#));
reg_q1604_init <= '0' ;
	p_reg_q1604: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1604 <= reg_q1604_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1604 <= reg_q1604_init;
        else
          reg_q1604 <= reg_q1604_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1664_in <= (reg_q1662 AND symb_decoder(16#2e#));
reg_q1664_init <= '0' ;
	p_reg_q1664: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1664 <= reg_q1664_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1664 <= reg_q1664_init;
        else
          reg_q1664 <= reg_q1664_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1932_in <= (reg_q1930 AND symb_decoder(16#73#)) OR
 					(reg_q1930 AND symb_decoder(16#53#));
reg_q1932_init <= '0' ;
	p_reg_q1932: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1932 <= reg_q1932_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1932 <= reg_q1932_init;
        else
          reg_q1932 <= reg_q1932_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2497_in <= (reg_q2495 AND symb_decoder(16#2a#));
reg_q2497_init <= '0' ;
	p_reg_q2497: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2497 <= reg_q2497_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2497 <= reg_q2497_init;
        else
          reg_q2497 <= reg_q2497_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q626_in <= (reg_q624 AND symb_decoder(16#76#)) OR
 					(reg_q624 AND symb_decoder(16#56#));
reg_q626_init <= '0' ;
	p_reg_q626: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q626 <= reg_q626_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q626 <= reg_q626_init;
        else
          reg_q626 <= reg_q626_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2109_in <= (reg_q2107 AND symb_decoder(16#78#)) OR
 					(reg_q2107 AND symb_decoder(16#58#));
reg_q2109_init <= '0' ;
	p_reg_q2109: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2109 <= reg_q2109_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2109 <= reg_q2109_init;
        else
          reg_q2109 <= reg_q2109_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2111_in <= (reg_q2109 AND symb_decoder(16#09#)) OR
 					(reg_q2109 AND symb_decoder(16#20#)) OR
 					(reg_q2109 AND symb_decoder(16#0d#)) OR
 					(reg_q2109 AND symb_decoder(16#0a#)) OR
 					(reg_q2109 AND symb_decoder(16#0c#)) OR
 					(reg_q2111 AND symb_decoder(16#0c#)) OR
 					(reg_q2111 AND symb_decoder(16#0d#)) OR
 					(reg_q2111 AND symb_decoder(16#0a#)) OR
 					(reg_q2111 AND symb_decoder(16#09#)) OR
 					(reg_q2111 AND symb_decoder(16#20#));
reg_q2111_init <= '0' ;
	p_reg_q2111: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2111 <= reg_q2111_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2111 <= reg_q2111_init;
        else
          reg_q2111 <= reg_q2111_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2585_in <= (reg_q2583 AND symb_decoder(16#0a#));
reg_q2585_init <= '0' ;
	p_reg_q2585: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2585 <= reg_q2585_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2585 <= reg_q2585_init;
        else
          reg_q2585 <= reg_q2585_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2587_in <= (reg_q2585 AND symb_decoder(16#63#)) OR
 					(reg_q2585 AND symb_decoder(16#43#));
reg_q2587_init <= '0' ;
	p_reg_q2587: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2587 <= reg_q2587_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2587 <= reg_q2587_init;
        else
          reg_q2587 <= reg_q2587_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q307_in <= (reg_q305 AND symb_decoder(16#4e#)) OR
 					(reg_q305 AND symb_decoder(16#6e#));
reg_q307_init <= '0' ;
	p_reg_q307: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q307 <= reg_q307_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q307 <= reg_q307_init;
        else
          reg_q307 <= reg_q307_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1533_in <= (reg_q1531 AND symb_decoder(16#53#)) OR
 					(reg_q1531 AND symb_decoder(16#73#));
reg_q1533_init <= '0' ;
	p_reg_q1533: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1533 <= reg_q1533_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1533 <= reg_q1533_init;
        else
          reg_q1533 <= reg_q1533_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2575_in <= (reg_q2573 AND symb_decoder(16#52#)) OR
 					(reg_q2573 AND symb_decoder(16#72#));
reg_q2575_init <= '0' ;
	p_reg_q2575: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2575 <= reg_q2575_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2575 <= reg_q2575_init;
        else
          reg_q2575 <= reg_q2575_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q518_in <= (reg_q516 AND symb_decoder(16#50#)) OR
 					(reg_q516 AND symb_decoder(16#70#));
reg_q518_init <= '0' ;
	p_reg_q518: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q518 <= reg_q518_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q518 <= reg_q518_init;
        else
          reg_q518 <= reg_q518_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q789_in <= (reg_q787 AND symb_decoder(16#66#)) OR
 					(reg_q787 AND symb_decoder(16#46#));
reg_q789_init <= '0' ;
	p_reg_q789: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q789 <= reg_q789_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q789 <= reg_q789_init;
        else
          reg_q789 <= reg_q789_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1734_in <= (reg_q1732 AND symb_decoder(16#70#)) OR
 					(reg_q1732 AND symb_decoder(16#50#));
reg_q1734_init <= '0' ;
	p_reg_q1734: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1734 <= reg_q1734_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1734 <= reg_q1734_init;
        else
          reg_q1734 <= reg_q1734_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1736_in <= (reg_q1734 AND symb_decoder(16#0a#)) OR
 					(reg_q1734 AND symb_decoder(16#20#)) OR
 					(reg_q1734 AND symb_decoder(16#09#)) OR
 					(reg_q1734 AND symb_decoder(16#0c#)) OR
 					(reg_q1734 AND symb_decoder(16#0d#)) OR
 					(reg_q1736 AND symb_decoder(16#0c#)) OR
 					(reg_q1736 AND symb_decoder(16#0d#)) OR
 					(reg_q1736 AND symb_decoder(16#20#)) OR
 					(reg_q1736 AND symb_decoder(16#0a#)) OR
 					(reg_q1736 AND symb_decoder(16#09#));
reg_q1736_init <= '0' ;
	p_reg_q1736: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1736 <= reg_q1736_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1736 <= reg_q1736_init;
        else
          reg_q1736 <= reg_q1736_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2221_in <= (reg_q2219 AND symb_decoder(16#72#)) OR
 					(reg_q2219 AND symb_decoder(16#52#));
reg_q2221_init <= '0' ;
	p_reg_q2221: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2221 <= reg_q2221_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2221 <= reg_q2221_init;
        else
          reg_q2221 <= reg_q2221_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2223_in <= (reg_q2221 AND symb_decoder(16#41#)) OR
 					(reg_q2221 AND symb_decoder(16#61#));
reg_q2223_init <= '0' ;
	p_reg_q2223: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2223 <= reg_q2223_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2223 <= reg_q2223_init;
        else
          reg_q2223 <= reg_q2223_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q598_in <= (reg_q596 AND symb_decoder(16#70#)) OR
 					(reg_q596 AND symb_decoder(16#50#));
reg_q598_init <= '0' ;
	p_reg_q598: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q598 <= reg_q598_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q598 <= reg_q598_init;
        else
          reg_q598 <= reg_q598_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q600_in <= (reg_q598 AND symb_decoder(16#72#)) OR
 					(reg_q598 AND symb_decoder(16#52#));
reg_q600_init <= '0' ;
	p_reg_q600: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q600 <= reg_q600_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q600 <= reg_q600_init;
        else
          reg_q600 <= reg_q600_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1832_in <= (reg_q1830 AND symb_decoder(16#48#)) OR
 					(reg_q1830 AND symb_decoder(16#68#));
reg_q1832_init <= '0' ;
	p_reg_q1832: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1832 <= reg_q1832_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1832 <= reg_q1832_init;
        else
          reg_q1832 <= reg_q1832_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1834_in <= (reg_q1832 AND symb_decoder(16#77#)) OR
 					(reg_q1832 AND symb_decoder(16#57#));
reg_q1834_init <= '0' ;
	p_reg_q1834: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1834 <= reg_q1834_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1834 <= reg_q1834_init;
        else
          reg_q1834 <= reg_q1834_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q64_in <= (reg_q62 AND symb_decoder(16#48#)) OR
 					(reg_q62 AND symb_decoder(16#68#));
reg_q64_init <= '0' ;
	p_reg_q64: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q64 <= reg_q64_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q64 <= reg_q64_init;
        else
          reg_q64 <= reg_q64_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q66_in <= (reg_q64 AND symb_decoder(16#74#)) OR
 					(reg_q64 AND symb_decoder(16#54#));
reg_q66_init <= '0' ;
	p_reg_q66: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q66 <= reg_q66_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q66 <= reg_q66_init;
        else
          reg_q66 <= reg_q66_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1015_in <= (reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q1014 AND symb_decoder(16#65#)) OR
 					(reg_q1014 AND symb_decoder(16#45#));
reg_q1015_init <= '0' ;
	p_reg_q1015: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1015 <= reg_q1015_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1015 <= reg_q1015_init;
        else
          reg_q1015 <= reg_q1015_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2413_in <= (reg_q2411 AND symb_decoder(16#53#)) OR
 					(reg_q2411 AND symb_decoder(16#73#));
reg_q2413_init <= '0' ;
	p_reg_q2413: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2413 <= reg_q2413_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2413 <= reg_q2413_init;
        else
          reg_q2413 <= reg_q2413_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2385_in <= (reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2383 AND symb_decoder(16#23#));
reg_q2385_init <= '0' ;
	p_reg_q2385: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2385 <= reg_q2385_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2385 <= reg_q2385_init;
        else
          reg_q2385 <= reg_q2385_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2387_in <= (reg_q2385 AND symb_decoder(16#31#));
reg_q2387_init <= '0' ;
	p_reg_q2387: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2387 <= reg_q2387_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2387 <= reg_q2387_init;
        else
          reg_q2387 <= reg_q2387_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q131_in <= (reg_q129 AND symb_decoder(16#43#)) OR
 					(reg_q129 AND symb_decoder(16#63#));
reg_q131_init <= '0' ;
	p_reg_q131: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q131 <= reg_q131_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q131 <= reg_q131_init;
        else
          reg_q131 <= reg_q131_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2217_in <= (reg_q2215 AND symb_decoder(16#6e#)) OR
 					(reg_q2215 AND symb_decoder(16#4e#));
reg_q2217_init <= '0' ;
	p_reg_q2217: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2217 <= reg_q2217_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2217 <= reg_q2217_init;
        else
          reg_q2217 <= reg_q2217_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q38_in <= (reg_q36 AND symb_decoder(16#64#)) OR
 					(reg_q36 AND symb_decoder(16#44#));
reg_q38_init <= '0' ;
	p_reg_q38: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q38 <= reg_q38_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q38 <= reg_q38_init;
        else
          reg_q38 <= reg_q38_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q40_in <= (reg_q38 AND symb_decoder(16#2e#));
reg_q40_init <= '0' ;
	p_reg_q40: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q40 <= reg_q40_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q40 <= reg_q40_init;
        else
          reg_q40 <= reg_q40_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q155_in <= (reg_q153 AND symb_decoder(16#63#)) OR
 					(reg_q153 AND symb_decoder(16#43#));
reg_q155_init <= '0' ;
	p_reg_q155: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q155 <= reg_q155_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q155 <= reg_q155_init;
        else
          reg_q155 <= reg_q155_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q157_in <= (reg_q155 AND symb_decoder(16#63#)) OR
 					(reg_q155 AND symb_decoder(16#43#));
reg_q157_init <= '0' ;
	p_reg_q157: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q157 <= reg_q157_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q157 <= reg_q157_init;
        else
          reg_q157 <= reg_q157_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q373_in <= (reg_q371 AND symb_decoder(16#22#));
reg_q373_init <= '0' ;
	p_reg_q373: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q373 <= reg_q373_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q373 <= reg_q373_init;
        else
          reg_q373 <= reg_q373_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q36_in <= (reg_q34 AND symb_decoder(16#45#)) OR
 					(reg_q34 AND symb_decoder(16#65#));
reg_q36_init <= '0' ;
	p_reg_q36: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q36 <= reg_q36_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q36 <= reg_q36_init;
        else
          reg_q36 <= reg_q36_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1550_in <= (reg_q1548 AND symb_decoder(16#74#)) OR
 					(reg_q1548 AND symb_decoder(16#54#));
reg_q1550_init <= '0' ;
	p_reg_q1550: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1550 <= reg_q1550_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1550 <= reg_q1550_init;
        else
          reg_q1550 <= reg_q1550_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1552_in <= (reg_q1550 AND symb_decoder(16#73#)) OR
 					(reg_q1550 AND symb_decoder(16#53#));
reg_q1552_init <= '0' ;
	p_reg_q1552: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1552 <= reg_q1552_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1552 <= reg_q1552_init;
        else
          reg_q1552 <= reg_q1552_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q834_in <= (reg_q832 AND symb_decoder(16#2e#));
reg_q834_init <= '0' ;
	p_reg_q834: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q834 <= reg_q834_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q834 <= reg_q834_init;
        else
          reg_q834 <= reg_q834_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q923_in <= (reg_q921 AND symb_decoder(16#45#)) OR
 					(reg_q921 AND symb_decoder(16#65#));
reg_q923_init <= '0' ;
	p_reg_q923: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q923 <= reg_q923_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q923 <= reg_q923_init;
        else
          reg_q923 <= reg_q923_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q925_in <= (reg_q923 AND symb_decoder(16#52#)) OR
 					(reg_q923 AND symb_decoder(16#72#));
reg_q925_init <= '0' ;
	p_reg_q925: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q925 <= reg_q925_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q925 <= reg_q925_init;
        else
          reg_q925 <= reg_q925_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1820_in <= (reg_q1818 AND symb_decoder(16#39#)) OR
 					(reg_q1818 AND symb_decoder(16#31#)) OR
 					(reg_q1818 AND symb_decoder(16#38#)) OR
 					(reg_q1818 AND symb_decoder(16#34#)) OR
 					(reg_q1818 AND symb_decoder(16#30#)) OR
 					(reg_q1818 AND symb_decoder(16#37#)) OR
 					(reg_q1818 AND symb_decoder(16#33#)) OR
 					(reg_q1818 AND symb_decoder(16#32#)) OR
 					(reg_q1818 AND symb_decoder(16#35#)) OR
 					(reg_q1818 AND symb_decoder(16#36#)) OR
 					(reg_q1820 AND symb_decoder(16#36#)) OR
 					(reg_q1820 AND symb_decoder(16#39#)) OR
 					(reg_q1820 AND symb_decoder(16#35#)) OR
 					(reg_q1820 AND symb_decoder(16#37#)) OR
 					(reg_q1820 AND symb_decoder(16#30#)) OR
 					(reg_q1820 AND symb_decoder(16#32#)) OR
 					(reg_q1820 AND symb_decoder(16#31#)) OR
 					(reg_q1820 AND symb_decoder(16#38#)) OR
 					(reg_q1820 AND symb_decoder(16#34#)) OR
 					(reg_q1820 AND symb_decoder(16#33#));
reg_q1820_init <= '0' ;
	p_reg_q1820: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1820 <= reg_q1820_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1820 <= reg_q1820_init;
        else
          reg_q1820 <= reg_q1820_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1143_in <= (reg_q1143 AND symb_decoder(16#34#)) OR
 					(reg_q1143 AND symb_decoder(16#32#)) OR
 					(reg_q1143 AND symb_decoder(16#38#)) OR
 					(reg_q1143 AND symb_decoder(16#39#)) OR
 					(reg_q1143 AND symb_decoder(16#33#)) OR
 					(reg_q1143 AND symb_decoder(16#30#)) OR
 					(reg_q1143 AND symb_decoder(16#37#)) OR
 					(reg_q1143 AND symb_decoder(16#31#)) OR
 					(reg_q1143 AND symb_decoder(16#36#)) OR
 					(reg_q1143 AND symb_decoder(16#35#)) OR
 					(reg_q1141 AND symb_decoder(16#37#)) OR
 					(reg_q1141 AND symb_decoder(16#34#)) OR
 					(reg_q1141 AND symb_decoder(16#35#)) OR
 					(reg_q1141 AND symb_decoder(16#36#)) OR
 					(reg_q1141 AND symb_decoder(16#38#)) OR
 					(reg_q1141 AND symb_decoder(16#30#)) OR
 					(reg_q1141 AND symb_decoder(16#31#)) OR
 					(reg_q1141 AND symb_decoder(16#32#)) OR
 					(reg_q1141 AND symb_decoder(16#39#)) OR
 					(reg_q1141 AND symb_decoder(16#33#));
reg_q1143_init <= '0' ;
	p_reg_q1143: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1143 <= reg_q1143_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1143 <= reg_q1143_init;
        else
          reg_q1143 <= reg_q1143_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1480_in <= (reg_q1478 AND symb_decoder(16#59#)) OR
 					(reg_q1478 AND symb_decoder(16#79#));
reg_q1480_init <= '0' ;
	p_reg_q1480: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1480 <= reg_q1480_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1480 <= reg_q1480_init;
        else
          reg_q1480 <= reg_q1480_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q638_in <= (reg_q636 AND symb_decoder(16#4c#)) OR
 					(reg_q636 AND symb_decoder(16#6c#));
reg_q638_init <= '0' ;
	p_reg_q638: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q638 <= reg_q638_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q638 <= reg_q638_init;
        else
          reg_q638 <= reg_q638_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q640_in <= (reg_q638 AND symb_decoder(16#49#)) OR
 					(reg_q638 AND symb_decoder(16#69#));
reg_q640_init <= '0' ;
	p_reg_q640: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q640 <= reg_q640_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q640 <= reg_q640_init;
        else
          reg_q640 <= reg_q640_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1179_in <= (reg_q1177 AND symb_decoder(16#4e#)) OR
 					(reg_q1177 AND symb_decoder(16#6e#));
reg_q1179_init <= '0' ;
	p_reg_q1179: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1179 <= reg_q1179_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1179 <= reg_q1179_init;
        else
          reg_q1179 <= reg_q1179_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1181_in <= (reg_q1179 AND symb_decoder(16#0a#)) OR
 					(reg_q1179 AND symb_decoder(16#0c#)) OR
 					(reg_q1179 AND symb_decoder(16#20#)) OR
 					(reg_q1179 AND symb_decoder(16#09#)) OR
 					(reg_q1179 AND symb_decoder(16#0d#)) OR
 					(reg_q1181 AND symb_decoder(16#09#)) OR
 					(reg_q1181 AND symb_decoder(16#20#)) OR
 					(reg_q1181 AND symb_decoder(16#0a#)) OR
 					(reg_q1181 AND symb_decoder(16#0d#)) OR
 					(reg_q1181 AND symb_decoder(16#0c#));
reg_q1181_init <= '0' ;
	p_reg_q1181: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1181 <= reg_q1181_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1181 <= reg_q1181_init;
        else
          reg_q1181 <= reg_q1181_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1375_in <= (reg_q1373 AND symb_decoder(16#66#)) OR
 					(reg_q1373 AND symb_decoder(16#46#));
reg_q1375_init <= '0' ;
	p_reg_q1375: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1375 <= reg_q1375_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1375 <= reg_q1375_init;
        else
          reg_q1375 <= reg_q1375_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2308_in <= (reg_q2306 AND symb_decoder(16#6c#)) OR
 					(reg_q2306 AND symb_decoder(16#4c#));
reg_q2308_init <= '0' ;
	p_reg_q2308: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2308 <= reg_q2308_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2308 <= reg_q2308_init;
        else
          reg_q2308 <= reg_q2308_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q750_in <= (reg_q750 AND symb_decoder(16#0c#)) OR
 					(reg_q750 AND symb_decoder(16#09#)) OR
 					(reg_q750 AND symb_decoder(16#0a#)) OR
 					(reg_q750 AND symb_decoder(16#20#)) OR
 					(reg_q750 AND symb_decoder(16#0d#)) OR
 					(reg_q748 AND symb_decoder(16#20#)) OR
 					(reg_q748 AND symb_decoder(16#0a#)) OR
 					(reg_q748 AND symb_decoder(16#0c#)) OR
 					(reg_q748 AND symb_decoder(16#0d#)) OR
 					(reg_q748 AND symb_decoder(16#09#));
reg_q750_init <= '0' ;
	p_reg_q750: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q750 <= reg_q750_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q750 <= reg_q750_init;
        else
          reg_q750 <= reg_q750_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1084_in <= (reg_q1084 AND symb_decoder(16#0d#)) OR
 					(reg_q1084 AND symb_decoder(16#09#)) OR
 					(reg_q1084 AND symb_decoder(16#20#)) OR
 					(reg_q1084 AND symb_decoder(16#0c#)) OR
 					(reg_q1084 AND symb_decoder(16#0a#)) OR
 					(reg_q1082 AND symb_decoder(16#09#)) OR
 					(reg_q1082 AND symb_decoder(16#0a#)) OR
 					(reg_q1082 AND symb_decoder(16#20#)) OR
 					(reg_q1082 AND symb_decoder(16#0c#)) OR
 					(reg_q1082 AND symb_decoder(16#0d#));
reg_q1084_init <= '0' ;
	p_reg_q1084: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1084 <= reg_q1084_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1084 <= reg_q1084_init;
        else
          reg_q1084 <= reg_q1084_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q333_in <= (reg_q331 AND symb_decoder(16#74#)) OR
 					(reg_q331 AND symb_decoder(16#54#));
reg_q333_init <= '0' ;
	p_reg_q333: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q333 <= reg_q333_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q333 <= reg_q333_init;
        else
          reg_q333 <= reg_q333_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q335_in <= (reg_q333 AND symb_decoder(16#43#)) OR
 					(reg_q333 AND symb_decoder(16#63#));
reg_q335_init <= '0' ;
	p_reg_q335: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q335 <= reg_q335_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q335 <= reg_q335_init;
        else
          reg_q335 <= reg_q335_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2288_in <= (reg_q2286 AND symb_decoder(16#0d#)) OR
 					(reg_q2286 AND symb_decoder(16#0c#)) OR
 					(reg_q2286 AND symb_decoder(16#20#)) OR
 					(reg_q2286 AND symb_decoder(16#0a#)) OR
 					(reg_q2286 AND symb_decoder(16#09#)) OR
 					(reg_q2288 AND symb_decoder(16#0a#)) OR
 					(reg_q2288 AND symb_decoder(16#0c#)) OR
 					(reg_q2288 AND symb_decoder(16#09#)) OR
 					(reg_q2288 AND symb_decoder(16#20#)) OR
 					(reg_q2288 AND symb_decoder(16#0d#));
reg_q2288_init <= '0' ;
	p_reg_q2288: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2288 <= reg_q2288_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2288 <= reg_q2288_init;
        else
          reg_q2288 <= reg_q2288_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q6_in <= (reg_q4 AND symb_decoder(16#30#));
reg_q6_init <= '0' ;
	p_reg_q6: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q6 <= reg_q6_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q6 <= reg_q6_init;
        else
          reg_q6 <= reg_q6_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q8_in <= (reg_q6 AND symb_decoder(16#46#)) OR
 					(reg_q6 AND symb_decoder(16#66#));
reg_q8_init <= '0' ;
	p_reg_q8: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q8 <= reg_q8_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q8 <= reg_q8_init;
        else
          reg_q8 <= reg_q8_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1560_in <= (reg_q1558 AND symb_decoder(16#76#)) OR
 					(reg_q1558 AND symb_decoder(16#56#));
reg_q1560_init <= '0' ;
	p_reg_q1560: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1560 <= reg_q1560_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1560 <= reg_q1560_init;
        else
          reg_q1560 <= reg_q1560_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2266_in <= (reg_q2264 AND symb_decoder(16#49#)) OR
 					(reg_q2264 AND symb_decoder(16#69#));
reg_q2266_init <= '0' ;
	p_reg_q2266: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2266 <= reg_q2266_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2266 <= reg_q2266_init;
        else
          reg_q2266 <= reg_q2266_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1141_in <= (reg_q1139 AND symb_decoder(16#2e#));
reg_q1141_init <= '0' ;
	p_reg_q1141: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1141 <= reg_q1141_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1141 <= reg_q1141_init;
        else
          reg_q1141 <= reg_q1141_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q329_in <= (reg_q327 AND symb_decoder(16#6e#)) OR
 					(reg_q327 AND symb_decoder(16#4e#));
reg_q329_init <= '0' ;
	p_reg_q329: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q329 <= reg_q329_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q329 <= reg_q329_init;
        else
          reg_q329 <= reg_q329_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q331_in <= (reg_q329 AND symb_decoder(16#65#)) OR
 					(reg_q329 AND symb_decoder(16#45#));
reg_q331_init <= '0' ;
	p_reg_q331: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q331 <= reg_q331_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q331 <= reg_q331_init;
        else
          reg_q331 <= reg_q331_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1488_in <= (reg_q1486 AND symb_decoder(16#3e#));
reg_q1488_init <= '0' ;
	p_reg_q1488: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1488 <= reg_q1488_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1488 <= reg_q1488_init;
        else
          reg_q1488 <= reg_q1488_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1337_in <= (reg_q1335 AND symb_decoder(16#2e#));
reg_q1337_init <= '0' ;
	p_reg_q1337: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1337 <= reg_q1337_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1337 <= reg_q1337_init;
        else
          reg_q1337 <= reg_q1337_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2274_in <= (reg_q2272 AND symb_decoder(16#52#)) OR
 					(reg_q2272 AND symb_decoder(16#72#));
reg_q2274_init <= '0' ;
	p_reg_q2274: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2274 <= reg_q2274_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2274 <= reg_q2274_init;
        else
          reg_q2274 <= reg_q2274_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1706_in <= (reg_q1704 AND symb_decoder(16#64#)) OR
 					(reg_q1704 AND symb_decoder(16#44#));
reg_q1706_init <= '0' ;
	p_reg_q1706: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1706 <= reg_q1706_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1706 <= reg_q1706_init;
        else
          reg_q1706 <= reg_q1706_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1708_in <= (reg_q1706 AND symb_decoder(16#0c#)) OR
 					(reg_q1706 AND symb_decoder(16#0d#)) OR
 					(reg_q1706 AND symb_decoder(16#20#)) OR
 					(reg_q1706 AND symb_decoder(16#0a#)) OR
 					(reg_q1706 AND symb_decoder(16#09#)) OR
 					(reg_q1708 AND symb_decoder(16#0d#)) OR
 					(reg_q1708 AND symb_decoder(16#0c#)) OR
 					(reg_q1708 AND symb_decoder(16#09#)) OR
 					(reg_q1708 AND symb_decoder(16#0a#)) OR
 					(reg_q1708 AND symb_decoder(16#20#));
reg_q1708_init <= '0' ;
	p_reg_q1708: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1708 <= reg_q1708_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1708 <= reg_q1708_init;
        else
          reg_q1708 <= reg_q1708_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1946_in <= (reg_q1944 AND symb_decoder(16#57#)) OR
 					(reg_q1944 AND symb_decoder(16#77#));
reg_q1946_init <= '0' ;
	p_reg_q1946: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1946 <= reg_q1946_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1946 <= reg_q1946_init;
        else
          reg_q1946 <= reg_q1946_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2435_in <= (reg_q2433 AND symb_decoder(16#45#)) OR
 					(reg_q2433 AND symb_decoder(16#65#));
reg_q2435_init <= '0' ;
	p_reg_q2435: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2435 <= reg_q2435_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2435 <= reg_q2435_init;
        else
          reg_q2435 <= reg_q2435_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2437_in <= (reg_q2435 AND symb_decoder(16#43#)) OR
 					(reg_q2435 AND symb_decoder(16#63#));
reg_q2437_init <= '0' ;
	p_reg_q2437: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2437 <= reg_q2437_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2437 <= reg_q2437_init;
        else
          reg_q2437 <= reg_q2437_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1464_in <= (reg_q1462 AND symb_decoder(16#41#)) OR
 					(reg_q1462 AND symb_decoder(16#61#));
reg_q1464_init <= '0' ;
	p_reg_q1464: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1464 <= reg_q1464_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1464 <= reg_q1464_init;
        else
          reg_q1464 <= reg_q1464_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1082_in <= (reg_q1080 AND symb_decoder(16#72#)) OR
 					(reg_q1080 AND symb_decoder(16#52#));
reg_q1082_init <= '0' ;
	p_reg_q1082: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1082 <= reg_q1082_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1082 <= reg_q1082_init;
        else
          reg_q1082 <= reg_q1082_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q770_in <= (reg_q768 AND symb_decoder(16#4f#)) OR
 					(reg_q768 AND symb_decoder(16#6f#));
reg_q770_init <= '0' ;
	p_reg_q770: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q770 <= reg_q770_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q770 <= reg_q770_init;
        else
          reg_q770 <= reg_q770_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1439_in <= (reg_q1437 AND symb_decoder(16#73#)) OR
 					(reg_q1437 AND symb_decoder(16#53#));
reg_q1439_init <= '0' ;
	p_reg_q1439: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1439 <= reg_q1439_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1439 <= reg_q1439_init;
        else
          reg_q1439 <= reg_q1439_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1744_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q1742 AND symb_decoder(16#09#)) OR
 					(reg_q1742 AND symb_decoder(16#20#)) OR
 					(reg_q1742 AND symb_decoder(16#0d#)) OR
 					(reg_q1742 AND symb_decoder(16#0a#)) OR
 					(reg_q1742 AND symb_decoder(16#0c#));
reg_q1744_init <= '0' ;
	p_reg_q1744: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1744 <= reg_q1744_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1744 <= reg_q1744_init;
        else
          reg_q1744 <= reg_q1744_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1598_in <= (reg_q1596 AND symb_decoder(16#65#)) OR
 					(reg_q1596 AND symb_decoder(16#45#));
reg_q1598_init <= '0' ;
	p_reg_q1598: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1598 <= reg_q1598_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1598 <= reg_q1598_init;
        else
          reg_q1598 <= reg_q1598_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1600_in <= (reg_q1598 AND symb_decoder(16#3a#));
reg_q1600_init <= '0' ;
	p_reg_q1600: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1600 <= reg_q1600_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1600 <= reg_q1600_init;
        else
          reg_q1600 <= reg_q1600_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1323_in <= (reg_q1321 AND symb_decoder(16#65#)) OR
 					(reg_q1321 AND symb_decoder(16#45#));
reg_q1323_init <= '0' ;
	p_reg_q1323: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1323 <= reg_q1323_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1323 <= reg_q1323_init;
        else
          reg_q1323 <= reg_q1323_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1325_in <= (reg_q1323 AND symb_decoder(16#52#)) OR
 					(reg_q1323 AND symb_decoder(16#72#));
reg_q1325_init <= '0' ;
	p_reg_q1325: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1325 <= reg_q1325_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1325 <= reg_q1325_init;
        else
          reg_q1325 <= reg_q1325_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1298_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1297 AND symb_decoder(16#0d#)) OR
 					(reg_q1297 AND symb_decoder(16#0a#));
reg_q1298_init <= '0' ;
	p_reg_q1298: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1298 <= reg_q1298_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1298 <= reg_q1298_init;
        else
          reg_q1298 <= reg_q1298_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2138_in <= (reg_q2138 AND symb_decoder(16#09#)) OR
 					(reg_q2138 AND symb_decoder(16#0c#)) OR
 					(reg_q2138 AND symb_decoder(16#0a#)) OR
 					(reg_q2138 AND symb_decoder(16#0d#)) OR
 					(reg_q2138 AND symb_decoder(16#20#)) OR
 					(reg_q2136 AND symb_decoder(16#0c#)) OR
 					(reg_q2136 AND symb_decoder(16#09#)) OR
 					(reg_q2136 AND symb_decoder(16#20#)) OR
 					(reg_q2136 AND symb_decoder(16#0d#)) OR
 					(reg_q2136 AND symb_decoder(16#0a#));
reg_q2138_init <= '0' ;
	p_reg_q2138: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2138 <= reg_q2138_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2138 <= reg_q2138_init;
        else
          reg_q2138 <= reg_q2138_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2140_in <= (reg_q2138 AND symb_decoder(16#54#)) OR
 					(reg_q2138 AND symb_decoder(16#74#));
reg_q2140_init <= '0' ;
	p_reg_q2140: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2140 <= reg_q2140_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2140 <= reg_q2140_init;
        else
          reg_q2140 <= reg_q2140_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q161_in <= (reg_q159 AND symb_decoder(16#73#)) OR
 					(reg_q159 AND symb_decoder(16#53#));
reg_q161_init <= '0' ;
	p_reg_q161: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q161 <= reg_q161_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q161 <= reg_q161_init;
        else
          reg_q161 <= reg_q161_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q163_in <= (reg_q161 AND symb_decoder(16#73#)) OR
 					(reg_q161 AND symb_decoder(16#53#));
reg_q163_init <= '0' ;
	p_reg_q163: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q163 <= reg_q163_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q163 <= reg_q163_init;
        else
          reg_q163 <= reg_q163_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2294_in <= (reg_q2292 AND symb_decoder(16#52#)) OR
 					(reg_q2292 AND symb_decoder(16#72#));
reg_q2294_init <= '0' ;
	p_reg_q2294: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2294 <= reg_q2294_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2294 <= reg_q2294_init;
        else
          reg_q2294 <= reg_q2294_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1367_in <= (reg_q1365 AND symb_decoder(16#65#)) OR
 					(reg_q1365 AND symb_decoder(16#45#));
reg_q1367_init <= '0' ;
	p_reg_q1367: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1367 <= reg_q1367_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1367 <= reg_q1367_init;
        else
          reg_q1367 <= reg_q1367_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1748_in <= (reg_q1746 AND symb_decoder(16#0a#)) OR
 					(reg_q1746 AND symb_decoder(16#0d#)) OR
 					(reg_q1746 AND symb_decoder(16#20#)) OR
 					(reg_q1746 AND symb_decoder(16#09#)) OR
 					(reg_q1746 AND symb_decoder(16#0c#));
reg_q1748_init <= '0' ;
	p_reg_q1748: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1748 <= reg_q1748_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1748 <= reg_q1748_init;
        else
          reg_q1748 <= reg_q1748_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2284_in <= (reg_q2282 AND symb_decoder(16#2e#));
reg_q2284_init <= '0' ;
	p_reg_q2284: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2284 <= reg_q2284_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2284 <= reg_q2284_init;
        else
          reg_q2284 <= reg_q2284_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q68_in <= (reg_q66 AND symb_decoder(16#45#)) OR
 					(reg_q66 AND symb_decoder(16#65#));
reg_q68_init <= '0' ;
	p_reg_q68: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q68 <= reg_q68_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q68 <= reg_q68_init;
        else
          reg_q68 <= reg_q68_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2329_in <= (reg_q2327 AND symb_decoder(16#4f#)) OR
 					(reg_q2327 AND symb_decoder(16#6f#));
reg_q2329_init <= '0' ;
	p_reg_q2329: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2329 <= reg_q2329_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2329 <= reg_q2329_init;
        else
          reg_q2329 <= reg_q2329_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2331_in <= (reg_q2329 AND symb_decoder(16#6c#)) OR
 					(reg_q2329 AND symb_decoder(16#4c#));
reg_q2331_init <= '0' ;
	p_reg_q2331: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2331 <= reg_q2331_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2331 <= reg_q2331_init;
        else
          reg_q2331 <= reg_q2331_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q984_in <= (reg_q982 AND symb_decoder(16#6f#)) OR
 					(reg_q982 AND symb_decoder(16#4f#));
reg_q984_init <= '0' ;
	p_reg_q984: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q984 <= reg_q984_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q984 <= reg_q984_init;
        else
          reg_q984 <= reg_q984_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q60_in <= (reg_q58 AND symb_decoder(16#65#)) OR
 					(reg_q58 AND symb_decoder(16#45#));
reg_q60_init <= '0' ;
	p_reg_q60: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q60 <= reg_q60_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q60 <= reg_q60_init;
        else
          reg_q60 <= reg_q60_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1692_in <= (reg_q1692 AND symb_decoder(16#20#)) OR
 					(reg_q1692 AND symb_decoder(16#09#)) OR
 					(reg_q1692 AND symb_decoder(16#0a#)) OR
 					(reg_q1692 AND symb_decoder(16#0d#)) OR
 					(reg_q1692 AND symb_decoder(16#0c#)) OR
 					(reg_q1690 AND symb_decoder(16#0d#)) OR
 					(reg_q1690 AND symb_decoder(16#20#)) OR
 					(reg_q1690 AND symb_decoder(16#0c#)) OR
 					(reg_q1690 AND symb_decoder(16#09#)) OR
 					(reg_q1690 AND symb_decoder(16#0a#));
reg_q1692_init <= '0' ;
	p_reg_q1692: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1692 <= reg_q1692_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1692 <= reg_q1692_init;
        else
          reg_q1692 <= reg_q1692_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q62_in <= (reg_q60 AND symb_decoder(16#43#)) OR
 					(reg_q60 AND symb_decoder(16#63#));
reg_q62_init <= '0' ;
	p_reg_q62: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q62 <= reg_q62_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q62 <= reg_q62_init;
        else
          reg_q62 <= reg_q62_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q395_in <= (reg_q393 AND symb_decoder(16#22#));
reg_q395_init <= '0' ;
	p_reg_q395: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q395 <= reg_q395_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q395 <= reg_q395_init;
        else
          reg_q395 <= reg_q395_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1688_in <= (reg_q1686 AND symb_decoder(16#6c#)) OR
 					(reg_q1686 AND symb_decoder(16#4c#));
reg_q1688_init <= '0' ;
	p_reg_q1688: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1688 <= reg_q1688_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1688 <= reg_q1688_init;
        else
          reg_q1688 <= reg_q1688_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1690_in <= (reg_q1688 AND symb_decoder(16#6c#)) OR
 					(reg_q1688 AND symb_decoder(16#4c#));
reg_q1690_init <= '0' ;
	p_reg_q1690: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1690 <= reg_q1690_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1690 <= reg_q1690_init;
        else
          reg_q1690 <= reg_q1690_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2134_in <= (reg_q2132 AND symb_decoder(16#4f#)) OR
 					(reg_q2132 AND symb_decoder(16#6f#));
reg_q2134_init <= '0' ;
	p_reg_q2134: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2134 <= reg_q2134_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2134 <= reg_q2134_init;
        else
          reg_q2134 <= reg_q2134_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2136_in <= (reg_q2134 AND symb_decoder(16#74#)) OR
 					(reg_q2134 AND symb_decoder(16#54#));
reg_q2136_init <= '0' ;
	p_reg_q2136: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2136 <= reg_q2136_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2136 <= reg_q2136_init;
        else
          reg_q2136 <= reg_q2136_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1910_in <= (reg_q1908 AND symb_decoder(16#6d#)) OR
 					(reg_q1908 AND symb_decoder(16#4d#));
reg_q1910_init <= '0' ;
	p_reg_q1910: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1910 <= reg_q1910_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1910 <= reg_q1910_init;
        else
          reg_q1910 <= reg_q1910_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1492_in <= (reg_q1490 AND symb_decoder(16#53#)) OR
 					(reg_q1490 AND symb_decoder(16#73#));
reg_q1492_init <= '0' ;
	p_reg_q1492: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1492 <= reg_q1492_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1492 <= reg_q1492_init;
        else
          reg_q1492 <= reg_q1492_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2117_in <= (reg_q2115 AND symb_decoder(16#6e#)) OR
 					(reg_q2115 AND symb_decoder(16#4e#));
reg_q2117_init <= '0' ;
	p_reg_q2117: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2117 <= reg_q2117_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2117 <= reg_q2117_init;
        else
          reg_q2117 <= reg_q2117_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2650_in <= (reg_q2648 AND symb_decoder(16#3a#));
reg_q2650_init <= '0' ;
	p_reg_q2650: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2650 <= reg_q2650_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2650 <= reg_q2650_init;
        else
          reg_q2650 <= reg_q2650_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q675_in <= (reg_q673 AND symb_decoder(16#3a#));
reg_q675_init <= '0' ;
	p_reg_q675: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q675 <= reg_q675_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q675 <= reg_q675_init;
        else
          reg_q675 <= reg_q675_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1531_in <= (reg_q1529 AND symb_decoder(16#75#)) OR
 					(reg_q1529 AND symb_decoder(16#55#));
reg_q1531_init <= '0' ;
	p_reg_q1531: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1531 <= reg_q1531_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1531 <= reg_q1531_init;
        else
          reg_q1531 <= reg_q1531_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1900_in <= (reg_q1898 AND symb_decoder(16#45#)) OR
 					(reg_q1898 AND symb_decoder(16#65#));
reg_q1900_init <= '0' ;
	p_reg_q1900: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1900 <= reg_q1900_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1900 <= reg_q1900_init;
        else
          reg_q1900 <= reg_q1900_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1411_in <= (reg_q1409 AND symb_decoder(16#4b#)) OR
 					(reg_q1409 AND symb_decoder(16#6b#));
reg_q1411_init <= '0' ;
	p_reg_q1411: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1411 <= reg_q1411_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1411 <= reg_q1411_init;
        else
          reg_q1411 <= reg_q1411_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1413_in <= (reg_q1411 AND symb_decoder(16#59#)) OR
 					(reg_q1411 AND symb_decoder(16#79#));
reg_q1413_init <= '0' ;
	p_reg_q1413: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1413 <= reg_q1413_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1413 <= reg_q1413_init;
        else
          reg_q1413 <= reg_q1413_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q105_in <= (reg_q103 AND symb_decoder(16#74#)) OR
 					(reg_q103 AND symb_decoder(16#54#));
reg_q105_init <= '0' ;
	p_reg_q105: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q105 <= reg_q105_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q105 <= reg_q105_init;
        else
          reg_q105 <= reg_q105_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q159_in <= (reg_q157 AND symb_decoder(16#65#)) OR
 					(reg_q157 AND symb_decoder(16#45#));
reg_q159_init <= '0' ;
	p_reg_q159: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q159 <= reg_q159_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q159 <= reg_q159_init;
        else
          reg_q159 <= reg_q159_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2107_in <= (reg_q2105 AND symb_decoder(16#48#)) OR
 					(reg_q2105 AND symb_decoder(16#68#));
reg_q2107_init <= '0' ;
	p_reg_q2107: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2107 <= reg_q2107_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2107 <= reg_q2107_init;
        else
          reg_q2107 <= reg_q2107_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1936_in <= (reg_q1934 AND symb_decoder(16#64#)) OR
 					(reg_q1934 AND symb_decoder(16#44#));
reg_q1936_init <= '0' ;
	p_reg_q1936: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1936 <= reg_q1936_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1936 <= reg_q1936_init;
        else
          reg_q1936 <= reg_q1936_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1676_in <= (reg_q1674 AND symb_decoder(16#66#)) OR
 					(reg_q1674 AND symb_decoder(16#46#));
reg_q1676_init <= '0' ;
	p_reg_q1676: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1676 <= reg_q1676_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1676 <= reg_q1676_init;
        else
          reg_q1676 <= reg_q1676_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1678_in <= (reg_q1676 AND symb_decoder(16#49#)) OR
 					(reg_q1676 AND symb_decoder(16#69#));
reg_q1678_init <= '0' ;
	p_reg_q1678: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1678 <= reg_q1678_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1678 <= reg_q1678_init;
        else
          reg_q1678 <= reg_q1678_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1502_in <= (reg_q1500 AND symb_decoder(16#52#)) OR
 					(reg_q1500 AND symb_decoder(16#72#));
reg_q1502_init <= '0' ;
	p_reg_q1502: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1502 <= reg_q1502_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1502 <= reg_q1502_init;
        else
          reg_q1502 <= reg_q1502_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1768_in <= (reg_q1766 AND symb_decoder(16#0a#)) OR
 					(reg_q1766 AND symb_decoder(16#09#)) OR
 					(reg_q1766 AND symb_decoder(16#20#)) OR
 					(reg_q1766 AND symb_decoder(16#0d#)) OR
 					(reg_q1766 AND symb_decoder(16#0c#));
reg_q1768_init <= '0' ;
	p_reg_q1768: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1768 <= reg_q1768_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1768 <= reg_q1768_init;
        else
          reg_q1768 <= reg_q1768_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q202_in <= (reg_q200 AND symb_decoder(16#53#)) OR
 					(reg_q200 AND symb_decoder(16#73#));
reg_q202_init <= '0' ;
	p_reg_q202: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q202 <= reg_q202_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q202 <= reg_q202_init;
        else
          reg_q202 <= reg_q202_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2510_in <= (reg_q2508 AND symb_decoder(16#54#));
reg_q2510_init <= '0' ;
	p_reg_q2510: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2510 <= reg_q2510_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2510 <= reg_q2510_init;
        else
          reg_q2510 <= reg_q2510_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2512_in <= (reg_q2510 AND symb_decoder(16#33#));
reg_q2512_init <= '0' ;
	p_reg_q2512: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2512 <= reg_q2512_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2512 <= reg_q2512_init;
        else
          reg_q2512 <= reg_q2512_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1527_in <= (reg_q1525 AND symb_decoder(16#74#)) OR
 					(reg_q1525 AND symb_decoder(16#54#));
reg_q1527_init <= '0' ;
	p_reg_q1527: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1527 <= reg_q1527_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1527 <= reg_q1527_init;
        else
          reg_q1527 <= reg_q1527_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1529_in <= (reg_q1527 AND symb_decoder(16#42#)) OR
 					(reg_q1527 AND symb_decoder(16#62#));
reg_q1529_init <= '0' ;
	p_reg_q1529: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1529 <= reg_q1529_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1529 <= reg_q1529_init;
        else
          reg_q1529 <= reg_q1529_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1496_in <= (reg_q1494 AND symb_decoder(16#72#)) OR
 					(reg_q1494 AND symb_decoder(16#52#));
reg_q1496_init <= '0' ;
	p_reg_q1496: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1496 <= reg_q1496_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1496 <= reg_q1496_init;
        else
          reg_q1496 <= reg_q1496_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2312_in <= (reg_q2310 AND symb_decoder(16#4e#)) OR
 					(reg_q2310 AND symb_decoder(16#6e#));
reg_q2312_init <= '0' ;
	p_reg_q2312: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2312 <= reg_q2312_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2312 <= reg_q2312_init;
        else
          reg_q2312 <= reg_q2312_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2314_in <= (reg_q2312 AND symb_decoder(16#65#)) OR
 					(reg_q2312 AND symb_decoder(16#45#));
reg_q2314_init <= '0' ;
	p_reg_q2314: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2314 <= reg_q2314_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2314 <= reg_q2314_init;
        else
          reg_q2314 <= reg_q2314_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1456_in <= (reg_q1454 AND symb_decoder(16#72#)) OR
 					(reg_q1454 AND symb_decoder(16#52#));
reg_q1456_init <= '0' ;
	p_reg_q1456: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1456 <= reg_q1456_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1456 <= reg_q1456_init;
        else
          reg_q1456 <= reg_q1456_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2692_in <= (reg_q2690 AND symb_decoder(16#21#));
reg_q2692_init <= '0' ;
	p_reg_q2692: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2692 <= reg_q2692_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2692 <= reg_q2692_init;
        else
          reg_q2692 <= reg_q2692_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2693_in <= (reg_q2692 AND symb_decoder(16#0d#));
reg_q2693_init <= '0' ;
	p_reg_q2693: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2693 <= reg_q2693_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2693 <= reg_q2693_init;
        else
          reg_q2693 <= reg_q2693_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q18_in <= (reg_q16 AND symb_decoder(16#49#)) OR
 					(reg_q16 AND symb_decoder(16#69#));
reg_q18_init <= '0' ;
	p_reg_q18: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q18 <= reg_q18_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q18 <= reg_q18_init;
        else
          reg_q18 <= reg_q18_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q959_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q958 AND symb_decoder(16#0d#)) OR
 					(reg_q958 AND symb_decoder(16#0a#));
reg_q959_init <= '0' ;
	p_reg_q959: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q959 <= reg_q959_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q959 <= reg_q959_init;
        else
          reg_q959 <= reg_q959_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q377_in <= (reg_q375 AND symb_decoder(16#68#)) OR
 					(reg_q375 AND symb_decoder(16#48#));
reg_q377_init <= '0' ;
	p_reg_q377: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q377 <= reg_q377_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q377 <= reg_q377_init;
        else
          reg_q377 <= reg_q377_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2597_in <= (reg_q2595 AND symb_decoder(16#6e#)) OR
 					(reg_q2595 AND symb_decoder(16#4e#));
reg_q2597_init <= '0' ;
	p_reg_q2597: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2597 <= reg_q2597_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2597 <= reg_q2597_init;
        else
          reg_q2597 <= reg_q2597_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q903_in <= (reg_q901 AND symb_decoder(16#0d#));
reg_q903_init <= '0' ;
	p_reg_q903: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q903 <= reg_q903_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q903 <= reg_q903_init;
        else
          reg_q903 <= reg_q903_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q905_in <= (reg_q903 AND symb_decoder(16#61#)) OR
 					(reg_q903 AND symb_decoder(16#41#));
reg_q905_init <= '0' ;
	p_reg_q905: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q905 <= reg_q905_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q905 <= reg_q905_init;
        else
          reg_q905 <= reg_q905_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1415_in <= (reg_q1413 AND symb_decoder(16#0d#));
reg_q1415_init <= '0' ;
	p_reg_q1415: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1415 <= reg_q1415_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1415 <= reg_q1415_init;
        else
          reg_q1415 <= reg_q1415_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1417_in <= (reg_q1415 AND symb_decoder(16#0a#));
reg_q1417_init <= '0' ;
	p_reg_q1417: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1417 <= reg_q1417_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1417 <= reg_q1417_init;
        else
          reg_q1417 <= reg_q1417_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2337_in <= (reg_q2335 AND symb_decoder(16#0d#)) OR
 					(reg_q2335 AND symb_decoder(16#0c#)) OR
 					(reg_q2335 AND symb_decoder(16#0a#)) OR
 					(reg_q2335 AND symb_decoder(16#09#)) OR
 					(reg_q2335 AND symb_decoder(16#20#)) OR
 					(reg_q2337 AND symb_decoder(16#20#)) OR
 					(reg_q2337 AND symb_decoder(16#0a#)) OR
 					(reg_q2337 AND symb_decoder(16#09#)) OR
 					(reg_q2337 AND symb_decoder(16#0c#)) OR
 					(reg_q2337 AND symb_decoder(16#0d#));
reg_q2337_init <= '0' ;
	p_reg_q2337: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2337 <= reg_q2337_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2337 <= reg_q2337_init;
        else
          reg_q2337 <= reg_q2337_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1151_in <= (reg_q1149 AND symb_decoder(16#0a#));
reg_q1151_init <= '0' ;
	p_reg_q1151: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1151 <= reg_q1151_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1151 <= reg_q1151_init;
        else
          reg_q1151 <= reg_q1151_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1153_in <= (reg_q1151 AND symb_decoder(16#0d#));
reg_q1153_init <= '0' ;
	p_reg_q1153: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1153 <= reg_q1153_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1153 <= reg_q1153_init;
        else
          reg_q1153 <= reg_q1153_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2662_in <= (reg_q2660 AND symb_decoder(16#6f#)) OR
 					(reg_q2660 AND symb_decoder(16#4f#));
reg_q2662_init <= '0' ;
	p_reg_q2662: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2662 <= reg_q2662_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2662 <= reg_q2662_init;
        else
          reg_q2662 <= reg_q2662_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2339_in <= (reg_q2337 AND symb_decoder(16#52#)) OR
 					(reg_q2337 AND symb_decoder(16#72#));
reg_q2339_init <= '0' ;
	p_reg_q2339: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2339 <= reg_q2339_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2339 <= reg_q2339_init;
        else
          reg_q2339 <= reg_q2339_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q705_in <= (reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q704 AND symb_decoder(16#43#)) OR
 					(reg_q704 AND symb_decoder(16#63#));
reg_q705_init <= '0' ;
	p_reg_q705: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q705 <= reg_q705_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q705 <= reg_q705_init;
        else
          reg_q705 <= reg_q705_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2345_in <= (reg_q2343 AND symb_decoder(16#4f#)) OR
 					(reg_q2343 AND symb_decoder(16#6f#));
reg_q2345_init <= '0' ;
	p_reg_q2345: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2345 <= reg_q2345_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2345 <= reg_q2345_init;
        else
          reg_q2345 <= reg_q2345_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1548_in <= (reg_q1546 AND symb_decoder(16#45#)) OR
 					(reg_q1546 AND symb_decoder(16#65#));
reg_q1548_init <= '0' ;
	p_reg_q1548: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1548 <= reg_q1548_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1548 <= reg_q1548_init;
        else
          reg_q1548 <= reg_q1548_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q337_in <= (reg_q335 AND symb_decoder(16#6f#)) OR
 					(reg_q335 AND symb_decoder(16#4f#));
reg_q337_init <= '0' ;
	p_reg_q337: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q337 <= reg_q337_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q337 <= reg_q337_init;
        else
          reg_q337 <= reg_q337_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q476_in <= (reg_q474 AND symb_decoder(16#30#));
reg_q476_init <= '0' ;
	p_reg_q476: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q476 <= reg_q476_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q476 <= reg_q476_init;
        else
          reg_q476 <= reg_q476_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1478_in <= (reg_q1476 AND symb_decoder(16#64#)) OR
 					(reg_q1476 AND symb_decoder(16#44#));
reg_q1478_init <= '0' ;
	p_reg_q1478: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1478 <= reg_q1478_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1478 <= reg_q1478_init;
        else
          reg_q1478 <= reg_q1478_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2272_in <= (reg_q2270 AND symb_decoder(16#50#)) OR
 					(reg_q2270 AND symb_decoder(16#70#));
reg_q2272_init <= '0' ;
	p_reg_q2272: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2272 <= reg_q2272_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2272 <= reg_q2272_init;
        else
          reg_q2272 <= reg_q2272_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1656_in <= (reg_q1654 AND symb_decoder(16#36#));
reg_q1656_init <= '0' ;
	p_reg_q1656: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1656 <= reg_q1656_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1656 <= reg_q1656_init;
        else
          reg_q1656 <= reg_q1656_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1658_in <= (reg_q1656 AND symb_decoder(16#36#));
reg_q1658_init <= '0' ;
	p_reg_q1658: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1658 <= reg_q1658_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1658 <= reg_q1658_init;
        else
          reg_q1658 <= reg_q1658_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q842_in <= (reg_q840 AND symb_decoder(16#2e#));
reg_q842_init <= '0' ;
	p_reg_q842: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q842 <= reg_q842_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q842 <= reg_q842_init;
        else
          reg_q842 <= reg_q842_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1321_in <= (reg_q1319 AND symb_decoder(16#73#)) OR
 					(reg_q1319 AND symb_decoder(16#53#));
reg_q1321_init <= '0' ;
	p_reg_q1321: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1321 <= reg_q1321_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1321 <= reg_q1321_init;
        else
          reg_q1321 <= reg_q1321_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1004_in <= (reg_q1002 AND symb_decoder(16#3a#));
reg_q1004_init <= '0' ;
	p_reg_q1004: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1004 <= reg_q1004_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1004 <= reg_q1004_init;
        else
          reg_q1004 <= reg_q1004_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q594_in <= (reg_q592 AND symb_decoder(16#58#)) OR
 					(reg_q592 AND symb_decoder(16#78#));
reg_q594_init <= '0' ;
	p_reg_q594: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q594 <= reg_q594_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q594 <= reg_q594_init;
        else
          reg_q594 <= reg_q594_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1051_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1050 AND symb_decoder(16#0d#)) OR
 					(reg_q1050 AND symb_decoder(16#0a#));
reg_q1051_init <= '0' ;
	p_reg_q1051: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1051 <= reg_q1051_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1051 <= reg_q1051_init;
        else
          reg_q1051 <= reg_q1051_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2196_in <= (reg_q2194 AND symb_decoder(16#64#)) OR
 					(reg_q2194 AND symb_decoder(16#44#));
reg_q2196_init <= '0' ;
	p_reg_q2196: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2196 <= reg_q2196_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2196 <= reg_q2196_init;
        else
          reg_q2196 <= reg_q2196_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2198_in <= (reg_q2196 AND symb_decoder(16#41#)) OR
 					(reg_q2196 AND symb_decoder(16#61#));
reg_q2198_init <= '0' ;
	p_reg_q2198: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2198 <= reg_q2198_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2198 <= reg_q2198_init;
        else
          reg_q2198 <= reg_q2198_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2231_in <= (reg_q2229 AND symb_decoder(16#73#)) OR
 					(reg_q2229 AND symb_decoder(16#53#));
reg_q2231_init <= '0' ;
	p_reg_q2231: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2231 <= reg_q2231_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2231 <= reg_q2231_init;
        else
          reg_q2231 <= reg_q2231_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2455_in <= (reg_q2453 AND symb_decoder(16#23#));
reg_q2455_init <= '0' ;
	p_reg_q2455: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2455 <= reg_q2455_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2455 <= reg_q2455_init;
        else
          reg_q2455 <= reg_q2455_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2457_in <= (reg_q2455 AND symb_decoder(16#33#));
reg_q2457_init <= '0' ;
	p_reg_q2457: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2457 <= reg_q2457_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2457 <= reg_q2457_init;
        else
          reg_q2457 <= reg_q2457_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q748_in <= (reg_q746 AND symb_decoder(16#54#)) OR
 					(reg_q746 AND symb_decoder(16#74#));
reg_q748_init <= '0' ;
	p_reg_q748: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q748 <= reg_q748_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q748 <= reg_q748_init;
        else
          reg_q748 <= reg_q748_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2557_in <= (reg_q2555 AND symb_decoder(16#45#)) OR
 					(reg_q2555 AND symb_decoder(16#65#));
reg_q2557_init <= '0' ;
	p_reg_q2557: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2557 <= reg_q2557_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2557 <= reg_q2557_init;
        else
          reg_q2557 <= reg_q2557_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2559_in <= (reg_q2557 AND symb_decoder(16#52#)) OR
 					(reg_q2557 AND symb_decoder(16#72#));
reg_q2559_init <= '0' ;
	p_reg_q2559: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2559 <= reg_q2559_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2559 <= reg_q2559_init;
        else
          reg_q2559 <= reg_q2559_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2668_in <= (reg_q2666 AND symb_decoder(16#69#)) OR
 					(reg_q2666 AND symb_decoder(16#49#));
reg_q2668_init <= '0' ;
	p_reg_q2668: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2668 <= reg_q2668_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2668 <= reg_q2668_init;
        else
          reg_q2668 <= reg_q2668_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2670_in <= (reg_q2668 AND symb_decoder(16#6e#)) OR
 					(reg_q2668 AND symb_decoder(16#4e#));
reg_q2670_init <= '0' ;
	p_reg_q2670: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2670 <= reg_q2670_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2670 <= reg_q2670_init;
        else
          reg_q2670 <= reg_q2670_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2310_in <= (reg_q2308 AND symb_decoder(16#49#)) OR
 					(reg_q2308 AND symb_decoder(16#69#));
reg_q2310_init <= '0' ;
	p_reg_q2310: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2310 <= reg_q2310_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2310 <= reg_q2310_init;
        else
          reg_q2310 <= reg_q2310_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2150_in <= (reg_q2148 AND symb_decoder(16#47#)) OR
 					(reg_q2148 AND symb_decoder(16#67#));
reg_q2150_init <= '0' ;
	p_reg_q2150: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2150 <= reg_q2150_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2150 <= reg_q2150_init;
        else
          reg_q2150 <= reg_q2150_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q466_in <= (reg_q464 AND symb_decoder(16#65#)) OR
 					(reg_q464 AND symb_decoder(16#45#));
reg_q466_init <= '0' ;
	p_reg_q466: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q466 <= reg_q466_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q466 <= reg_q466_init;
        else
          reg_q466 <= reg_q466_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q468_in <= (reg_q466 AND symb_decoder(16#61#)) OR
 					(reg_q466 AND symb_decoder(16#41#));
reg_q468_init <= '0' ;
	p_reg_q468: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q468 <= reg_q468_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q468 <= reg_q468_init;
        else
          reg_q468 <= reg_q468_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q852_in <= (reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q850 AND symb_decoder(16#5b#));
reg_q852_init <= '0' ;
	p_reg_q852: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q852 <= reg_q852_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q852 <= reg_q852_init;
        else
          reg_q852 <= reg_q852_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q854_in <= (reg_q852 AND symb_decoder(16#64#)) OR
 					(reg_q852 AND symb_decoder(16#44#));
reg_q854_init <= '0' ;
	p_reg_q854: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q854 <= reg_q854_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q854 <= reg_q854_init;
        else
          reg_q854 <= reg_q854_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q415_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q414 AND symb_decoder(16#0a#)) OR
 					(reg_q414 AND symb_decoder(16#0d#));
reg_q415_init <= '0' ;
	p_reg_q415: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q415 <= reg_q415_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q415 <= reg_q415_init;
        else
          reg_q415 <= reg_q415_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q416_in <= (reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q415 AND symb_decoder(16#62#)) OR
 					(reg_q415 AND symb_decoder(16#42#));
reg_q416_init <= '0' ;
	p_reg_q416: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q416 <= reg_q416_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q416 <= reg_q416_init;
        else
          reg_q416 <= reg_q416_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1914_in <= (reg_q1912 AND symb_decoder(16#74#)) OR
 					(reg_q1912 AND symb_decoder(16#54#));
reg_q1914_init <= '0' ;
	p_reg_q1914: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1914 <= reg_q1914_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1914 <= reg_q1914_init;
        else
          reg_q1914 <= reg_q1914_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2439_in <= (reg_q2437 AND symb_decoder(16#54#)) OR
 					(reg_q2437 AND symb_decoder(16#74#));
reg_q2439_init <= '0' ;
	p_reg_q2439: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2439 <= reg_q2439_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2439 <= reg_q2439_init;
        else
          reg_q2439 <= reg_q2439_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1307_in <= (reg_q1305 AND symb_decoder(16#46#)) OR
 					(reg_q1305 AND symb_decoder(16#66#));
reg_q1307_init <= '0' ;
	p_reg_q1307: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1307 <= reg_q1307_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1307 <= reg_q1307_init;
        else
          reg_q1307 <= reg_q1307_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q628_in <= (reg_q626 AND symb_decoder(16#45#)) OR
 					(reg_q626 AND symb_decoder(16#65#));
reg_q628_init <= '0' ;
	p_reg_q628: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q628 <= reg_q628_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q628 <= reg_q628_init;
        else
          reg_q628 <= reg_q628_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2132_in <= (reg_q2130 AND symb_decoder(16#47#)) OR
 					(reg_q2130 AND symb_decoder(16#67#));
reg_q2132_init <= '0' ;
	p_reg_q2132: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2132 <= reg_q2132_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2132 <= reg_q2132_init;
        else
          reg_q2132 <= reg_q2132_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2459_in <= (reg_q2457 AND symb_decoder(16#23#));
reg_q2459_init <= '0' ;
	p_reg_q2459: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2459 <= reg_q2459_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2459 <= reg_q2459_init;
        else
          reg_q2459 <= reg_q2459_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1726_in <= (reg_q1724 AND symb_decoder(16#75#)) OR
 					(reg_q1724 AND symb_decoder(16#55#));
reg_q1726_init <= '0' ;
	p_reg_q1726: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1726 <= reg_q1726_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1726 <= reg_q1726_init;
        else
          reg_q1726 <= reg_q1726_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q538_in <= (reg_q536 AND symb_decoder(16#25#));
reg_q538_init <= '0' ;
	p_reg_q538: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q538 <= reg_q538_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q538 <= reg_q538_init;
        else
          reg_q538 <= reg_q538_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q540_in <= (reg_q538 AND symb_decoder(16#32#));
reg_q540_init <= '0' ;
	p_reg_q540: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q540 <= reg_q540_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q540 <= reg_q540_init;
        else
          reg_q540 <= reg_q540_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2583_in <= (reg_q2615 AND symb_decoder(16#0d#)) OR
 					(reg_q2579 AND symb_decoder(16#0d#));
reg_q2583_init <= '0' ;
	p_reg_q2583: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2583 <= reg_q2583_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2583 <= reg_q2583_init;
        else
          reg_q2583 <= reg_q2583_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q588_in <= (reg_q586 AND symb_decoder(16#70#)) OR
 					(reg_q586 AND symb_decoder(16#50#));
reg_q588_init <= '0' ;
	p_reg_q588: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q588 <= reg_q588_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q588 <= reg_q588_init;
        else
          reg_q588 <= reg_q588_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1684_in <= (reg_q1682 AND symb_decoder(16#57#)) OR
 					(reg_q1682 AND symb_decoder(16#77#));
reg_q1684_init <= '0' ;
	p_reg_q1684: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1684 <= reg_q1684_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1684 <= reg_q1684_init;
        else
          reg_q1684 <= reg_q1684_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1686_in <= (reg_q1684 AND symb_decoder(16#41#)) OR
 					(reg_q1684 AND symb_decoder(16#61#));
reg_q1686_init <= '0' ;
	p_reg_q1686: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1686 <= reg_q1686_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1686 <= reg_q1686_init;
        else
          reg_q1686 <= reg_q1686_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q403_in <= (reg_q401 AND symb_decoder(16#6f#)) OR
 					(reg_q401 AND symb_decoder(16#4f#));
reg_q403_init <= '0' ;
	p_reg_q403: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q403 <= reg_q403_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q403 <= reg_q403_init;
        else
          reg_q403 <= reg_q403_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q405_in <= (reg_q403 AND symb_decoder(16#4a#)) OR
 					(reg_q403 AND symb_decoder(16#6a#));
reg_q405_init <= '0' ;
	p_reg_q405: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q405 <= reg_q405_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q405 <= reg_q405_init;
        else
          reg_q405 <= reg_q405_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2347_in <= (reg_q2345 AND symb_decoder(16#74#)) OR
 					(reg_q2345 AND symb_decoder(16#54#));
reg_q2347_init <= '0' ;
	p_reg_q2347: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2347 <= reg_q2347_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2347 <= reg_q2347_init;
        else
          reg_q2347 <= reg_q2347_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q446_in <= (reg_q444 AND symb_decoder(16#72#)) OR
 					(reg_q444 AND symb_decoder(16#52#));
reg_q446_init <= '0' ;
	p_reg_q446: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q446 <= reg_q446_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q446 <= reg_q446_init;
        else
          reg_q446 <= reg_q446_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1014_in <= (reg_q1013 AND symb_decoder(16#0d#)) OR
 					(reg_q1013 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#));
reg_q1014_init <= '0' ;
	p_reg_q1014: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1014 <= reg_q1014_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1014 <= reg_q1014_init;
        else
          reg_q1014 <= reg_q1014_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q570_in <= (reg_q568 AND symb_decoder(16#32#));
reg_q570_init <= '0' ;
	p_reg_q570: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q570 <= reg_q570_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q570 <= reg_q570_init;
        else
          reg_q570 <= reg_q570_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1183_in <= (reg_q1181 AND symb_decoder(16#73#)) OR
 					(reg_q1181 AND symb_decoder(16#53#));
reg_q1183_init <= '0' ;
	p_reg_q1183: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1183 <= reg_q1183_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1183 <= reg_q1183_init;
        else
          reg_q1183 <= reg_q1183_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1185_in <= (reg_q1183 AND symb_decoder(16#54#)) OR
 					(reg_q1183 AND symb_decoder(16#74#));
reg_q1185_init <= '0' ;
	p_reg_q1185: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1185 <= reg_q1185_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1185 <= reg_q1185_init;
        else
          reg_q1185 <= reg_q1185_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q194_in <= (reg_q192 AND symb_decoder(16#47#)) OR
 					(reg_q192 AND symb_decoder(16#67#));
reg_q194_init <= '0' ;
	p_reg_q194: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q194 <= reg_q194_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q194 <= reg_q194_init;
        else
          reg_q194 <= reg_q194_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q196_in <= (reg_q194 AND symb_decoder(16#45#)) OR
 					(reg_q194 AND symb_decoder(16#65#));
reg_q196_init <= '0' ;
	p_reg_q196: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q196 <= reg_q196_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q196 <= reg_q196_init;
        else
          reg_q196 <= reg_q196_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1331_in <= (reg_q1329 AND symb_decoder(16#72#)) OR
 					(reg_q1329 AND symb_decoder(16#52#));
reg_q1331_init <= '0' ;
	p_reg_q1331: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1331 <= reg_q1331_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1331 <= reg_q1331_init;
        else
          reg_q1331 <= reg_q1331_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q294_in <= (reg_q292 AND symb_decoder(16#63#)) OR
 					(reg_q292 AND symb_decoder(16#43#));
reg_q294_init <= '0' ;
	p_reg_q294: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q294 <= reg_q294_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q294 <= reg_q294_init;
        else
          reg_q294 <= reg_q294_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q296_in <= (reg_q294 AND symb_decoder(16#4f#)) OR
 					(reg_q294 AND symb_decoder(16#6f#));
reg_q296_init <= '0' ;
	p_reg_q296: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q296 <= reg_q296_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q296 <= reg_q296_init;
        else
          reg_q296 <= reg_q296_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1615_in <= (reg_q1613 AND symb_decoder(16#46#)) OR
 					(reg_q1613 AND symb_decoder(16#66#));
reg_q1615_init <= '0' ;
	p_reg_q1615: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1615 <= reg_q1615_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1615 <= reg_q1615_init;
        else
          reg_q1615 <= reg_q1615_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1617_in <= (reg_q1615 AND symb_decoder(16#72#)) OR
 					(reg_q1615 AND symb_decoder(16#52#));
reg_q1617_init <= '0' ;
	p_reg_q1617: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1617 <= reg_q1617_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1617 <= reg_q1617_init;
        else
          reg_q1617 <= reg_q1617_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1682_in <= (reg_q1680 AND symb_decoder(16#45#)) OR
 					(reg_q1680 AND symb_decoder(16#65#));
reg_q1682_init <= '0' ;
	p_reg_q1682: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1682 <= reg_q1682_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1682 <= reg_q1682_init;
        else
          reg_q1682 <= reg_q1682_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1892_in <= (reg_q1890 AND symb_decoder(16#44#)) OR
 					(reg_q1890 AND symb_decoder(16#64#));
reg_q1892_init <= '0' ;
	p_reg_q1892: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1892 <= reg_q1892_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1892 <= reg_q1892_init;
        else
          reg_q1892 <= reg_q1892_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q502_in <= (reg_q500 AND symb_decoder(16#4e#)) OR
 					(reg_q500 AND symb_decoder(16#6e#));
reg_q502_init <= '0' ;
	p_reg_q502: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q502 <= reg_q502_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q502 <= reg_q502_init;
        else
          reg_q502 <= reg_q502_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q504_in <= (reg_q502 AND symb_decoder(16#45#)) OR
 					(reg_q502 AND symb_decoder(16#65#));
reg_q504_init <= '0' ;
	p_reg_q504: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q504 <= reg_q504_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q504 <= reg_q504_init;
        else
          reg_q504 <= reg_q504_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1957_in <= (reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q1956 AND symb_decoder(16#73#)) OR
 					(reg_q1956 AND symb_decoder(16#53#));
reg_q1957_init <= '0' ;
	p_reg_q1957: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1957 <= reg_q1957_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1957 <= reg_q1957_init;
        else
          reg_q1957 <= reg_q1957_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1959_in <= (reg_q1957 AND symb_decoder(16#69#)) OR
 					(reg_q1957 AND symb_decoder(16#49#));
reg_q1959_init <= '0' ;
	p_reg_q1959: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1959 <= reg_q1959_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1959 <= reg_q1959_init;
        else
          reg_q1959 <= reg_q1959_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1035_in <= (reg_q1035 AND symb_decoder(16#0a#)) OR
 					(reg_q1035 AND symb_decoder(16#0d#)) OR
 					(reg_q1035 AND symb_decoder(16#09#)) OR
 					(reg_q1035 AND symb_decoder(16#0c#)) OR
 					(reg_q1035 AND symb_decoder(16#20#)) OR
 					(reg_q1033 AND symb_decoder(16#0c#)) OR
 					(reg_q1033 AND symb_decoder(16#20#)) OR
 					(reg_q1033 AND symb_decoder(16#09#)) OR
 					(reg_q1033 AND symb_decoder(16#0d#)) OR
 					(reg_q1033 AND symb_decoder(16#0a#));
reg_q1035_init <= '0' ;
	p_reg_q1035: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1035 <= reg_q1035_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1035 <= reg_q1035_init;
        else
          reg_q1035 <= reg_q1035_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2425_in <= (reg_q2423 AND symb_decoder(16#41#)) OR
 					(reg_q2423 AND symb_decoder(16#61#));
reg_q2425_init <= '0' ;
	p_reg_q2425: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2425 <= reg_q2425_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2425 <= reg_q2425_init;
        else
          reg_q2425 <= reg_q2425_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1017_in <= (reg_q1015 AND symb_decoder(16#72#)) OR
 					(reg_q1015 AND symb_decoder(16#52#));
reg_q1017_init <= '0' ;
	p_reg_q1017: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1017 <= reg_q1017_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1017 <= reg_q1017_init;
        else
          reg_q1017 <= reg_q1017_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1019_in <= (reg_q1017 AND symb_decoder(16#61#)) OR
 					(reg_q1017 AND symb_decoder(16#41#));
reg_q1019_init <= '0' ;
	p_reg_q1019: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1019 <= reg_q1019_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1019 <= reg_q1019_init;
        else
          reg_q1019 <= reg_q1019_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q361_in <= (reg_q359 AND symb_decoder(16#72#)) OR
 					(reg_q359 AND symb_decoder(16#52#));
reg_q361_init <= '0' ;
	p_reg_q361: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q361 <= reg_q361_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q361 <= reg_q361_init;
        else
          reg_q361 <= reg_q361_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q141_in <= (reg_q139 AND symb_decoder(16#43#)) OR
 					(reg_q139 AND symb_decoder(16#63#));
reg_q141_init <= '0' ;
	p_reg_q141: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q141 <= reg_q141_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q141 <= reg_q141_init;
        else
          reg_q141 <= reg_q141_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q50_in <= (reg_q48 AND symb_decoder(16#30#));
reg_q50_init <= '0' ;
	p_reg_q50: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q50 <= reg_q50_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q50 <= reg_q50_init;
        else
          reg_q50 <= reg_q50_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2522_in <= (reg_q2520 AND symb_decoder(16#67#)) OR
 					(reg_q2520 AND symb_decoder(16#47#));
reg_q2522_init <= '0' ;
	p_reg_q2522: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2522 <= reg_q2522_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2522 <= reg_q2522_init;
        else
          reg_q2522 <= reg_q2522_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q586_in <= (reg_q584 AND symb_decoder(16#6f#)) OR
 					(reg_q584 AND symb_decoder(16#4f#));
reg_q586_init <= '0' ;
	p_reg_q586: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q586 <= reg_q586_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q586 <= reg_q586_init;
        else
          reg_q586 <= reg_q586_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q724_in <= (reg_q722 AND symb_decoder(16#74#)) OR
 					(reg_q722 AND symb_decoder(16#54#));
reg_q724_init <= '0' ;
	p_reg_q724: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q724 <= reg_q724_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q724 <= reg_q724_init;
        else
          reg_q724 <= reg_q724_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q968_in <= (reg_q966 AND symb_decoder(16#65#)) OR
 					(reg_q966 AND symb_decoder(16#45#));
reg_q968_init <= '0' ;
	p_reg_q968: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q968 <= reg_q968_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q968 <= reg_q968_init;
        else
          reg_q968 <= reg_q968_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q970_in <= (reg_q968 AND symb_decoder(16#4c#)) OR
 					(reg_q968 AND symb_decoder(16#6c#));
reg_q970_init <= '0' ;
	p_reg_q970: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q970 <= reg_q970_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q970 <= reg_q970_init;
        else
          reg_q970 <= reg_q970_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1023_in <= (reg_q1021 AND symb_decoder(16#45#)) OR
 					(reg_q1021 AND symb_decoder(16#65#));
reg_q1023_init <= '0' ;
	p_reg_q1023: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1023 <= reg_q1023_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1023 <= reg_q1023_init;
        else
          reg_q1023 <= reg_q1023_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1159_in <= (reg_q1157 AND symb_decoder(16#0a#));
reg_q1159_init <= '0' ;
	p_reg_q1159: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1159 <= reg_q1159_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1159 <= reg_q1159_init;
        else
          reg_q1159 <= reg_q1159_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2534_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2533 AND symb_decoder(16#0a#)) OR
 					(reg_q2533 AND symb_decoder(16#0d#));
reg_q2534_init <= '0' ;
	p_reg_q2534: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2534 <= reg_q2534_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2534 <= reg_q2534_init;
        else
          reg_q2534 <= reg_q2534_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1169_in <= (reg_q1167 AND symb_decoder(16#65#)) OR
 					(reg_q1167 AND symb_decoder(16#45#));
reg_q1169_init <= '0' ;
	p_reg_q1169: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1169 <= reg_q1169_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1169 <= reg_q1169_init;
        else
          reg_q1169 <= reg_q1169_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q349_in <= (reg_q347 AND symb_decoder(16#2e#));
reg_q349_init <= '0' ;
	p_reg_q349: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q349 <= reg_q349_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q349 <= reg_q349_init;
        else
          reg_q349 <= reg_q349_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2403_in <= (reg_q2401 AND symb_decoder(16#6f#)) OR
 					(reg_q2401 AND symb_decoder(16#4f#));
reg_q2403_init <= '0' ;
	p_reg_q2403: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2403 <= reg_q2403_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2403 <= reg_q2403_init;
        else
          reg_q2403 <= reg_q2403_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2182_in <= (reg_q2180 AND symb_decoder(16#54#)) OR
 					(reg_q2180 AND symb_decoder(16#74#));
reg_q2182_init <= '0' ;
	p_reg_q2182: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2182 <= reg_q2182_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2182 <= reg_q2182_init;
        else
          reg_q2182 <= reg_q2182_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1033_in <= (reg_q1031 AND symb_decoder(16#6e#)) OR
 					(reg_q1031 AND symb_decoder(16#4e#));
reg_q1033_init <= '0' ;
	p_reg_q1033: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1033 <= reg_q1033_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1033 <= reg_q1033_init;
        else
          reg_q1033 <= reg_q1033_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2445_in <= (reg_q2443 AND symb_decoder(16#6f#)) OR
 					(reg_q2443 AND symb_decoder(16#4f#));
reg_q2445_init <= '0' ;
	p_reg_q2445: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2445 <= reg_q2445_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2445 <= reg_q2445_init;
        else
          reg_q2445 <= reg_q2445_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2447_in <= (reg_q2445 AND symb_decoder(16#41#)) OR
 					(reg_q2445 AND symb_decoder(16#61#));
reg_q2447_init <= '0' ;
	p_reg_q2447: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2447 <= reg_q2447_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2447 <= reg_q2447_init;
        else
          reg_q2447 <= reg_q2447_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1971_in <= (reg_q1969 AND symb_decoder(16#45#)) OR
 					(reg_q1969 AND symb_decoder(16#65#));
reg_q1971_init <= '0' ;
	p_reg_q1971: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1971 <= reg_q1971_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1971 <= reg_q1971_init;
        else
          reg_q1971 <= reg_q1971_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1973_in <= (reg_q1971 AND symb_decoder(16#72#)) OR
 					(reg_q1971 AND symb_decoder(16#52#));
reg_q1973_init <= '0' ;
	p_reg_q1973: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1973 <= reg_q1973_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1973 <= reg_q1973_init;
        else
          reg_q1973 <= reg_q1973_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2640_in <= (reg_q2638 AND symb_decoder(16#72#)) OR
 					(reg_q2638 AND symb_decoder(16#52#));
reg_q2640_init <= '0' ;
	p_reg_q2640: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2640 <= reg_q2640_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2640 <= reg_q2640_init;
        else
          reg_q2640 <= reg_q2640_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q399_in <= (reg_q397 AND symb_decoder(16#50#)) OR
 					(reg_q397 AND symb_decoder(16#70#));
reg_q399_init <= '0' ;
	p_reg_q399: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q399 <= reg_q399_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q399 <= reg_q399_init;
        else
          reg_q399 <= reg_q399_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q401_in <= (reg_q399 AND symb_decoder(16#72#)) OR
 					(reg_q399 AND symb_decoder(16#52#));
reg_q401_init <= '0' ;
	p_reg_q401: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q401 <= reg_q401_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q401 <= reg_q401_init;
        else
          reg_q401 <= reg_q401_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1447_in <= (reg_q1445 AND symb_decoder(16#65#)) OR
 					(reg_q1445 AND symb_decoder(16#45#));
reg_q1447_init <= '0' ;
	p_reg_q1447: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1447 <= reg_q1447_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1447 <= reg_q1447_init;
        else
          reg_q1447 <= reg_q1447_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1449_in <= (reg_q1447 AND symb_decoder(16#6d#)) OR
 					(reg_q1447 AND symb_decoder(16#4d#));
reg_q1449_init <= '0' ;
	p_reg_q1449: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1449 <= reg_q1449_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1449 <= reg_q1449_init;
        else
          reg_q1449 <= reg_q1449_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1716_in <= (reg_q1714 AND symb_decoder(16#74#)) OR
 					(reg_q1714 AND symb_decoder(16#54#));
reg_q1716_init <= '0' ;
	p_reg_q1716: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1716 <= reg_q1716_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1716 <= reg_q1716_init;
        else
          reg_q1716 <= reg_q1716_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q580_in <= (reg_q578 AND symb_decoder(16#25#));
reg_q580_init <= '0' ;
	p_reg_q580: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q580 <= reg_q580_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q580 <= reg_q580_init;
        else
          reg_q580 <= reg_q580_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q582_in <= (reg_q580 AND symb_decoder(16#32#));
reg_q582_init <= '0' ;
	p_reg_q582: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q582 <= reg_q582_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q582 <= reg_q582_init;
        else
          reg_q582 <= reg_q582_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1710_in <= (reg_q1708 AND symb_decoder(16#50#)) OR
 					(reg_q1708 AND symb_decoder(16#70#));
reg_q1710_init <= '0' ;
	p_reg_q1710: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1710 <= reg_q1710_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1710 <= reg_q1710_init;
        else
          reg_q1710 <= reg_q1710_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2474_in <= (reg_q2472 AND symb_decoder(16#52#));
reg_q2474_init <= '0' ;
	p_reg_q2474: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2474 <= reg_q2474_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2474 <= reg_q2474_init;
        else
          reg_q2474 <= reg_q2474_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2476_in <= (reg_q2474 AND symb_decoder(16#54#));
reg_q2476_init <= '0' ;
	p_reg_q2476: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2476 <= reg_q2476_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2476 <= reg_q2476_init;
        else
          reg_q2476 <= reg_q2476_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q758_in <= (reg_q756 AND symb_decoder(16#64#)) OR
 					(reg_q756 AND symb_decoder(16#44#));
reg_q758_init <= '0' ;
	p_reg_q758: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q758 <= reg_q758_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q758 <= reg_q758_init;
        else
          reg_q758 <= reg_q758_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q760_in <= (reg_q758 AND symb_decoder(16#69#)) OR
 					(reg_q758 AND symb_decoder(16#49#));
reg_q760_init <= '0' ;
	p_reg_q760: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q760 <= reg_q760_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q760 <= reg_q760_init;
        else
          reg_q760 <= reg_q760_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q820_in <= (reg_q818 AND symb_decoder(16#6d#)) OR
 					(reg_q818 AND symb_decoder(16#4d#));
reg_q820_init <= '0' ;
	p_reg_q820: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q820 <= reg_q820_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q820 <= reg_q820_init;
        else
          reg_q820 <= reg_q820_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q822_in <= (reg_q820 AND symb_decoder(16#49#)) OR
 					(reg_q820 AND symb_decoder(16#69#));
reg_q822_init <= '0' ;
	p_reg_q822: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q822 <= reg_q822_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q822 <= reg_q822_init;
        else
          reg_q822 <= reg_q822_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2010_in <= (reg_q2008 AND symb_decoder(16#61#)) OR
 					(reg_q2008 AND symb_decoder(16#41#));
reg_q2010_init <= '0' ;
	p_reg_q2010: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2010 <= reg_q2010_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2010 <= reg_q2010_init;
        else
          reg_q2010 <= reg_q2010_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2012_in <= (reg_q2010 AND symb_decoder(16#6e#)) OR
 					(reg_q2010 AND symb_decoder(16#4e#));
reg_q2012_init <= '0' ;
	p_reg_q2012: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2012 <= reg_q2012_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2012 <= reg_q2012_init;
        else
          reg_q2012 <= reg_q2012_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q496_in <= (reg_q494 AND symb_decoder(16#6e#)) OR
 					(reg_q494 AND symb_decoder(16#4e#));
reg_q496_init <= '0' ;
	p_reg_q496: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q496 <= reg_q496_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q496 <= reg_q496_init;
        else
          reg_q496 <= reg_q496_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q498_in <= (reg_q496 AND symb_decoder(16#6c#)) OR
 					(reg_q496 AND symb_decoder(16#4c#));
reg_q498_init <= '0' ;
	p_reg_q498: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q498 <= reg_q498_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q498 <= reg_q498_init;
        else
          reg_q498 <= reg_q498_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q972_in <= (reg_q970 AND symb_decoder(16#63#)) OR
 					(reg_q970 AND symb_decoder(16#43#));
reg_q972_init <= '0' ;
	p_reg_q972: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q972 <= reg_q972_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q972 <= reg_q972_init;
        else
          reg_q972 <= reg_q972_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q730_in <= (reg_q728 AND symb_decoder(16#4e#)) OR
 					(reg_q728 AND symb_decoder(16#6e#));
reg_q730_init <= '0' ;
	p_reg_q730: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q730 <= reg_q730_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q730 <= reg_q730_init;
        else
          reg_q730 <= reg_q730_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1260_in <= (reg_q1258 AND symb_decoder(16#20#)) OR
 					(reg_q1258 AND symb_decoder(16#0a#)) OR
 					(reg_q1258 AND symb_decoder(16#0c#)) OR
 					(reg_q1258 AND symb_decoder(16#09#)) OR
 					(reg_q1258 AND symb_decoder(16#0d#)) OR
 					(reg_q1260 AND symb_decoder(16#0a#)) OR
 					(reg_q1260 AND symb_decoder(16#20#)) OR
 					(reg_q1260 AND symb_decoder(16#0c#)) OR
 					(reg_q1260 AND symb_decoder(16#09#)) OR
 					(reg_q1260 AND symb_decoder(16#0d#));
reg_q1260_init <= '0' ;
	p_reg_q1260: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1260 <= reg_q1260_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1260 <= reg_q1260_init;
        else
          reg_q1260 <= reg_q1260_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1387_in <= (reg_q1385 AND symb_decoder(16#61#)) OR
 					(reg_q1385 AND symb_decoder(16#41#));
reg_q1387_init <= '0' ;
	p_reg_q1387: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1387 <= reg_q1387_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1387 <= reg_q1387_init;
        else
          reg_q1387 <= reg_q1387_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1389_in <= (reg_q1387 AND symb_decoder(16#6d#)) OR
 					(reg_q1387 AND symb_decoder(16#4d#));
reg_q1389_init <= '0' ;
	p_reg_q1389: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1389 <= reg_q1389_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1389 <= reg_q1389_init;
        else
          reg_q1389 <= reg_q1389_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1979_in <= (reg_q1997 AND symb_decoder(16#23#)) OR
 					(reg_q1975 AND symb_decoder(16#23#));
reg_q1979_init <= '0' ;
	p_reg_q1979: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1979 <= reg_q1979_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1979 <= reg_q1979_init;
        else
          reg_q1979 <= reg_q1979_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q442_in <= (reg_q440 AND symb_decoder(16#76#)) OR
 					(reg_q440 AND symb_decoder(16#56#));
reg_q442_init <= '0' ;
	p_reg_q442: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q442 <= reg_q442_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q442 <= reg_q442_init;
        else
          reg_q442 <= reg_q442_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q444_in <= (reg_q442 AND symb_decoder(16#65#)) OR
 					(reg_q442 AND symb_decoder(16#45#));
reg_q444_init <= '0' ;
	p_reg_q444: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q444 <= reg_q444_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q444 <= reg_q444_init;
        else
          reg_q444 <= reg_q444_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1092_in <= (reg_q1090 AND symb_decoder(16#0c#)) OR
 					(reg_q1090 AND symb_decoder(16#0d#)) OR
 					(reg_q1090 AND symb_decoder(16#0a#)) OR
 					(reg_q1090 AND symb_decoder(16#20#)) OR
 					(reg_q1090 AND symb_decoder(16#09#)) OR
 					(reg_q1092 AND symb_decoder(16#20#)) OR
 					(reg_q1092 AND symb_decoder(16#09#)) OR
 					(reg_q1092 AND symb_decoder(16#0c#)) OR
 					(reg_q1092 AND symb_decoder(16#0d#)) OR
 					(reg_q1092 AND symb_decoder(16#0a#));
reg_q1092_init <= '0' ;
	p_reg_q1092: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1092 <= reg_q1092_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1092 <= reg_q1092_init;
        else
          reg_q1092 <= reg_q1092_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1594_in <= (reg_q1592 AND symb_decoder(16#49#)) OR
 					(reg_q1592 AND symb_decoder(16#69#));
reg_q1594_init <= '0' ;
	p_reg_q1594: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1594 <= reg_q1594_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1594 <= reg_q1594_init;
        else
          reg_q1594 <= reg_q1594_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1596_in <= (reg_q1594 AND symb_decoder(16#43#)) OR
 					(reg_q1594 AND symb_decoder(16#63#));
reg_q1596_init <= '0' ;
	p_reg_q1596: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1596 <= reg_q1596_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1596 <= reg_q1596_init;
        else
          reg_q1596 <= reg_q1596_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2260_in <= (reg_q2258 AND symb_decoder(16#4f#)) OR
 					(reg_q2258 AND symb_decoder(16#6f#));
reg_q2260_init <= '0' ;
	p_reg_q2260: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2260 <= reg_q2260_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2260 <= reg_q2260_init;
        else
          reg_q2260 <= reg_q2260_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1956_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1955 AND symb_decoder(16#0a#)) OR
 					(reg_q1955 AND symb_decoder(16#0d#));
reg_q1956_init <= '0' ;
	p_reg_q1956: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1956 <= reg_q1956_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1956 <= reg_q1956_init;
        else
          reg_q1956 <= reg_q1956_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1858_in <= (reg_q1856 AND symb_decoder(16#49#)) OR
 					(reg_q1856 AND symb_decoder(16#69#));
reg_q1858_init <= '0' ;
	p_reg_q1858: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1858 <= reg_q1858_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1858 <= reg_q1858_init;
        else
          reg_q1858 <= reg_q1858_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1860_in <= (reg_q1858 AND symb_decoder(16#44#)) OR
 					(reg_q1858 AND symb_decoder(16#64#));
reg_q1860_init <= '0' ;
	p_reg_q1860: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1860 <= reg_q1860_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1860 <= reg_q1860_init;
        else
          reg_q1860 <= reg_q1860_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1397_in <= (reg_q1395 AND symb_decoder(16#63#)) OR
 					(reg_q1395 AND symb_decoder(16#43#));
reg_q1397_init <= '0' ;
	p_reg_q1397: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1397 <= reg_q1397_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1397 <= reg_q1397_init;
        else
          reg_q1397 <= reg_q1397_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q78_in <= (reg_q76 AND symb_decoder(16#72#)) OR
 					(reg_q76 AND symb_decoder(16#52#));
reg_q78_init <= '0' ;
	p_reg_q78: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q78 <= reg_q78_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q78 <= reg_q78_init;
        else
          reg_q78 <= reg_q78_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q229_in <= (reg_q227 AND symb_decoder(16#36#));
reg_q229_init <= '0' ;
	p_reg_q229: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q229 <= reg_q229_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q229 <= reg_q229_init;
        else
          reg_q229 <= reg_q229_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q666_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q665 AND symb_decoder(16#0a#)) OR
 					(reg_q665 AND symb_decoder(16#0d#));
reg_q666_init <= '0' ;
	p_reg_q666: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q666 <= reg_q666_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q666 <= reg_q666_init;
        else
          reg_q666 <= reg_q666_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1619_in <= (reg_q1617 AND symb_decoder(16#45#)) OR
 					(reg_q1617 AND symb_decoder(16#65#));
reg_q1619_init <= '0' ;
	p_reg_q1619: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1619 <= reg_q1619_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1619 <= reg_q1619_init;
        else
          reg_q1619 <= reg_q1619_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q10_in <= (reg_q8 AND symb_decoder(16#69#)) OR
 					(reg_q8 AND symb_decoder(16#49#));
reg_q10_init <= '0' ;
	p_reg_q10: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q10 <= reg_q10_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q10 <= reg_q10_init;
        else
          reg_q10 <= reg_q10_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1872_in <= (reg_q1870 AND symb_decoder(16#6f#)) OR
 					(reg_q1870 AND symb_decoder(16#4f#));
reg_q1872_init <= '0' ;
	p_reg_q1872: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1872 <= reg_q1872_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1872 <= reg_q1872_init;
        else
          reg_q1872 <= reg_q1872_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1874_in <= (reg_q1872 AND symb_decoder(16#52#)) OR
 					(reg_q1872 AND symb_decoder(16#72#));
reg_q1874_init <= '0' ;
	p_reg_q1874: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1874 <= reg_q1874_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1874 <= reg_q1874_init;
        else
          reg_q1874 <= reg_q1874_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1299_in <= (reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1298 AND symb_decoder(16#67#)) OR
 					(reg_q1298 AND symb_decoder(16#47#));
reg_q1299_init <= '0' ;
	p_reg_q1299: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1299 <= reg_q1299_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1299 <= reg_q1299_init;
        else
          reg_q1299 <= reg_q1299_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q93_in <= (reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q92 AND symb_decoder(16#30#));
reg_q93_init <= '0' ;
	p_reg_q93: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q93 <= reg_q93_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q93 <= reg_q93_init;
        else
          reg_q93 <= reg_q93_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q95_in <= (reg_q93 AND symb_decoder(16#30#));
reg_q95_init <= '0' ;
	p_reg_q95: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q95 <= reg_q95_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q95 <= reg_q95_init;
        else
          reg_q95 <= reg_q95_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q391_in <= (reg_q389 AND symb_decoder(16#45#)) OR
 					(reg_q389 AND symb_decoder(16#65#));
reg_q391_init <= '0' ;
	p_reg_q391: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q391 <= reg_q391_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q391 <= reg_q391_init;
        else
          reg_q391 <= reg_q391_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q393_in <= (reg_q391 AND symb_decoder(16#4e#)) OR
 					(reg_q391 AND symb_decoder(16#6e#));
reg_q393_init <= '0' ;
	p_reg_q393: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q393 <= reg_q393_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q393 <= reg_q393_init;
        else
          reg_q393 <= reg_q393_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q28_in <= (reg_q26 AND symb_decoder(16#45#)) OR
 					(reg_q26 AND symb_decoder(16#65#));
reg_q28_init <= '0' ;
	p_reg_q28: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q28 <= reg_q28_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q28 <= reg_q28_init;
        else
          reg_q28 <= reg_q28_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1961_in <= (reg_q1959 AND symb_decoder(16#23#));
reg_q1961_init <= '0' ;
	p_reg_q1961: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1961 <= reg_q1961_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1961 <= reg_q1961_init;
        else
          reg_q1961 <= reg_q1961_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q389_in <= (reg_q387 AND symb_decoder(16#65#)) OR
 					(reg_q387 AND symb_decoder(16#45#));
reg_q389_init <= '0' ;
	p_reg_q389: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q389 <= reg_q389_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q389 <= reg_q389_init;
        else
          reg_q389 <= reg_q389_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q756_in <= (reg_q754 AND symb_decoder(16#0d#)) OR
 					(reg_q754 AND symb_decoder(16#0a#)) OR
 					(reg_q754 AND symb_decoder(16#20#)) OR
 					(reg_q754 AND symb_decoder(16#09#)) OR
 					(reg_q754 AND symb_decoder(16#0c#)) OR
 					(reg_q756 AND symb_decoder(16#20#)) OR
 					(reg_q756 AND symb_decoder(16#0c#)) OR
 					(reg_q756 AND symb_decoder(16#0a#)) OR
 					(reg_q756 AND symb_decoder(16#0d#)) OR
 					(reg_q756 AND symb_decoder(16#09#));
reg_q756_init <= '0' ;
	p_reg_q756: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q756 <= reg_q756_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q756 <= reg_q756_init;
        else
          reg_q756 <= reg_q756_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1760_in <= (reg_q1758 AND symb_decoder(16#20#)) OR
 					(reg_q1758 AND symb_decoder(16#0c#)) OR
 					(reg_q1758 AND symb_decoder(16#0d#)) OR
 					(reg_q1758 AND symb_decoder(16#0a#)) OR
 					(reg_q1758 AND symb_decoder(16#09#));
reg_q1760_init <= '0' ;
	p_reg_q1760: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1760 <= reg_q1760_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1760 <= reg_q1760_init;
        else
          reg_q1760 <= reg_q1760_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q838_in <= (reg_q836 AND symb_decoder(16#2e#));
reg_q838_init <= '0' ;
	p_reg_q838: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q838 <= reg_q838_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q838 <= reg_q838_init;
        else
          reg_q838 <= reg_q838_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q824_in <= (reg_q822 AND symb_decoder(16#6e#)) OR
 					(reg_q822 AND symb_decoder(16#4e#));
reg_q824_init <= '0' ;
	p_reg_q824: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q824 <= reg_q824_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q824 <= reg_q824_init;
        else
          reg_q824 <= reg_q824_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q826_in <= (reg_q824 AND symb_decoder(16#46#)) OR
 					(reg_q824 AND symb_decoder(16#66#));
reg_q826_init <= '0' ;
	p_reg_q826: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q826 <= reg_q826_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q826 <= reg_q826_init;
        else
          reg_q826 <= reg_q826_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2680_in <= (reg_q2678 AND symb_decoder(16#61#)) OR
 					(reg_q2678 AND symb_decoder(16#41#));
reg_q2680_init <= '0' ;
	p_reg_q2680: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2680 <= reg_q2680_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2680 <= reg_q2680_init;
        else
          reg_q2680 <= reg_q2680_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2682_in <= (reg_q2680 AND symb_decoder(16#52#)) OR
 					(reg_q2680 AND symb_decoder(16#72#));
reg_q2682_init <= '0' ;
	p_reg_q2682: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2682 <= reg_q2682_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2682 <= reg_q2682_init;
        else
          reg_q2682 <= reg_q2682_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q858_in <= (reg_q856 AND symb_decoder(16#69#)) OR
 					(reg_q856 AND symb_decoder(16#49#));
reg_q858_init <= '0' ;
	p_reg_q858: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q858 <= reg_q858_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q858 <= reg_q858_init;
        else
          reg_q858 <= reg_q858_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q860_in <= (reg_q858 AND symb_decoder(16#76#)) OR
 					(reg_q858 AND symb_decoder(16#56#));
reg_q860_init <= '0' ;
	p_reg_q860: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q860 <= reg_q860_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q860 <= reg_q860_init;
        else
          reg_q860 <= reg_q860_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q874_in <= (reg_q872 AND symb_decoder(16#5c#));
reg_q874_init <= '0' ;
	p_reg_q874: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q874 <= reg_q874_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q874 <= reg_q874_init;
        else
          reg_q874 <= reg_q874_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2656_in <= (reg_q2654 AND symb_decoder(16#45#)) OR
 					(reg_q2654 AND symb_decoder(16#65#));
reg_q2656_init <= '0' ;
	p_reg_q2656: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2656 <= reg_q2656_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2656 <= reg_q2656_init;
        else
          reg_q2656 <= reg_q2656_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q656_in <= (reg_q654 AND symb_decoder(16#31#));
reg_q656_init <= '0' ;
	p_reg_q656: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q656 <= reg_q656_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q656 <= reg_q656_init;
        else
          reg_q656 <= reg_q656_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q407_in <= (reg_q405 AND symb_decoder(16#45#)) OR
 					(reg_q405 AND symb_decoder(16#65#));
reg_q407_init <= '0' ;
	p_reg_q407: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q407 <= reg_q407_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q407 <= reg_q407_init;
        else
          reg_q407 <= reg_q407_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1466_in <= (reg_q1464 AND symb_decoder(16#72#)) OR
 					(reg_q1464 AND symb_decoder(16#52#));
reg_q1466_init <= '0' ;
	p_reg_q1466: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1466 <= reg_q1466_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1466 <= reg_q1466_init;
        else
          reg_q1466 <= reg_q1466_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2349_in <= (reg_q2347 AND symb_decoder(16#65#)) OR
 					(reg_q2347 AND symb_decoder(16#45#));
reg_q2349_init <= '0' ;
	p_reg_q2349: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2349 <= reg_q2349_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2349 <= reg_q2349_init;
        else
          reg_q2349 <= reg_q2349_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1525_in <= (reg_q1523 AND symb_decoder(16#45#)) OR
 					(reg_q1523 AND symb_decoder(16#65#));
reg_q1525_init <= '0' ;
	p_reg_q1525: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1525 <= reg_q1525_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1525 <= reg_q1525_init;
        else
          reg_q1525 <= reg_q1525_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1351_in <= (reg_q1349 AND symb_decoder(16#72#)) OR
 					(reg_q1349 AND symb_decoder(16#52#));
reg_q1351_init <= '0' ;
	p_reg_q1351: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1351 <= reg_q1351_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1351 <= reg_q1351_init;
        else
          reg_q1351 <= reg_q1351_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1353_in <= (reg_q1351 AND symb_decoder(16#54#)) OR
 					(reg_q1351 AND symb_decoder(16#74#));
reg_q1353_init <= '0' ;
	p_reg_q1353: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1353 <= reg_q1353_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1353 <= reg_q1353_init;
        else
          reg_q1353 <= reg_q1353_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1564_in <= (reg_q1562 AND symb_decoder(16#72#)) OR
 					(reg_q1562 AND symb_decoder(16#52#));
reg_q1564_init <= '0' ;
	p_reg_q1564: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1564 <= reg_q1564_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1564 <= reg_q1564_init;
        else
          reg_q1564 <= reg_q1564_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q115_in <= (reg_q113 AND symb_decoder(16#72#)) OR
 					(reg_q113 AND symb_decoder(16#52#));
reg_q115_init <= '0' ;
	p_reg_q115: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q115 <= reg_q115_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q115 <= reg_q115_init;
        else
          reg_q115 <= reg_q115_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q117_in <= (reg_q115 AND symb_decoder(16#4f#)) OR
 					(reg_q115 AND symb_decoder(16#6f#));
reg_q117_init <= '0' ;
	p_reg_q117: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q117 <= reg_q117_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q117 <= reg_q117_init;
        else
          reg_q117 <= reg_q117_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1123_in <= (reg_q1121 AND symb_decoder(16#64#)) OR
 					(reg_q1121 AND symb_decoder(16#44#));
reg_q1123_init <= '0' ;
	p_reg_q1123: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1123 <= reg_q1123_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1123 <= reg_q1123_init;
        else
          reg_q1123 <= reg_q1123_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q550_in <= (reg_q548 AND symb_decoder(16#72#)) OR
 					(reg_q548 AND symb_decoder(16#52#));
reg_q550_init <= '0' ;
	p_reg_q550: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q550 <= reg_q550_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q550 <= reg_q550_init;
        else
          reg_q550 <= reg_q550_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q552_in <= (reg_q550 AND symb_decoder(16#74#)) OR
 					(reg_q550 AND symb_decoder(16#54#));
reg_q552_init <= '0' ;
	p_reg_q552: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q552 <= reg_q552_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q552 <= reg_q552_init;
        else
          reg_q552 <= reg_q552_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2026_in <= (reg_q2024 AND symb_decoder(16#6e#)) OR
 					(reg_q2024 AND symb_decoder(16#4e#));
reg_q2026_init <= '0' ;
	p_reg_q2026: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2026 <= reg_q2026_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2026 <= reg_q2026_init;
        else
          reg_q2026 <= reg_q2026_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q317_in <= (reg_q315 AND symb_decoder(16#00#));
reg_q317_init <= '0' ;
	p_reg_q317: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q317 <= reg_q317_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q317 <= reg_q317_init;
        else
          reg_q317 <= reg_q317_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q319_in <= (reg_q317 AND symb_decoder(16#00#));
reg_q319_init <= '0' ;
	p_reg_q319: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q319 <= reg_q319_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q319 <= reg_q319_init;
        else
          reg_q319 <= reg_q319_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1225_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1224 AND symb_decoder(16#0d#)) OR
 					(reg_q1224 AND symb_decoder(16#0a#));
reg_q1225_init <= '0' ;
	p_reg_q1225: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1225 <= reg_q1225_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1225 <= reg_q1225_init;
        else
          reg_q1225 <= reg_q1225_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1782_in <= (reg_q1780 AND symb_decoder(16#20#)) OR
 					(reg_q1780 AND symb_decoder(16#0d#)) OR
 					(reg_q1780 AND symb_decoder(16#0c#)) OR
 					(reg_q1780 AND symb_decoder(16#0a#)) OR
 					(reg_q1780 AND symb_decoder(16#09#));
reg_q1782_init <= '0' ;
	p_reg_q1782: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1782 <= reg_q1782_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1782 <= reg_q1782_init;
        else
          reg_q1782 <= reg_q1782_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q409_in <= (reg_q407 AND symb_decoder(16#63#)) OR
 					(reg_q407 AND symb_decoder(16#43#));
reg_q409_init <= '0' ;
	p_reg_q409: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q409 <= reg_q409_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q409 <= reg_q409_init;
        else
          reg_q409 <= reg_q409_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q411_in <= (reg_q409 AND symb_decoder(16#54#)) OR
 					(reg_q409 AND symb_decoder(16#74#));
reg_q411_init <= '0' ;
	p_reg_q411: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q411 <= reg_q411_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q411 <= reg_q411_init;
        else
          reg_q411 <= reg_q411_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2188_in <= (reg_q2186 AND symb_decoder(16#4e#)) OR
 					(reg_q2186 AND symb_decoder(16#6e#));
reg_q2188_init <= '0' ;
	p_reg_q2188: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2188 <= reg_q2188_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2188 <= reg_q2188_init;
        else
          reg_q2188 <= reg_q2188_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2190_in <= (reg_q2188 AND symb_decoder(16#41#)) OR
 					(reg_q2188 AND symb_decoder(16#61#));
reg_q2190_init <= '0' ;
	p_reg_q2190: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2190 <= reg_q2190_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2190 <= reg_q2190_init;
        else
          reg_q2190 <= reg_q2190_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1177_in <= (reg_q1175 AND symb_decoder(16#6f#)) OR
 					(reg_q1175 AND symb_decoder(16#4f#));
reg_q1177_init <= '0' ;
	p_reg_q1177: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1177 <= reg_q1177_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1177 <= reg_q1177_init;
        else
          reg_q1177 <= reg_q1177_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2672_in <= (reg_q2670 AND symb_decoder(16#47#)) OR
 					(reg_q2670 AND symb_decoder(16#67#));
reg_q2672_init <= '0' ;
	p_reg_q2672: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2672 <= reg_q2672_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2672 <= reg_q2672_init;
        else
          reg_q2672 <= reg_q2672_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2674_in <= (reg_q2672 AND symb_decoder(16#0c#)) OR
 					(reg_q2672 AND symb_decoder(16#0d#)) OR
 					(reg_q2672 AND symb_decoder(16#20#)) OR
 					(reg_q2672 AND symb_decoder(16#0a#)) OR
 					(reg_q2672 AND symb_decoder(16#09#));
reg_q2674_init <= '0' ;
	p_reg_q2674: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2674 <= reg_q2674_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2674 <= reg_q2674_init;
        else
          reg_q2674 <= reg_q2674_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q634_in <= (reg_q632 AND symb_decoder(16#4f#)) OR
 					(reg_q632 AND symb_decoder(16#6f#));
reg_q634_init <= '0' ;
	p_reg_q634: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q634 <= reg_q634_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q634 <= reg_q634_init;
        else
          reg_q634 <= reg_q634_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2125_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2124 AND symb_decoder(16#0d#)) OR
 					(reg_q2124 AND symb_decoder(16#0a#));
reg_q2125_init <= '0' ;
	p_reg_q2125: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2125 <= reg_q2125_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2125 <= reg_q2125_init;
        else
          reg_q2125 <= reg_q2125_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2126_in <= (reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2125 AND symb_decoder(16#57#)) OR
 					(reg_q2125 AND symb_decoder(16#77#));
reg_q2126_init <= '0' ;
	p_reg_q2126: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2126 <= reg_q2126_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2126 <= reg_q2126_init;
        else
          reg_q2126 <= reg_q2126_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1878_in <= (reg_q1876 AND symb_decoder(16#61#)) OR
 					(reg_q1876 AND symb_decoder(16#41#));
reg_q1878_init <= '0' ;
	p_reg_q1878: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1878 <= reg_q1878_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1878 <= reg_q1878_init;
        else
          reg_q1878 <= reg_q1878_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q681_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q680 AND symb_decoder(16#0a#)) OR
 					(reg_q680 AND symb_decoder(16#0d#));
reg_q681_init <= '0' ;
	p_reg_q681: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q681 <= reg_q681_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q681 <= reg_q681_init;
        else
          reg_q681 <= reg_q681_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1836_in <= (reg_q1834 AND symb_decoder(16#49#)) OR
 					(reg_q1834 AND symb_decoder(16#69#));
reg_q1836_init <= '0' ;
	p_reg_q1836: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1836 <= reg_q1836_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1836 <= reg_q1836_init;
        else
          reg_q1836 <= reg_q1836_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1838_in <= (reg_q1836 AND symb_decoder(16#4e#)) OR
 					(reg_q1836 AND symb_decoder(16#6e#));
reg_q1838_init <= '0' ;
	p_reg_q1838: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1838 <= reg_q1838_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1838 <= reg_q1838_init;
        else
          reg_q1838 <= reg_q1838_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1458_in <= (reg_q1456 AND symb_decoder(16#41#)) OR
 					(reg_q1456 AND symb_decoder(16#61#));
reg_q1458_init <= '0' ;
	p_reg_q1458: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1458 <= reg_q1458_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1458 <= reg_q1458_init;
        else
          reg_q1458 <= reg_q1458_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q787_in <= (reg_q785 AND symb_decoder(16#6e#)) OR
 					(reg_q785 AND symb_decoder(16#4e#));
reg_q787_init <= '0' ;
	p_reg_q787: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q787 <= reg_q787_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q787 <= reg_q787_init;
        else
          reg_q787 <= reg_q787_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1391_in <= (reg_q1389 AND symb_decoder(16#45#)) OR
 					(reg_q1389 AND symb_decoder(16#65#));
reg_q1391_init <= '0' ;
	p_reg_q1391: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1391 <= reg_q1391_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1391 <= reg_q1391_init;
        else
          reg_q1391 <= reg_q1391_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1888_in <= (reg_q1886 AND symb_decoder(16#68#)) OR
 					(reg_q1886 AND symb_decoder(16#48#));
reg_q1888_init <= '0' ;
	p_reg_q1888: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1888 <= reg_q1888_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1888 <= reg_q1888_init;
        else
          reg_q1888 <= reg_q1888_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1876_in <= (reg_q1874 AND symb_decoder(16#74#)) OR
 					(reg_q1874 AND symb_decoder(16#54#));
reg_q1876_init <= '0' ;
	p_reg_q1876: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1876 <= reg_q1876_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1876 <= reg_q1876_init;
        else
          reg_q1876 <= reg_q1876_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1898_in <= (reg_q1896 AND symb_decoder(16#6e#)) OR
 					(reg_q1896 AND symb_decoder(16#4e#));
reg_q1898_init <= '0' ;
	p_reg_q1898: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1898 <= reg_q1898_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1898 <= reg_q1898_init;
        else
          reg_q1898 <= reg_q1898_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2176_in <= (reg_q2172 AND symb_decoder(16#66#)) OR
 					(reg_q2172 AND symb_decoder(16#46#)) OR
 					(reg_q2208 AND symb_decoder(16#66#)) OR
 					(reg_q2208 AND symb_decoder(16#46#));
reg_q2176_init <= '0' ;
	p_reg_q2176: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2176 <= reg_q2176_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2176 <= reg_q2176_init;
        else
          reg_q2176 <= reg_q2176_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q434_in <= (reg_q432 AND symb_decoder(16#4e#)) OR
 					(reg_q432 AND symb_decoder(16#6e#));
reg_q434_init <= '0' ;
	p_reg_q434: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q434 <= reg_q434_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q434 <= reg_q434_init;
        else
          reg_q434 <= reg_q434_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q436_in <= (reg_q434 AND symb_decoder(16#65#)) OR
 					(reg_q434 AND symb_decoder(16#45#));
reg_q436_init <= '0' ;
	p_reg_q436: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q436 <= reg_q436_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q436 <= reg_q436_init;
        else
          reg_q436 <= reg_q436_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1494_in <= (reg_q1492 AND symb_decoder(16#45#)) OR
 					(reg_q1492 AND symb_decoder(16#65#));
reg_q1494_init <= '0' ;
	p_reg_q1494: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1494 <= reg_q1494_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1494 <= reg_q1494_init;
        else
          reg_q1494 <= reg_q1494_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2146_in <= (reg_q2144 AND symb_decoder(16#73#)) OR
 					(reg_q2144 AND symb_decoder(16#53#));
reg_q2146_init <= '0' ;
	p_reg_q2146: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2146 <= reg_q2146_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2146 <= reg_q2146_init;
        else
          reg_q2146 <= reg_q2146_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1788_in <= (reg_q1786 AND symb_decoder(16#20#)) OR
 					(reg_q1786 AND symb_decoder(16#0a#)) OR
 					(reg_q1786 AND symb_decoder(16#09#)) OR
 					(reg_q1786 AND symb_decoder(16#0c#)) OR
 					(reg_q1786 AND symb_decoder(16#0d#));
reg_q1788_init <= '0' ;
	p_reg_q1788: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1788 <= reg_q1788_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1788 <= reg_q1788_init;
        else
          reg_q1788 <= reg_q1788_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q270_in <= (reg_q268 AND symb_decoder(16#31#));
reg_q270_init <= '0' ;
	p_reg_q270: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q270 <= reg_q270_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q270 <= reg_q270_init;
        else
          reg_q270 <= reg_q270_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1347_in <= (reg_q1345 AND symb_decoder(16#70#)) OR
 					(reg_q1345 AND symb_decoder(16#50#));
reg_q1347_init <= '0' ;
	p_reg_q1347: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1347 <= reg_q1347_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1347 <= reg_q1347_init;
        else
          reg_q1347 <= reg_q1347_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1349_in <= (reg_q1347 AND symb_decoder(16#4f#)) OR
 					(reg_q1347 AND symb_decoder(16#6f#));
reg_q1349_init <= '0' ;
	p_reg_q1349: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1349 <= reg_q1349_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1349 <= reg_q1349_init;
        else
          reg_q1349 <= reg_q1349_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1238_in <= (reg_q1236 AND symb_decoder(16#41#)) OR
 					(reg_q1236 AND symb_decoder(16#61#));
reg_q1238_init <= '0' ;
	p_reg_q1238: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1238 <= reg_q1238_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1238 <= reg_q1238_init;
        else
          reg_q1238 <= reg_q1238_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1240_in <= (reg_q1238 AND symb_decoder(16#53#)) OR
 					(reg_q1238 AND symb_decoder(16#73#));
reg_q1240_init <= '0' ;
	p_reg_q1240: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1240 <= reg_q1240_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1240 <= reg_q1240_init;
        else
          reg_q1240 <= reg_q1240_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q422_in <= (reg_q420 AND symb_decoder(16#64#)) OR
 					(reg_q420 AND symb_decoder(16#44#));
reg_q422_init <= '0' ;
	p_reg_q422: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q422 <= reg_q422_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q422 <= reg_q422_init;
        else
          reg_q422 <= reg_q422_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q982_in <= (reg_q980 AND symb_decoder(16#54#)) OR
 					(reg_q980 AND symb_decoder(16#74#));
reg_q982_init <= '0' ;
	p_reg_q982: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q982 <= reg_q982_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q982 <= reg_q982_init;
        else
          reg_q982 <= reg_q982_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1562_in <= (reg_q1560 AND symb_decoder(16#65#)) OR
 					(reg_q1560 AND symb_decoder(16#45#));
reg_q1562_init <= '0' ;
	p_reg_q1562: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1562 <= reg_q1562_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1562 <= reg_q1562_init;
        else
          reg_q1562 <= reg_q1562_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q817_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q816 AND symb_decoder(16#0a#)) OR
 					(reg_q816 AND symb_decoder(16#0d#));
reg_q817_init <= '0' ;
	p_reg_q817: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q817 <= reg_q817_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q817 <= reg_q817_init;
        else
          reg_q817 <= reg_q817_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q818_in <= (reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q817 AND symb_decoder(16#64#)) OR
 					(reg_q817 AND symb_decoder(16#44#));
reg_q818_init <= '0' ;
	p_reg_q818: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q818 <= reg_q818_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q818 <= reg_q818_init;
        else
          reg_q818 <= reg_q818_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q263_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q262 AND symb_decoder(16#0d#)) OR
 					(reg_q262 AND symb_decoder(16#0a#));
reg_q263_init <= '0' ;
	p_reg_q263: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q263 <= reg_q263_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q263 <= reg_q263_init;
        else
          reg_q263 <= reg_q263_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q264_in <= (reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q263 AND symb_decoder(16#41#)) OR
 					(reg_q263 AND symb_decoder(16#61#));
reg_q264_init <= '0' ;
	p_reg_q264: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q264 <= reg_q264_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q264 <= reg_q264_init;
        else
          reg_q264 <= reg_q264_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q470_in <= (reg_q468 AND symb_decoder(16#72#)) OR
 					(reg_q468 AND symb_decoder(16#52#));
reg_q470_init <= '0' ;
	p_reg_q470: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q470 <= reg_q470_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q470 <= reg_q470_init;
        else
          reg_q470 <= reg_q470_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1096_in <= (reg_q1096 AND symb_decoder(16#09#)) OR
 					(reg_q1096 AND symb_decoder(16#0a#)) OR
 					(reg_q1096 AND symb_decoder(16#0d#)) OR
 					(reg_q1096 AND symb_decoder(16#20#)) OR
 					(reg_q1096 AND symb_decoder(16#0c#)) OR
 					(reg_q1094 AND symb_decoder(16#09#)) OR
 					(reg_q1094 AND symb_decoder(16#0c#)) OR
 					(reg_q1094 AND symb_decoder(16#0d#)) OR
 					(reg_q1094 AND symb_decoder(16#20#)) OR
 					(reg_q1094 AND symb_decoder(16#0a#));
reg_q1096_init <= '0' ;
	p_reg_q1096: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1096 <= reg_q1096_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1096 <= reg_q1096_init;
        else
          reg_q1096 <= reg_q1096_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2441_in <= (reg_q2439 AND symb_decoder(16#41#)) OR
 					(reg_q2439 AND symb_decoder(16#61#));
reg_q2441_init <= '0' ;
	p_reg_q2441: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2441 <= reg_q2441_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2441 <= reg_q2441_init;
        else
          reg_q2441 <= reg_q2441_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2443_in <= (reg_q2441 AND symb_decoder(16#64#)) OR
 					(reg_q2441 AND symb_decoder(16#44#));
reg_q2443_init <= '0' ;
	p_reg_q2443: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2443 <= reg_q2443_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2443 <= reg_q2443_init;
        else
          reg_q2443 <= reg_q2443_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1590_in <= (reg_q1588 AND symb_decoder(16#72#)) OR
 					(reg_q1588 AND symb_decoder(16#52#));
reg_q1590_init <= '0' ;
	p_reg_q1590: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1590 <= reg_q1590_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1590 <= reg_q1590_init;
        else
          reg_q1590 <= reg_q1590_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1592_in <= (reg_q1590 AND symb_decoder(16#76#)) OR
 					(reg_q1590 AND symb_decoder(16#56#));
reg_q1592_init <= '0' ;
	p_reg_q1592: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1592 <= reg_q1592_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1592 <= reg_q1592_init;
        else
          reg_q1592 <= reg_q1592_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1774_in <= (reg_q1772 AND symb_decoder(16#0d#)) OR
 					(reg_q1772 AND symb_decoder(16#0c#)) OR
 					(reg_q1772 AND symb_decoder(16#0a#)) OR
 					(reg_q1772 AND symb_decoder(16#09#)) OR
 					(reg_q1772 AND symb_decoder(16#20#));
reg_q1774_init <= '0' ;
	p_reg_q1774: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1774 <= reg_q1774_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1774 <= reg_q1774_init;
        else
          reg_q1774 <= reg_q1774_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1776_in <= (reg_q1774 AND symb_decoder(16#0d#)) OR
 					(reg_q1774 AND symb_decoder(16#0a#)) OR
 					(reg_q1774 AND symb_decoder(16#0c#)) OR
 					(reg_q1774 AND symb_decoder(16#20#)) OR
 					(reg_q1774 AND symb_decoder(16#09#));
reg_q1776_init <= '0' ;
	p_reg_q1776: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1776 <= reg_q1776_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1776 <= reg_q1776_init;
        else
          reg_q1776 <= reg_q1776_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1094_in <= (reg_q1092 AND symb_decoder(16#2e#));
reg_q1094_init <= '0' ;
	p_reg_q1094: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1094 <= reg_q1094_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1094 <= reg_q1094_init;
        else
          reg_q1094 <= reg_q1094_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q927_in <= (reg_q925 AND symb_decoder(16#76#)) OR
 					(reg_q925 AND symb_decoder(16#56#));
reg_q927_init <= '0' ;
	p_reg_q927: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q927 <= reg_q927_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q927 <= reg_q927_init;
        else
          reg_q927 <= reg_q927_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q785_in <= (reg_q783 AND symb_decoder(16#49#)) OR
 					(reg_q783 AND symb_decoder(16#69#));
reg_q785_init <= '0' ;
	p_reg_q785: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q785 <= reg_q785_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q785 <= reg_q785_init;
        else
          reg_q785 <= reg_q785_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2611_in <= (reg_q2609 AND symb_decoder(16#3a#));
reg_q2611_init <= '0' ;
	p_reg_q2611: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2611 <= reg_q2611_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2611 <= reg_q2611_init;
        else
          reg_q2611 <= reg_q2611_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2423_in <= (reg_q2421 AND symb_decoder(16#74#)) OR
 					(reg_q2421 AND symb_decoder(16#54#));
reg_q2423_init <= '0' ;
	p_reg_q2423: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2423 <= reg_q2423_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2423 <= reg_q2423_init;
        else
          reg_q2423 <= reg_q2423_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1230_in <= (reg_q1228 AND symb_decoder(16#54#)) OR
 					(reg_q1228 AND symb_decoder(16#74#));
reg_q1230_init <= '0' ;
	p_reg_q1230: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1230 <= reg_q1230_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1230 <= reg_q1230_init;
        else
          reg_q1230 <= reg_q1230_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q994_in <= (reg_q992 AND symb_decoder(16#6c#)) OR
 					(reg_q992 AND symb_decoder(16#4c#));
reg_q994_init <= '0' ;
	p_reg_q994: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q994 <= reg_q994_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q994 <= reg_q994_init;
        else
          reg_q994 <= reg_q994_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q996_in <= (reg_q994 AND symb_decoder(16#46#)) OR
 					(reg_q994 AND symb_decoder(16#66#));
reg_q996_init <= '0' ;
	p_reg_q996: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q996 <= reg_q996_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q996 <= reg_q996_init;
        else
          reg_q996 <= reg_q996_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2144_in <= (reg_q2142 AND symb_decoder(16#69#)) OR
 					(reg_q2142 AND symb_decoder(16#49#));
reg_q2144_init <= '0' ;
	p_reg_q2144: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2144 <= reg_q2144_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2144 <= reg_q2144_init;
        else
          reg_q2144 <= reg_q2144_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1234_in <= (reg_q1232 AND symb_decoder(16#63#)) OR
 					(reg_q1232 AND symb_decoder(16#43#));
reg_q1234_init <= '0' ;
	p_reg_q1234: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1234 <= reg_q1234_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1234 <= reg_q1234_init;
        else
          reg_q1234 <= reg_q1234_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1236_in <= (reg_q1234 AND symb_decoder(16#52#)) OR
 					(reg_q1234 AND symb_decoder(16#72#));
reg_q1236_init <= '0' ;
	p_reg_q1236: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1236 <= reg_q1236_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1236 <= reg_q1236_init;
        else
          reg_q1236 <= reg_q1236_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2239_in <= (reg_q2237 AND symb_decoder(16#45#)) OR
 					(reg_q2237 AND symb_decoder(16#65#));
reg_q2239_init <= '0' ;
	p_reg_q2239: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2239 <= reg_q2239_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2239 <= reg_q2239_init;
        else
          reg_q2239 <= reg_q2239_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q992_in <= (reg_q990 AND symb_decoder(16#49#)) OR
 					(reg_q990 AND symb_decoder(16#69#));
reg_q992_init <= '0' ;
	p_reg_q992: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q992 <= reg_q992_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q992 <= reg_q992_init;
        else
          reg_q992 <= reg_q992_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q186_in <= (reg_q184 AND symb_decoder(16#30#));
reg_q186_init <= '0' ;
	p_reg_q186: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q186 <= reg_q186_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q186 <= reg_q186_init;
        else
          reg_q186 <= reg_q186_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q188_in <= (reg_q186 AND symb_decoder(16#31#));
reg_q188_init <= '0' ;
	p_reg_q188: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q188 <= reg_q188_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q188 <= reg_q188_init;
        else
          reg_q188 <= reg_q188_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1862_in <= (reg_q1860 AND symb_decoder(16#6f#)) OR
 					(reg_q1860 AND symb_decoder(16#4f#));
reg_q1862_init <= '0' ;
	p_reg_q1862: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1862 <= reg_q1862_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1862 <= reg_q1862_init;
        else
          reg_q1862 <= reg_q1862_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q153_in <= (reg_q151 AND symb_decoder(16#55#)) OR
 					(reg_q151 AND symb_decoder(16#75#));
reg_q153_init <= '0' ;
	p_reg_q153: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q153 <= reg_q153_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q153 <= reg_q153_init;
        else
          reg_q153 <= reg_q153_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1738_in <= (reg_q1736 AND symb_decoder(16#49#)) OR
 					(reg_q1736 AND symb_decoder(16#69#));
reg_q1738_init <= '0' ;
	p_reg_q1738: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1738 <= reg_q1738_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1738 <= reg_q1738_init;
        else
          reg_q1738 <= reg_q1738_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1740_in <= (reg_q1738 AND symb_decoder(16#53#)) OR
 					(reg_q1738 AND symb_decoder(16#73#));
reg_q1740_init <= '0' ;
	p_reg_q1740: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1740 <= reg_q1740_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1740 <= reg_q1740_init;
        else
          reg_q1740 <= reg_q1740_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q282_in <= (reg_q280 AND symb_decoder(16#74#)) OR
 					(reg_q280 AND symb_decoder(16#54#));
reg_q282_init <= '0' ;
	p_reg_q282: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q282 <= reg_q282_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q282 <= reg_q282_init;
        else
          reg_q282 <= reg_q282_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q284_in <= (reg_q282 AND symb_decoder(16#48#)) OR
 					(reg_q282 AND symb_decoder(16#68#));
reg_q284_init <= '0' ;
	p_reg_q284: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q284 <= reg_q284_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q284 <= reg_q284_init;
        else
          reg_q284 <= reg_q284_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2688_in <= (reg_q2686 AND symb_decoder(16#44#)) OR
 					(reg_q2686 AND symb_decoder(16#64#));
reg_q2688_init <= '0' ;
	p_reg_q2688: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2688 <= reg_q2688_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2688 <= reg_q2688_init;
        else
          reg_q2688 <= reg_q2688_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1280_in <= (reg_q1278 AND symb_decoder(16#2d#));
reg_q1280_init <= '0' ;
	p_reg_q1280: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1280 <= reg_q1280_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1280 <= reg_q1280_init;
        else
          reg_q1280 <= reg_q1280_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1282_in <= (reg_q1280 AND symb_decoder(16#4c#)) OR
 					(reg_q1280 AND symb_decoder(16#6c#));
reg_q1282_init <= '0' ;
	p_reg_q1282: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1282 <= reg_q1282_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1282 <= reg_q1282_init;
        else
          reg_q1282 <= reg_q1282_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q494_in <= (reg_q492 AND symb_decoder(16#6f#)) OR
 					(reg_q492 AND symb_decoder(16#4f#));
reg_q494_init <= '0' ;
	p_reg_q494: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q494 <= reg_q494_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q494 <= reg_q494_init;
        else
          reg_q494 <= reg_q494_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1694_in <= (reg_q1692 AND symb_decoder(16#67#)) OR
 					(reg_q1692 AND symb_decoder(16#47#));
reg_q1694_init <= '0' ;
	p_reg_q1694: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1694 <= reg_q1694_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1694 <= reg_q1694_init;
        else
          reg_q1694 <= reg_q1694_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1431_in <= (reg_q1429 AND symb_decoder(16#69#)) OR
 					(reg_q1429 AND symb_decoder(16#49#));
reg_q1431_init <= '0' ;
	p_reg_q1431: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1431 <= reg_q1431_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1431 <= reg_q1431_init;
        else
          reg_q1431 <= reg_q1431_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2325_in <= (reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2324 AND symb_decoder(16#22#));
reg_q2325_init <= '0' ;
	p_reg_q2325: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2325 <= reg_q2325_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2325 <= reg_q2325_init;
        else
          reg_q2325 <= reg_q2325_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2421_in <= (reg_q2419 AND symb_decoder(16#53#)) OR
 					(reg_q2419 AND symb_decoder(16#73#));
reg_q2421_init <= '0' ;
	p_reg_q2421: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2421 <= reg_q2421_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2421 <= reg_q2421_init;
        else
          reg_q2421 <= reg_q2421_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q290_in <= (reg_q288 AND symb_decoder(16#65#)) OR
 					(reg_q288 AND symb_decoder(16#45#));
reg_q290_init <= '0' ;
	p_reg_q290: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q290 <= reg_q290_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q290 <= reg_q290_init;
        else
          reg_q290 <= reg_q290_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1570_in <= (reg_q1568 AND symb_decoder(16#4f#)) OR
 					(reg_q1568 AND symb_decoder(16#6f#));
reg_q1570_init <= '0' ;
	p_reg_q1570: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1570 <= reg_q1570_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1570 <= reg_q1570_init;
        else
          reg_q1570 <= reg_q1570_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1662_in <= (reg_q1660 AND symb_decoder(16#76#)) OR
 					(reg_q1660 AND symb_decoder(16#56#));
reg_q1662_init <= '0' ;
	p_reg_q1662: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1662 <= reg_q1662_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1662 <= reg_q1662_init;
        else
          reg_q1662 <= reg_q1662_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2219_in <= (reg_q2217 AND symb_decoder(16#43#)) OR
 					(reg_q2217 AND symb_decoder(16#63#));
reg_q2219_init <= '0' ;
	p_reg_q2219: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2219 <= reg_q2219_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2219 <= reg_q2219_init;
        else
          reg_q2219 <= reg_q2219_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2605_in <= (reg_q2603 AND symb_decoder(16#73#)) OR
 					(reg_q2603 AND symb_decoder(16#53#));
reg_q2605_init <= '0' ;
	p_reg_q2605: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2605 <= reg_q2605_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2605 <= reg_q2605_init;
        else
          reg_q2605 <= reg_q2605_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2607_in <= (reg_q2605 AND symb_decoder(16#65#)) OR
 					(reg_q2605 AND symb_decoder(16#45#));
reg_q2607_init <= '0' ;
	p_reg_q2607: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2607 <= reg_q2607_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2607 <= reg_q2607_init;
        else
          reg_q2607 <= reg_q2607_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q32_in <= (reg_q30 AND symb_decoder(16#75#)) OR
 					(reg_q30 AND symb_decoder(16#55#));
reg_q32_init <= '0' ;
	p_reg_q32: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q32 <= reg_q32_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q32 <= reg_q32_init;
        else
          reg_q32 <= reg_q32_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q34_in <= (reg_q32 AND symb_decoder(16#74#)) OR
 					(reg_q32 AND symb_decoder(16#54#));
reg_q34_init <= '0' ;
	p_reg_q34: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q34 <= reg_q34_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q34 <= reg_q34_init;
        else
          reg_q34 <= reg_q34_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q339_in <= (reg_q337 AND symb_decoder(16#4e#)) OR
 					(reg_q337 AND symb_decoder(16#6e#));
reg_q339_init <= '0' ;
	p_reg_q339: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q339 <= reg_q339_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q339 <= reg_q339_init;
        else
          reg_q339 <= reg_q339_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q165_in <= (reg_q163 AND symb_decoder(16#66#)) OR
 					(reg_q163 AND symb_decoder(16#46#));
reg_q165_init <= '0' ;
	p_reg_q165: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q165 <= reg_q165_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q165 <= reg_q165_init;
        else
          reg_q165 <= reg_q165_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1508_in <= (reg_q1506 AND symb_decoder(16#45#)) OR
 					(reg_q1506 AND symb_decoder(16#65#));
reg_q1508_init <= '0' ;
	p_reg_q1508: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1508 <= reg_q1508_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1508 <= reg_q1508_init;
        else
          reg_q1508 <= reg_q1508_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q167_in <= (reg_q165 AND symb_decoder(16#55#)) OR
 					(reg_q165 AND symb_decoder(16#75#));
reg_q167_init <= '0' ;
	p_reg_q167: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q167 <= reg_q167_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q167 <= reg_q167_init;
        else
          reg_q167 <= reg_q167_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q169_in <= (reg_q167 AND symb_decoder(16#4c#)) OR
 					(reg_q167 AND symb_decoder(16#6c#));
reg_q169_init <= '0' ;
	p_reg_q169: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q169 <= reg_q169_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q169 <= reg_q169_init;
        else
          reg_q169 <= reg_q169_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q536_in <= (reg_q534 AND symb_decoder(16#5d#));
reg_q536_init <= '0' ;
	p_reg_q536: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q536 <= reg_q536_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q536 <= reg_q536_init;
        else
          reg_q536 <= reg_q536_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1232_in <= (reg_q1230 AND symb_decoder(16#45#)) OR
 					(reg_q1230 AND symb_decoder(16#65#));
reg_q1232_init <= '0' ;
	p_reg_q1232: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1232 <= reg_q1232_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1232 <= reg_q1232_init;
        else
          reg_q1232 <= reg_q1232_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q184_in <= (reg_q182 AND symb_decoder(16#30#));
reg_q184_init <= '0' ;
	p_reg_q184: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q184 <= reg_q184_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q184 <= reg_q184_init;
        else
          reg_q184 <= reg_q184_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q856_in <= (reg_q854 AND symb_decoder(16#72#)) OR
 					(reg_q854 AND symb_decoder(16#52#));
reg_q856_init <= '0' ;
	p_reg_q856: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q856 <= reg_q856_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q856 <= reg_q856_init;
        else
          reg_q856 <= reg_q856_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q718_in <= (reg_q716 AND symb_decoder(16#69#)) OR
 					(reg_q716 AND symb_decoder(16#49#));
reg_q718_init <= '0' ;
	p_reg_q718: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q718 <= reg_q718_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q718 <= reg_q718_init;
        else
          reg_q718 <= reg_q718_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1605_in <= (reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q1604 AND symb_decoder(16#4e#)) OR
 					(reg_q1604 AND symb_decoder(16#6e#));
reg_q1605_init <= '0' ;
	p_reg_q1605: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1605 <= reg_q1605_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1605 <= reg_q1605_init;
        else
          reg_q1605 <= reg_q1605_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2678_in <= (reg_q2676 AND symb_decoder(16#74#)) OR
 					(reg_q2676 AND symb_decoder(16#54#));
reg_q2678_init <= '0' ;
	p_reg_q2678: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2678 <= reg_q2678_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2678 <= reg_q2678_init;
        else
          reg_q2678 <= reg_q2678_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q917_in <= (reg_q915 AND symb_decoder(16#61#)) OR
 					(reg_q915 AND symb_decoder(16#41#));
reg_q917_init <= '0' ;
	p_reg_q917: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q917 <= reg_q917_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q917 <= reg_q917_init;
        else
          reg_q917 <= reg_q917_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q919_in <= (reg_q917 AND symb_decoder(16#20#)) OR
 					(reg_q917 AND symb_decoder(16#0d#)) OR
 					(reg_q917 AND symb_decoder(16#0a#)) OR
 					(reg_q917 AND symb_decoder(16#09#)) OR
 					(reg_q917 AND symb_decoder(16#0c#)) OR
 					(reg_q919 AND symb_decoder(16#0a#)) OR
 					(reg_q919 AND symb_decoder(16#09#)) OR
 					(reg_q919 AND symb_decoder(16#0d#)) OR
 					(reg_q919 AND symb_decoder(16#20#)) OR
 					(reg_q919 AND symb_decoder(16#0c#));
reg_q919_init <= '0' ;
	p_reg_q919: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q919 <= reg_q919_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q919 <= reg_q919_init;
        else
          reg_q919 <= reg_q919_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2001_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2000 AND symb_decoder(16#0d#)) OR
 					(reg_q2000 AND symb_decoder(16#0a#));
reg_q2001_init <= '0' ;
	p_reg_q2001: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2001 <= reg_q2001_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2001 <= reg_q2001_init;
        else
          reg_q2001 <= reg_q2001_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2036_in <= (reg_q2034 AND symb_decoder(16#4c#)) OR
 					(reg_q2034 AND symb_decoder(16#6c#));
reg_q2036_init <= '0' ;
	p_reg_q2036: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2036 <= reg_q2036_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2036 <= reg_q2036_init;
        else
          reg_q2036 <= reg_q2036_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q546_in <= (reg_q544 AND symb_decoder(16#70#)) OR
 					(reg_q544 AND symb_decoder(16#50#));
reg_q546_init <= '0' ;
	p_reg_q546: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q546 <= reg_q546_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q546 <= reg_q546_init;
        else
          reg_q546 <= reg_q546_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q548_in <= (reg_q546 AND symb_decoder(16#6f#)) OR
 					(reg_q546 AND symb_decoder(16#4f#));
reg_q548_init <= '0' ;
	p_reg_q548: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q548 <= reg_q548_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q548 <= reg_q548_init;
        else
          reg_q548 <= reg_q548_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2634_in <= (reg_q2632 AND symb_decoder(16#c0#));
reg_q2634_init <= '0' ;
	p_reg_q2634: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2634 <= reg_q2634_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2634 <= reg_q2634_init;
        else
          reg_q2634 <= reg_q2634_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2162_in <= (reg_q2160 AND symb_decoder(16#44#)) OR
 					(reg_q2160 AND symb_decoder(16#64#));
reg_q2162_init <= '0' ;
	p_reg_q2162: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2162 <= reg_q2162_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2162 <= reg_q2162_init;
        else
          reg_q2162 <= reg_q2162_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2365_in <= (reg_q2363 AND symb_decoder(16#52#)) OR
 					(reg_q2363 AND symb_decoder(16#72#));
reg_q2365_init <= '0' ;
	p_reg_q2365: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2365 <= reg_q2365_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2365 <= reg_q2365_init;
        else
          reg_q2365 <= reg_q2365_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q762_in <= (reg_q760 AND symb_decoder(16#52#)) OR
 					(reg_q760 AND symb_decoder(16#72#));
reg_q762_init <= '0' ;
	p_reg_q762: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q762 <= reg_q762_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q762 <= reg_q762_init;
        else
          reg_q762 <= reg_q762_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q764_in <= (reg_q762 AND symb_decoder(16#45#)) OR
 					(reg_q762 AND symb_decoder(16#65#));
reg_q764_init <= '0' ;
	p_reg_q764: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q764 <= reg_q764_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q764 <= reg_q764_init;
        else
          reg_q764 <= reg_q764_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q218_in <= (reg_q216 AND symb_decoder(16#6c#)) OR
 					(reg_q216 AND symb_decoder(16#4c#));
reg_q218_init <= '0' ;
	p_reg_q218: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q218 <= reg_q218_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q218 <= reg_q218_init;
        else
          reg_q218 <= reg_q218_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q220_in <= (reg_q218 AND symb_decoder(16#69#)) OR
 					(reg_q218 AND symb_decoder(16#49#));
reg_q220_init <= '0' ;
	p_reg_q220: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q220 <= reg_q220_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q220 <= reg_q220_init;
        else
          reg_q220 <= reg_q220_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1357_in <= (reg_q1355 AND symb_decoder(16#32#)) OR
 					(reg_q1355 AND symb_decoder(16#39#)) OR
 					(reg_q1355 AND symb_decoder(16#36#)) OR
 					(reg_q1355 AND symb_decoder(16#33#)) OR
 					(reg_q1355 AND symb_decoder(16#30#)) OR
 					(reg_q1355 AND symb_decoder(16#37#)) OR
 					(reg_q1355 AND symb_decoder(16#31#)) OR
 					(reg_q1355 AND symb_decoder(16#38#)) OR
 					(reg_q1355 AND symb_decoder(16#34#)) OR
 					(reg_q1355 AND symb_decoder(16#35#));
reg_q1357_init <= '0' ;
	p_reg_q1357: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1357 <= reg_q1357_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1357 <= reg_q1357_init;
        else
          reg_q1357 <= reg_q1357_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1995_in <= (reg_q1993 AND symb_decoder(16#23#));
reg_q1995_init <= '0' ;
	p_reg_q1995: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1995 <= reg_q1995_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1995 <= reg_q1995_init;
        else
          reg_q1995 <= reg_q1995_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2024_in <= (reg_q2022 AND symb_decoder(16#49#)) OR
 					(reg_q2022 AND symb_decoder(16#69#));
reg_q2024_init <= '0' ;
	p_reg_q2024: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2024 <= reg_q2024_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2024 <= reg_q2024_init;
        else
          reg_q2024 <= reg_q2024_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1934_in <= (reg_q1932 AND symb_decoder(16#45#)) OR
 					(reg_q1932 AND symb_decoder(16#65#));
reg_q1934_init <= '0' ;
	p_reg_q1934: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1934 <= reg_q1934_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1934 <= reg_q1934_init;
        else
          reg_q1934 <= reg_q1934_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q375_in <= (reg_q373 AND symb_decoder(16#54#)) OR
 					(reg_q373 AND symb_decoder(16#74#));
reg_q375_init <= '0' ;
	p_reg_q375: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q375 <= reg_q375_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q375 <= reg_q375_init;
        else
          reg_q375 <= reg_q375_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2472_in <= (reg_q2470 AND symb_decoder(16#4f#));
reg_q2472_init <= '0' ;
	p_reg_q2472: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2472 <= reg_q2472_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2472 <= reg_q2472_init;
        else
          reg_q2472 <= reg_q2472_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2628_in <= (reg_q2626 AND symb_decoder(16#74#)) OR
 					(reg_q2626 AND symb_decoder(16#54#));
reg_q2628_init <= '0' ;
	p_reg_q2628: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2628 <= reg_q2628_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2628 <= reg_q2628_init;
        else
          reg_q2628 <= reg_q2628_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q292_in <= (reg_q290 AND symb_decoder(16#4c#)) OR
 					(reg_q290 AND symb_decoder(16#6c#));
reg_q292_init <= '0' ;
	p_reg_q292: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q292 <= reg_q292_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q292 <= reg_q292_init;
        else
          reg_q292 <= reg_q292_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1702_in <= (reg_q1700 AND symb_decoder(16#64#)) OR
 					(reg_q1700 AND symb_decoder(16#44#));
reg_q1702_init <= '0' ;
	p_reg_q1702: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1702 <= reg_q1702_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1702 <= reg_q1702_init;
        else
          reg_q1702 <= reg_q1702_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1704_in <= (reg_q1702 AND symb_decoder(16#45#)) OR
 					(reg_q1702 AND symb_decoder(16#65#));
reg_q1704_init <= '0' ;
	p_reg_q1704: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1704 <= reg_q1704_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1704 <= reg_q1704_init;
        else
          reg_q1704 <= reg_q1704_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2491_in <= (reg_q2489 AND symb_decoder(16#52#));
reg_q2491_init <= '0' ;
	p_reg_q2491: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2491 <= reg_q2491_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2491 <= reg_q2491_init;
        else
          reg_q2491 <= reg_q2491_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2493_in <= (reg_q2491 AND symb_decoder(16#54#));
reg_q2493_init <= '0' ;
	p_reg_q2493: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2493 <= reg_q2493_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2493 <= reg_q2493_init;
        else
          reg_q2493 <= reg_q2493_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2451_in <= (reg_q2449 AND symb_decoder(16#32#));
reg_q2451_init <= '0' ;
	p_reg_q2451: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2451 <= reg_q2451_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2451 <= reg_q2451_init;
        else
          reg_q2451 <= reg_q2451_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2453_in <= (reg_q2451 AND symb_decoder(16#23#));
reg_q2453_init <= '0' ;
	p_reg_q2453: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2453 <= reg_q2453_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2453 <= reg_q2453_init;
        else
          reg_q2453 <= reg_q2453_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1722_in <= (reg_q1720 AND symb_decoder(16#59#)) OR
 					(reg_q1720 AND symb_decoder(16#79#));
reg_q1722_init <= '0' ;
	p_reg_q1722: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1722 <= reg_q1722_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1722 <= reg_q1722_init;
        else
          reg_q1722 <= reg_q1722_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1724_in <= (reg_q1722 AND symb_decoder(16#6f#)) OR
 					(reg_q1722 AND symb_decoder(16#4f#));
reg_q1724_init <= '0' ;
	p_reg_q1724: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1724 <= reg_q1724_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1724 <= reg_q1724_init;
        else
          reg_q1724 <= reg_q1724_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2101_in <= (reg_q2099 AND symb_decoder(16#61#)) OR
 					(reg_q2099 AND symb_decoder(16#41#));
reg_q2101_init <= '0' ;
	p_reg_q2101: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2101 <= reg_q2101_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2101 <= reg_q2101_init;
        else
          reg_q2101 <= reg_q2101_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1510_in <= (reg_q1508 AND symb_decoder(16#72#)) OR
 					(reg_q1508 AND symb_decoder(16#52#));
reg_q1510_init <= '0' ;
	p_reg_q1510: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1510 <= reg_q1510_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1510 <= reg_q1510_init;
        else
          reg_q1510 <= reg_q1510_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1512_in <= (reg_q1510 AND symb_decoder(16#73#)) OR
 					(reg_q1510 AND symb_decoder(16#53#));
reg_q1512_init <= '0' ;
	p_reg_q1512: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1512 <= reg_q1512_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1512 <= reg_q1512_init;
        else
          reg_q1512 <= reg_q1512_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1607_in <= (reg_q1605 AND symb_decoder(16#49#)) OR
 					(reg_q1605 AND symb_decoder(16#69#));
reg_q1607_init <= '0' ;
	p_reg_q1607: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1607 <= reg_q1607_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1607 <= reg_q1607_init;
        else
          reg_q1607 <= reg_q1607_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q720_in <= (reg_q718 AND symb_decoder(16#67#)) OR
 					(reg_q718 AND symb_decoder(16#47#));
reg_q720_init <= '0' ;
	p_reg_q720: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q720 <= reg_q720_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q720 <= reg_q720_init;
        else
          reg_q720 <= reg_q720_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q722_in <= (reg_q720 AND symb_decoder(16#65#)) OR
 					(reg_q720 AND symb_decoder(16#45#));
reg_q722_init <= '0' ;
	p_reg_q722: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q722 <= reg_q722_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q722 <= reg_q722_init;
        else
          reg_q722 <= reg_q722_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1572_in <= (reg_q1570 AND symb_decoder(16#6e#)) OR
 					(reg_q1570 AND symb_decoder(16#4e#));
reg_q1572_init <= '0' ;
	p_reg_q1572: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1572 <= reg_q1572_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1572 <= reg_q1572_init;
        else
          reg_q1572 <= reg_q1572_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q562_in <= (reg_q560 AND symb_decoder(16#64#)) OR
 					(reg_q560 AND symb_decoder(16#44#));
reg_q562_init <= '0' ;
	p_reg_q562: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q562 <= reg_q562_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q562 <= reg_q562_init;
        else
          reg_q562 <= reg_q562_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q564_in <= (reg_q562 AND symb_decoder(16#79#)) OR
 					(reg_q562 AND symb_decoder(16#59#));
reg_q564_init <= '0' ;
	p_reg_q564: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q564 <= reg_q564_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q564 <= reg_q564_init;
        else
          reg_q564 <= reg_q564_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1680_in <= (reg_q1678 AND symb_decoder(16#72#)) OR
 					(reg_q1678 AND symb_decoder(16#52#));
reg_q1680_init <= '0' ;
	p_reg_q1680: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1680 <= reg_q1680_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1680 <= reg_q1680_init;
        else
          reg_q1680 <= reg_q1680_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q736_in <= (reg_q734 AND symb_decoder(16#63#)) OR
 					(reg_q734 AND symb_decoder(16#43#));
reg_q736_init <= '0' ;
	p_reg_q736: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q736 <= reg_q736_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q736 <= reg_q736_init;
        else
          reg_q736 <= reg_q736_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q738_in <= (reg_q736 AND symb_decoder(16#4f#)) OR
 					(reg_q736 AND symb_decoder(16#6f#));
reg_q738_init <= '0' ;
	p_reg_q738: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q738 <= reg_q738_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q738 <= reg_q738_init;
        else
          reg_q738 <= reg_q738_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q486_in <= (reg_q484 AND symb_decoder(16#30#));
reg_q486_init <= '0' ;
	p_reg_q486: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q486 <= reg_q486_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q486 <= reg_q486_init;
        else
          reg_q486 <= reg_q486_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q488_in <= (reg_q486 AND symb_decoder(16#25#));
reg_q488_init <= '0' ;
	p_reg_q488: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q488 <= reg_q488_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q488 <= reg_q488_init;
        else
          reg_q488 <= reg_q488_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2142_in <= (reg_q2140 AND symb_decoder(16#68#)) OR
 					(reg_q2140 AND symb_decoder(16#48#));
reg_q2142_init <= '0' ;
	p_reg_q2142: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2142 <= reg_q2142_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2142 <= reg_q2142_init;
        else
          reg_q2142 <= reg_q2142_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1276_in <= (reg_q1274 AND symb_decoder(16#4f#)) OR
 					(reg_q1274 AND symb_decoder(16#6f#));
reg_q1276_init <= '0' ;
	p_reg_q1276: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1276 <= reg_q1276_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1276 <= reg_q1276_init;
        else
          reg_q1276 <= reg_q1276_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2237_in <= (reg_q2235 AND symb_decoder(16#56#)) OR
 					(reg_q2235 AND symb_decoder(16#76#));
reg_q2237_init <= '0' ;
	p_reg_q2237: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2237 <= reg_q2237_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2237 <= reg_q2237_init;
        else
          reg_q2237 <= reg_q2237_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1890_in <= (reg_q1888 AND symb_decoder(16#41#)) OR
 					(reg_q1888 AND symb_decoder(16#61#));
reg_q1890_init <= '0' ;
	p_reg_q1890: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1890 <= reg_q1890_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1890 <= reg_q1890_init;
        else
          reg_q1890 <= reg_q1890_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2014_in <= (reg_q2012 AND symb_decoder(16#53#)) OR
 					(reg_q2012 AND symb_decoder(16#73#));
reg_q2014_init <= '0' ;
	p_reg_q2014: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2014 <= reg_q2014_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2014 <= reg_q2014_init;
        else
          reg_q2014 <= reg_q2014_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1305_in <= (reg_q1303 AND symb_decoder(16#4c#)) OR
 					(reg_q1303 AND symb_decoder(16#6c#));
reg_q1305_init <= '0' ;
	p_reg_q1305: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1305 <= reg_q1305_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1305 <= reg_q1305_init;
        else
          reg_q1305 <= reg_q1305_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2549_in <= (reg_q2547 AND symb_decoder(16#47#)) OR
 					(reg_q2547 AND symb_decoder(16#67#));
reg_q2549_init <= '0' ;
	p_reg_q2549: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2549 <= reg_q2549_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2549 <= reg_q2549_init;
        else
          reg_q2549 <= reg_q2549_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2551_in <= (reg_q2549 AND symb_decoder(16#49#)) OR
 					(reg_q2549 AND symb_decoder(16#69#));
reg_q2551_init <= '0' ;
	p_reg_q2551: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2551 <= reg_q2551_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2551 <= reg_q2551_init;
        else
          reg_q2551 <= reg_q2551_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1804_in <= (reg_q1802 AND symb_decoder(16#53#)) OR
 					(reg_q1802 AND symb_decoder(16#73#));
reg_q1804_init <= '0' ;
	p_reg_q1804: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1804 <= reg_q1804_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1804 <= reg_q1804_init;
        else
          reg_q1804 <= reg_q1804_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1098_in <= (reg_q1096 AND symb_decoder(16#70#)) OR
 					(reg_q1096 AND symb_decoder(16#50#));
reg_q1098_init <= '0' ;
	p_reg_q1098: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1098 <= reg_q1098_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1098 <= reg_q1098_init;
        else
          reg_q1098 <= reg_q1098_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2200_in <= (reg_q2198 AND symb_decoder(16#65#)) OR
 					(reg_q2198 AND symb_decoder(16#45#));
reg_q2200_init <= '0' ;
	p_reg_q2200: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2200 <= reg_q2200_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2200 <= reg_q2200_init;
        else
          reg_q2200 <= reg_q2200_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q182_in <= (reg_q180 AND symb_decoder(16#30#));
reg_q182_init <= '0' ;
	p_reg_q182: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q182 <= reg_q182_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q182 <= reg_q182_init;
        else
          reg_q182 <= reg_q182_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2567_in <= (reg_q2565 AND symb_decoder(16#6f#)) OR
 					(reg_q2565 AND symb_decoder(16#4f#));
reg_q2567_init <= '0' ;
	p_reg_q2567: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2567 <= reg_q2567_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2567 <= reg_q2567_init;
        else
          reg_q2567 <= reg_q2567_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q654_in <= (reg_q652 AND symb_decoder(16#32#));
reg_q654_init <= '0' ;
	p_reg_q654: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q654 <= reg_q654_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q654 <= reg_q654_init;
        else
          reg_q654 <= reg_q654_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q278_in <= (reg_q276 AND symb_decoder(16#45#)) OR
 					(reg_q276 AND symb_decoder(16#65#));
reg_q278_init <= '0' ;
	p_reg_q278: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q278 <= reg_q278_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q278 <= reg_q278_init;
        else
          reg_q278 <= reg_q278_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q280_in <= (reg_q278 AND symb_decoder(16#61#)) OR
 					(reg_q278 AND symb_decoder(16#41#));
reg_q280_init <= '0' ;
	p_reg_q280: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q280 <= reg_q280_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q280 <= reg_q280_init;
        else
          reg_q280 <= reg_q280_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q584_in <= (reg_q582 AND symb_decoder(16#31#));
reg_q584_init <= '0' ;
	p_reg_q584: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q584 <= reg_q584_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q584 <= reg_q584_init;
        else
          reg_q584 <= reg_q584_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1625_in <= (reg_q1623 AND symb_decoder(16#5f#));
reg_q1625_init <= '0' ;
	p_reg_q1625: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1625 <= reg_q1625_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1625 <= reg_q1625_init;
        else
          reg_q1625 <= reg_q1625_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1627_in <= (reg_q1625 AND symb_decoder(16#56#)) OR
 					(reg_q1625 AND symb_decoder(16#76#));
reg_q1627_init <= '0' ;
	p_reg_q1627: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1627 <= reg_q1627_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1627 <= reg_q1627_init;
        else
          reg_q1627 <= reg_q1627_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1441_in <= (reg_q1439 AND symb_decoder(16#59#)) OR
 					(reg_q1439 AND symb_decoder(16#79#));
reg_q1441_init <= '0' ;
	p_reg_q1441: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1441 <= reg_q1441_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1441 <= reg_q1441_init;
        else
          reg_q1441 <= reg_q1441_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q456_in <= (reg_q454 AND symb_decoder(16#4f#)) OR
 					(reg_q454 AND symb_decoder(16#6f#));
reg_q456_init <= '0' ;
	p_reg_q456: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q456 <= reg_q456_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q456 <= reg_q456_init;
        else
          reg_q456 <= reg_q456_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q458_in <= (reg_q456 AND symb_decoder(16#64#)) OR
 					(reg_q456 AND symb_decoder(16#44#));
reg_q458_init <= '0' ;
	p_reg_q458: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q458 <= reg_q458_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q458 <= reg_q458_init;
        else
          reg_q458 <= reg_q458_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1732_in <= (reg_q1730 AND symb_decoder(16#69#)) OR
 					(reg_q1730 AND symb_decoder(16#49#));
reg_q1732_init <= '0' ;
	p_reg_q1732: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1732 <= reg_q1732_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1732 <= reg_q1732_init;
        else
          reg_q1732 <= reg_q1732_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q4_in <= (reg_q2 AND symb_decoder(16#30#));
reg_q4_init <= '0' ;
	p_reg_q4: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q4 <= reg_q4_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q4 <= reg_q4_init;
        else
          reg_q4 <= reg_q4_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q212_in <= (reg_q210 AND symb_decoder(16#4d#)) OR
 					(reg_q210 AND symb_decoder(16#6d#));
reg_q212_init <= '0' ;
	p_reg_q212: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q212 <= reg_q212_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q212 <= reg_q212_init;
        else
          reg_q212 <= reg_q212_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2419_in <= (reg_q2417 AND symb_decoder(16#45#)) OR
 					(reg_q2417 AND symb_decoder(16#65#));
reg_q2419_init <= '0' ;
	p_reg_q2419: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2419 <= reg_q2419_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2419 <= reg_q2419_init;
        else
          reg_q2419 <= reg_q2419_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q276_in <= (reg_q274 AND symb_decoder(16#44#)) OR
 					(reg_q274 AND symb_decoder(16#64#));
reg_q276_init <= '0' ;
	p_reg_q276: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q276 <= reg_q276_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q276 <= reg_q276_init;
        else
          reg_q276 <= reg_q276_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q345_in <= (reg_q343 AND symb_decoder(16#6f#)) OR
 					(reg_q343 AND symb_decoder(16#4f#));
reg_q345_init <= '0' ;
	p_reg_q345: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q345 <= reg_q345_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q345 <= reg_q345_init;
        else
          reg_q345 <= reg_q345_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1290_in <= (reg_q1288 AND symb_decoder(16#2e#));
reg_q1290_init <= '0' ;
	p_reg_q1290: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1290 <= reg_q1290_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1290 <= reg_q1290_init;
        else
          reg_q1290 <= reg_q1290_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1292_in <= (reg_q1290 AND symb_decoder(16#2e#));
reg_q1292_init <= '0' ;
	p_reg_q1292: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1292 <= reg_q1292_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1292 <= reg_q1292_init;
        else
          reg_q1292 <= reg_q1292_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2078_in <= (reg_q2076 AND symb_decoder(16#65#));
reg_q2078_init <= '0' ;
	p_reg_q2078: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2078 <= reg_q2078_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2078 <= reg_q2078_init;
        else
          reg_q2078 <= reg_q2078_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2080_in <= (reg_q2078 AND symb_decoder(16#72#));
reg_q2080_init <= '0' ;
	p_reg_q2080: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2080 <= reg_q2080_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2080 <= reg_q2080_init;
        else
          reg_q2080 <= reg_q2080_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1830_in <= (reg_q1828 AND symb_decoder(16#43#)) OR
 					(reg_q1828 AND symb_decoder(16#63#));
reg_q1830_init <= '0' ;
	p_reg_q1830: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1830 <= reg_q1830_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1830 <= reg_q1830_init;
        else
          reg_q1830 <= reg_q1830_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1798_in <= (reg_q1796 AND symb_decoder(16#75#)) OR
 					(reg_q1796 AND symb_decoder(16#55#));
reg_q1798_init <= '0' ;
	p_reg_q1798: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1798 <= reg_q1798_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1798 <= reg_q1798_init;
        else
          reg_q1798 <= reg_q1798_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2020_in <= (reg_q2018 AND symb_decoder(16#72#)) OR
 					(reg_q2018 AND symb_decoder(16#52#));
reg_q2020_init <= '0' ;
	p_reg_q2020: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2020 <= reg_q2020_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2020 <= reg_q2020_init;
        else
          reg_q2020 <= reg_q2020_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2539_in <= (reg_q2537 AND symb_decoder(16#46#)) OR
 					(reg_q2537 AND symb_decoder(16#66#));
reg_q2539_init <= '0' ;
	p_reg_q2539: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2539 <= reg_q2539_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2539 <= reg_q2539_init;
        else
          reg_q2539 <= reg_q2539_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2541_in <= (reg_q2539 AND symb_decoder(16#4f#)) OR
 					(reg_q2539 AND symb_decoder(16#6f#));
reg_q2541_init <= '0' ;
	p_reg_q2541: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2541 <= reg_q2541_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2541 <= reg_q2541_init;
        else
          reg_q2541 <= reg_q2541_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2316_in <= (reg_q2314 AND symb_decoder(16#21#));
reg_q2316_init <= '0' ;
	p_reg_q2316: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2316 <= reg_q2316_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2316 <= reg_q2316_init;
        else
          reg_q2316 <= reg_q2316_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2318_in <= (reg_q2316 AND symb_decoder(16#21#));
reg_q2318_init <= '0' ;
	p_reg_q2318: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2318 <= reg_q2318_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2318 <= reg_q2318_init;
        else
          reg_q2318 <= reg_q2318_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q931_in <= (reg_q929 AND symb_decoder(16#52#)) OR
 					(reg_q929 AND symb_decoder(16#72#));
reg_q931_init <= '0' ;
	p_reg_q931: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q931 <= reg_q931_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q931 <= reg_q931_init;
        else
          reg_q931 <= reg_q931_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1629_in <= (reg_q1627 AND symb_decoder(16#69#)) OR
 					(reg_q1627 AND symb_decoder(16#49#));
reg_q1629_init <= '0' ;
	p_reg_q1629: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1629 <= reg_q1629_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1629 <= reg_q1629_init;
        else
          reg_q1629 <= reg_q1629_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2465_in <= (reg_q2463 AND symb_decoder(16#23#));
reg_q2465_init <= '0' ;
	p_reg_q2465: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2465 <= reg_q2465_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2465 <= reg_q2465_init;
        else
          reg_q2465 <= reg_q2465_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2056_in <= (reg_q2054 AND symb_decoder(16#68#));
reg_q2056_init <= '0' ;
	p_reg_q2056: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2056 <= reg_q2056_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2056 <= reg_q2056_init;
        else
          reg_q2056 <= reg_q2056_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2058_in <= (reg_q2056 AND symb_decoder(16#65#));
reg_q2058_init <= '0' ;
	p_reg_q2058: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2058 <= reg_q2058_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2058 <= reg_q2058_init;
        else
          reg_q2058 <= reg_q2058_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2022_in <= (reg_q2020 AND symb_decoder(16#52#)) OR
 					(reg_q2020 AND symb_decoder(16#72#));
reg_q2022_init <= '0' ;
	p_reg_q2022: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2022 <= reg_q2022_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2022 <= reg_q2022_init;
        else
          reg_q2022 <= reg_q2022_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1948_in <= (reg_q1946 AND symb_decoder(16#41#)) OR
 					(reg_q1946 AND symb_decoder(16#61#));
reg_q1948_init <= '0' ;
	p_reg_q1948: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1948 <= reg_q1948_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1948 <= reg_q1948_init;
        else
          reg_q1948 <= reg_q1948_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1950_in <= (reg_q1948 AND symb_decoder(16#52#)) OR
 					(reg_q1948 AND symb_decoder(16#72#));
reg_q1950_init <= '0' ;
	p_reg_q1950: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1950 <= reg_q1950_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1950 <= reg_q1950_init;
        else
          reg_q1950 <= reg_q1950_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2168_in <= (reg_q2166 AND symb_decoder(16#6d#)) OR
 					(reg_q2166 AND symb_decoder(16#4d#));
reg_q2168_init <= '0' ;
	p_reg_q2168: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2168 <= reg_q2168_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2168 <= reg_q2168_init;
        else
          reg_q2168 <= reg_q2168_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q636_in <= (reg_q634 AND symb_decoder(16#6e#)) OR
 					(reg_q634 AND symb_decoder(16#4e#));
reg_q636_init <= '0' ;
	p_reg_q636: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q636 <= reg_q636_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q636 <= reg_q636_init;
        else
          reg_q636 <= reg_q636_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1484_in <= (reg_q1482 AND symb_decoder(16#2d#));
reg_q1484_init <= '0' ;
	p_reg_q1484: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1484 <= reg_q1484_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1484 <= reg_q1484_init;
        else
          reg_q1484 <= reg_q1484_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q929_in <= (reg_q927 AND symb_decoder(16#45#)) OR
 					(reg_q927 AND symb_decoder(16#65#));
reg_q929_init <= '0' ;
	p_reg_q929: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q929 <= reg_q929_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q929 <= reg_q929_init;
        else
          reg_q929 <= reg_q929_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q460_in <= (reg_q458 AND symb_decoder(16#59#)) OR
 					(reg_q458 AND symb_decoder(16#79#));
reg_q460_init <= '0' ;
	p_reg_q460: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q460 <= reg_q460_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q460 <= reg_q460_init;
        else
          reg_q460 <= reg_q460_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1700_in <= (reg_q1698 AND symb_decoder(16#72#)) OR
 					(reg_q1698 AND symb_decoder(16#52#));
reg_q1700_init <= '0' ;
	p_reg_q1700: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1700 <= reg_q1700_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1700 <= reg_q1700_init;
        else
          reg_q1700 <= reg_q1700_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2084_in <= (reg_q2082 AND symb_decoder(16#65#));
reg_q2084_init <= '0' ;
	p_reg_q2084: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2084 <= reg_q2084_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2084 <= reg_q2084_init;
        else
          reg_q2084 <= reg_q2084_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2086_in <= (reg_q2084 AND symb_decoder(16#72#));
reg_q2086_init <= '0' ;
	p_reg_q2086: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2086 <= reg_q2086_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2086 <= reg_q2086_init;
        else
          reg_q2086 <= reg_q2086_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1474_in <= (reg_q1472 AND symb_decoder(16#45#)) OR
 					(reg_q1472 AND symb_decoder(16#65#));
reg_q1474_init <= '0' ;
	p_reg_q1474: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1474 <= reg_q1474_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1474 <= reg_q1474_init;
        else
          reg_q1474 <= reg_q1474_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1476_in <= (reg_q1474 AND symb_decoder(16#61#)) OR
 					(reg_q1474 AND symb_decoder(16#41#));
reg_q1476_init <= '0' ;
	p_reg_q1476: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1476 <= reg_q1476_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1476 <= reg_q1476_init;
        else
          reg_q1476 <= reg_q1476_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1052_in <= (reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q1051 AND symb_decoder(16#45#)) OR
 					(reg_q1051 AND symb_decoder(16#65#));
reg_q1052_init <= '0' ;
	p_reg_q1052: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1052 <= reg_q1052_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1052 <= reg_q1052_init;
        else
          reg_q1052 <= reg_q1052_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1054_in <= (reg_q1052 AND symb_decoder(16#58#)) OR
 					(reg_q1052 AND symb_decoder(16#78#));
reg_q1054_init <= '0' ;
	p_reg_q1054: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1054 <= reg_q1054_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1054 <= reg_q1054_init;
        else
          reg_q1054 <= reg_q1054_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2619_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2618 AND symb_decoder(16#0a#)) OR
 					(reg_q2618 AND symb_decoder(16#0d#));
reg_q2619_init <= '0' ;
	p_reg_q2619: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2619 <= reg_q2619_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2619 <= reg_q2619_init;
        else
          reg_q2619 <= reg_q2619_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1856_in <= (reg_q1854 AND symb_decoder(16#56#)) OR
 					(reg_q1854 AND symb_decoder(16#76#));
reg_q1856_init <= '0' ;
	p_reg_q1856: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1856 <= reg_q1856_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1856 <= reg_q1856_init;
        else
          reg_q1856 <= reg_q1856_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2363_in <= (reg_q2361 AND symb_decoder(16#45#)) OR
 					(reg_q2361 AND symb_decoder(16#65#));
reg_q2363_init <= '0' ;
	p_reg_q2363: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2363 <= reg_q2363_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2363 <= reg_q2363_init;
        else
          reg_q2363 <= reg_q2363_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2327_in <= (reg_q2325 AND symb_decoder(16#57#)) OR
 					(reg_q2325 AND symb_decoder(16#77#));
reg_q2327_init <= '0' ;
	p_reg_q2327: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2327 <= reg_q2327_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2327 <= reg_q2327_init;
        else
          reg_q2327 <= reg_q2327_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q222_in <= (reg_q220 AND symb_decoder(16#6e#)) OR
 					(reg_q220 AND symb_decoder(16#4e#));
reg_q222_init <= '0' ;
	p_reg_q222: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q222 <= reg_q222_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q222 <= reg_q222_init;
        else
          reg_q222 <= reg_q222_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1155_in <= (reg_q1153 AND symb_decoder(16#0a#));
reg_q1155_init <= '0' ;
	p_reg_q1155: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1155 <= reg_q1155_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1155 <= reg_q1155_init;
        else
          reg_q1155 <= reg_q1155_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1746_in <= (reg_q1744 AND symb_decoder(16#0c#)) OR
 					(reg_q1744 AND symb_decoder(16#0a#)) OR
 					(reg_q1744 AND symb_decoder(16#20#)) OR
 					(reg_q1744 AND symb_decoder(16#09#)) OR
 					(reg_q1744 AND symb_decoder(16#0d#));
reg_q1746_init <= '0' ;
	p_reg_q1746: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1746 <= reg_q1746_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1746 <= reg_q1746_init;
        else
          reg_q1746 <= reg_q1746_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1262_in <= (reg_q1260 AND symb_decoder(16#53#)) OR
 					(reg_q1260 AND symb_decoder(16#73#));
reg_q1262_init <= '0' ;
	p_reg_q1262: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1262 <= reg_q1262_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1262 <= reg_q1262_init;
        else
          reg_q1262 <= reg_q1262_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2389_in <= (reg_q2387 AND symb_decoder(16#23#));
reg_q2389_init <= '0' ;
	p_reg_q2389: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2389 <= reg_q2389_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2389 <= reg_q2389_init;
        else
          reg_q2389 <= reg_q2389_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2391_in <= (reg_q2389 AND symb_decoder(16#41#)) OR
 					(reg_q2389 AND symb_decoder(16#61#));
reg_q2391_init <= '0' ;
	p_reg_q2391: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2391 <= reg_q2391_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2391 <= reg_q2391_init;
        else
          reg_q2391 <= reg_q2391_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2359_in <= (reg_q2357 AND symb_decoder(16#61#)) OR
 					(reg_q2357 AND symb_decoder(16#41#));
reg_q2359_init <= '0' ;
	p_reg_q2359: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2359 <= reg_q2359_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2359 <= reg_q2359_init;
        else
          reg_q2359 <= reg_q2359_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1952_in <= (reg_q1950 AND symb_decoder(16#45#)) OR
 					(reg_q1950 AND symb_decoder(16#65#));
reg_q1952_init <= '0' ;
	p_reg_q1952: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1952 <= reg_q1952_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1952 <= reg_q1952_init;
        else
          reg_q1952 <= reg_q1952_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2563_in <= (reg_q2561 AND symb_decoder(16#44#)) OR
 					(reg_q2561 AND symb_decoder(16#64#));
reg_q2563_init <= '0' ;
	p_reg_q2563: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2563 <= reg_q2563_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2563 <= reg_q2563_init;
        else
          reg_q2563 <= reg_q2563_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2593_in <= (reg_q2591 AND symb_decoder(16#72#)) OR
 					(reg_q2591 AND symb_decoder(16#52#));
reg_q2593_init <= '0' ;
	p_reg_q2593: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2593 <= reg_q2593_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2593 <= reg_q2593_init;
        else
          reg_q2593 <= reg_q2593_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2595_in <= (reg_q2593 AND symb_decoder(16#65#)) OR
 					(reg_q2593 AND symb_decoder(16#45#));
reg_q2595_init <= '0' ;
	p_reg_q2595: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2595 <= reg_q2595_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2595 <= reg_q2595_init;
        else
          reg_q2595 <= reg_q2595_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q313_in <= (reg_q311 AND symb_decoder(16#65#)) OR
 					(reg_q311 AND symb_decoder(16#45#));
reg_q313_init <= '0' ;
	p_reg_q313: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q313 <= reg_q313_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q313 <= reg_q313_init;
        else
          reg_q313 <= reg_q313_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q315_in <= (reg_q313 AND symb_decoder(16#52#)) OR
 					(reg_q313 AND symb_decoder(16#72#));
reg_q315_init <= '0' ;
	p_reg_q315: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q315 <= reg_q315_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q315 <= reg_q315_init;
        else
          reg_q315 <= reg_q315_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q576_in <= (reg_q574 AND symb_decoder(16#32#));
reg_q576_init <= '0' ;
	p_reg_q576: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q576 <= reg_q576_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q576 <= reg_q576_init;
        else
          reg_q576 <= reg_q576_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q578_in <= (reg_q576 AND symb_decoder(16#31#));
reg_q578_init <= '0' ;
	p_reg_q578: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q578 <= reg_q578_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q578 <= reg_q578_init;
        else
          reg_q578 <= reg_q578_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1472_in <= (reg_q1470 AND symb_decoder(16#52#)) OR
 					(reg_q1470 AND symb_decoder(16#72#));
reg_q1472_init <= '0' ;
	p_reg_q1472: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1472 <= reg_q1472_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1472 <= reg_q1472_init;
        else
          reg_q1472 <= reg_q1472_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2603_in <= (reg_q2601 AND symb_decoder(16#55#)) OR
 					(reg_q2601 AND symb_decoder(16#75#));
reg_q2603_init <= '0' ;
	p_reg_q2603: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2603 <= reg_q2603_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2603 <= reg_q2603_init;
        else
          reg_q2603 <= reg_q2603_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1588_in <= (reg_q1586 AND symb_decoder(16#65#)) OR
 					(reg_q1586 AND symb_decoder(16#45#));
reg_q1588_init <= '0' ;
	p_reg_q1588: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1588 <= reg_q1588_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1588 <= reg_q1588_init;
        else
          reg_q1588 <= reg_q1588_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2076_in <= (reg_q2074 AND symb_decoder(16#53#));
reg_q2076_init <= '0' ;
	p_reg_q2076: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2076 <= reg_q2076_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2076 <= reg_q2076_init;
        else
          reg_q2076 <= reg_q2076_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2206_in <= (reg_q2204 AND symb_decoder(16#6e#)) OR
 					(reg_q2204 AND symb_decoder(16#4e#));
reg_q2206_init <= '0' ;
	p_reg_q2206: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2206 <= reg_q2206_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2206 <= reg_q2206_init;
        else
          reg_q2206 <= reg_q2206_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2212_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2211 AND symb_decoder(16#0a#)) OR
 					(reg_q2211 AND symb_decoder(16#0d#));
reg_q2212_init <= '0' ;
	p_reg_q2212: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2212 <= reg_q2212_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2212 <= reg_q2212_init;
        else
          reg_q2212 <= reg_q2212_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2006_in <= (reg_q2004 AND symb_decoder(16#54#)) OR
 					(reg_q2004 AND symb_decoder(16#74#));
reg_q2006_init <= '0' ;
	p_reg_q2006: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2006 <= reg_q2006_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2006 <= reg_q2006_init;
        else
          reg_q2006 <= reg_q2006_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2008_in <= (reg_q2006 AND symb_decoder(16#72#)) OR
 					(reg_q2006 AND symb_decoder(16#52#));
reg_q2008_init <= '0' ;
	p_reg_q2008: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2008 <= reg_q2008_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2008 <= reg_q2008_init;
        else
          reg_q2008 <= reg_q2008_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q355_in <= (reg_q353 AND symb_decoder(16#72#)) OR
 					(reg_q353 AND symb_decoder(16#52#));
reg_q355_init <= '0' ;
	p_reg_q355: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q355 <= reg_q355_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q355 <= reg_q355_init;
        else
          reg_q355 <= reg_q355_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1074_in <= (reg_q1072 AND symb_decoder(16#65#)) OR
 					(reg_q1072 AND symb_decoder(16#45#));
reg_q1074_init <= '0' ;
	p_reg_q1074: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1074 <= reg_q1074_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1074 <= reg_q1074_init;
        else
          reg_q1074 <= reg_q1074_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2225_in <= (reg_q2223 AND symb_decoder(16#53#)) OR
 					(reg_q2223 AND symb_decoder(16#73#));
reg_q2225_init <= '0' ;
	p_reg_q2225: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2225 <= reg_q2225_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2225 <= reg_q2225_init;
        else
          reg_q2225 <= reg_q2225_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1385_in <= (reg_q1383 AND symb_decoder(16#6e#)) OR
 					(reg_q1383 AND symb_decoder(16#4e#));
reg_q1385_init <= '0' ;
	p_reg_q1385: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1385 <= reg_q1385_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1385 <= reg_q1385_init;
        else
          reg_q1385 <= reg_q1385_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1119_in <= (reg_q1117 AND symb_decoder(16#63#)) OR
 					(reg_q1117 AND symb_decoder(16#43#));
reg_q1119_init <= '0' ;
	p_reg_q1119: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1119 <= reg_q1119_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1119 <= reg_q1119_init;
        else
          reg_q1119 <= reg_q1119_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q274_in <= (reg_q272 AND symb_decoder(16#20#));
reg_q274_init <= '0' ;
	p_reg_q274: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q274 <= reg_q274_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q274 <= reg_q274_init;
        else
          reg_q274 <= reg_q274_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q650_in <= (reg_q648 AND symb_decoder(16#31#));
reg_q650_init <= '0' ;
	p_reg_q650: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q650 <= reg_q650_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q650 <= reg_q650_init;
        else
          reg_q650 <= reg_q650_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q652_in <= (reg_q650 AND symb_decoder(16#25#));
reg_q652_init <= '0' ;
	p_reg_q652: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q652 <= reg_q652_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q652 <= reg_q652_init;
        else
          reg_q652 <= reg_q652_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2609_in <= (reg_q2607 AND symb_decoder(16#72#)) OR
 					(reg_q2607 AND symb_decoder(16#52#));
reg_q2609_init <= '0' ;
	p_reg_q2609: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2609 <= reg_q2609_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2609 <= reg_q2609_init;
        else
          reg_q2609 <= reg_q2609_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1635_in <= (reg_q1633 AND symb_decoder(16#69#)) OR
 					(reg_q1633 AND symb_decoder(16#49#));
reg_q1635_init <= '0' ;
	p_reg_q1635: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1635 <= reg_q1635_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1635 <= reg_q1635_init;
        else
          reg_q1635 <= reg_q1635_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q667_in <= (reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q666 AND symb_decoder(16#42#)) OR
 					(reg_q666 AND symb_decoder(16#62#));
reg_q667_init <= '0' ;
	p_reg_q667: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q667 <= reg_q667_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q667 <= reg_q667_init;
        else
          reg_q667 <= reg_q667_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1912_in <= (reg_q1910 AND symb_decoder(16#6f#)) OR
 					(reg_q1910 AND symb_decoder(16#4f#));
reg_q1912_init <= '0' ;
	p_reg_q1912: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1912 <= reg_q1912_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1912 <= reg_q1912_init;
        else
          reg_q1912 <= reg_q1912_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1514_in <= (reg_q1512 AND symb_decoder(16#69#)) OR
 					(reg_q1512 AND symb_decoder(16#49#));
reg_q1514_init <= '0' ;
	p_reg_q1514: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1514 <= reg_q1514_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1514 <= reg_q1514_init;
        else
          reg_q1514 <= reg_q1514_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1516_in <= (reg_q1514 AND symb_decoder(16#4f#)) OR
 					(reg_q1514 AND symb_decoder(16#6f#));
reg_q1516_init <= '0' ;
	p_reg_q1516: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1516 <= reg_q1516_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1516 <= reg_q1516_init;
        else
          reg_q1516 <= reg_q1516_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1940_in <= (reg_q1938 AND symb_decoder(16#53#)) OR
 					(reg_q1938 AND symb_decoder(16#73#));
reg_q1940_init <= '0' ;
	p_reg_q1940: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1940 <= reg_q1940_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1940 <= reg_q1940_init;
        else
          reg_q1940 <= reg_q1940_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1100_in <= (reg_q1098 AND symb_decoder(16#4f#)) OR
 					(reg_q1098 AND symb_decoder(16#6f#));
reg_q1100_init <= '0' ;
	p_reg_q1100: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1100 <= reg_q1100_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1100 <= reg_q1100_init;
        else
          reg_q1100 <= reg_q1100_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q227_in <= (reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q226 AND symb_decoder(16#36#));
reg_q227_init <= '0' ;
	p_reg_q227: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q227 <= reg_q227_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q227 <= reg_q227_init;
        else
          reg_q227 <= reg_q227_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q506_in <= (reg_q504 AND symb_decoder(16#3a#));
reg_q506_init <= '0' ;
	p_reg_q506: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q506 <= reg_q506_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q506 <= reg_q506_init;
        else
          reg_q506 <= reg_q506_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q682_in <= (reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q681 AND symb_decoder(16#43#)) OR
 					(reg_q681 AND symb_decoder(16#63#));
reg_q682_init <= '0' ;
	p_reg_q682: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q682 <= reg_q682_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q682 <= reg_q682_init;
        else
          reg_q682 <= reg_q682_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1021_in <= (reg_q1019 AND symb_decoder(16#7a#)) OR
 					(reg_q1019 AND symb_decoder(16#5a#));
reg_q1021_init <= '0' ;
	p_reg_q1021: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1021 <= reg_q1021_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1021 <= reg_q1021_init;
        else
          reg_q1021 <= reg_q1021_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q190_in <= (reg_q188 AND symb_decoder(16#33#));
reg_q190_init <= '0' ;
	p_reg_q190: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q190 <= reg_q190_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q190 <= reg_q190_init;
        else
          reg_q190 <= reg_q190_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q192_in <= (reg_q190 AND symb_decoder(16#41#)) OR
 					(reg_q190 AND symb_decoder(16#61#));
reg_q192_init <= '0' ;
	p_reg_q192: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q192 <= reg_q192_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q192 <= reg_q192_init;
        else
          reg_q192 <= reg_q192_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2433_in <= (reg_q2431 AND symb_decoder(16#4e#)) OR
 					(reg_q2431 AND symb_decoder(16#6e#));
reg_q2433_init <= '0' ;
	p_reg_q2433: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2433 <= reg_q2433_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2433 <= reg_q2433_init;
        else
          reg_q2433 <= reg_q2433_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q921_in <= (reg_q919 AND symb_decoder(16#73#)) OR
 					(reg_q919 AND symb_decoder(16#53#));
reg_q921_init <= '0' ;
	p_reg_q921: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q921 <= reg_q921_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q921 <= reg_q921_init;
        else
          reg_q921 <= reg_q921_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1278_in <= (reg_q1276 AND symb_decoder(16#4e#)) OR
 					(reg_q1276 AND symb_decoder(16#6e#));
reg_q1278_init <= '0' ;
	p_reg_q1278: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1278 <= reg_q1278_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1278 <= reg_q1278_init;
        else
          reg_q1278 <= reg_q1278_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q214_in <= (reg_q212 AND symb_decoder(16#45#)) OR
 					(reg_q212 AND symb_decoder(16#65#));
reg_q214_init <= '0' ;
	p_reg_q214: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q214 <= reg_q214_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q214 <= reg_q214_init;
        else
          reg_q214 <= reg_q214_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q347_in <= (reg_q345 AND symb_decoder(16#6c#)) OR
 					(reg_q345 AND symb_decoder(16#4c#));
reg_q347_init <= '0' ;
	p_reg_q347: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q347 <= reg_q347_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q347 <= reg_q347_init;
        else
          reg_q347 <= reg_q347_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2664_in <= (reg_q2662 AND symb_decoder(16#67#)) OR
 					(reg_q2662 AND symb_decoder(16#47#));
reg_q2664_init <= '0' ;
	p_reg_q2664: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2664 <= reg_q2664_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2664 <= reg_q2664_init;
        else
          reg_q2664 <= reg_q2664_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2676_in <= (reg_q2674 AND symb_decoder(16#73#)) OR
 					(reg_q2674 AND symb_decoder(16#53#));
reg_q2676_init <= '0' ;
	p_reg_q2676: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2676 <= reg_q2676_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2676 <= reg_q2676_init;
        else
          reg_q2676 <= reg_q2676_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2666_in <= (reg_q2664 AND symb_decoder(16#47#)) OR
 					(reg_q2664 AND symb_decoder(16#67#));
reg_q2666_init <= '0' ;
	p_reg_q2666: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2666 <= reg_q2666_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2666 <= reg_q2666_init;
        else
          reg_q2666 <= reg_q2666_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q428_in <= (reg_q426 AND symb_decoder(16#72#)) OR
 					(reg_q426 AND symb_decoder(16#52#));
reg_q428_init <= '0' ;
	p_reg_q428: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q428 <= reg_q428_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q428 <= reg_q428_init;
        else
          reg_q428 <= reg_q428_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2485_in <= (reg_q2695 AND symb_decoder(16#2a#));
reg_q2485_init <= '0' ;
	p_reg_q2485: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2485 <= reg_q2485_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2485 <= reg_q2485_init;
        else
          reg_q2485 <= reg_q2485_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1637_in <= (reg_q1635 AND symb_decoder(16#6d#)) OR
 					(reg_q1635 AND symb_decoder(16#4d#));
reg_q1637_init <= '0' ;
	p_reg_q1637: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1637 <= reg_q1637_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1637 <= reg_q1637_init;
        else
          reg_q1637 <= reg_q1637_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2361_in <= (reg_q2359 AND symb_decoder(16#67#)) OR
 					(reg_q2359 AND symb_decoder(16#47#));
reg_q2361_init <= '0' ;
	p_reg_q2361: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2361 <= reg_q2361_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2361 <= reg_q2361_init;
        else
          reg_q2361 <= reg_q2361_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1187_in <= (reg_q1185 AND symb_decoder(16#41#)) OR
 					(reg_q1185 AND symb_decoder(16#61#));
reg_q1187_init <= '0' ;
	p_reg_q1187: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1187 <= reg_q1187_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1187 <= reg_q1187_init;
        else
          reg_q1187 <= reg_q1187_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1294_in <= (reg_q1292 AND symb_decoder(16#2e#));
reg_q1294_init <= '0' ;
	p_reg_q1294: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1294 <= reg_q1294_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1294 <= reg_q1294_init;
        else
          reg_q1294 <= reg_q1294_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q478_in <= (reg_q476 AND symb_decoder(16#30#));
reg_q478_init <= '0' ;
	p_reg_q478: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q478 <= reg_q478_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q478 <= reg_q478_init;
        else
          reg_q478 <= reg_q478_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1864_in <= (reg_q1862 AND symb_decoder(16#72#)) OR
 					(reg_q1862 AND symb_decoder(16#52#));
reg_q1864_init <= '0' ;
	p_reg_q1864: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1864 <= reg_q1864_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1864 <= reg_q1864_init;
        else
          reg_q1864 <= reg_q1864_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1203_in <= (reg_q1201 AND symb_decoder(16#4f#)) OR
 					(reg_q1201 AND symb_decoder(16#6f#));
reg_q1203_init <= '0' ;
	p_reg_q1203: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1203 <= reg_q1203_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1203 <= reg_q1203_init;
        else
          reg_q1203 <= reg_q1203_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q500_in <= (reg_q498 AND symb_decoder(16#69#)) OR
 					(reg_q498 AND symb_decoder(16#49#));
reg_q500_init <= '0' ;
	p_reg_q500: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q500 <= reg_q500_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q500 <= reg_q500_init;
        else
          reg_q500 <= reg_q500_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q998_in <= (reg_q996 AND symb_decoder(16#74#)) OR
 					(reg_q996 AND symb_decoder(16#54#));
reg_q998_init <= '0' ;
	p_reg_q998: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q998 <= reg_q998_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q998 <= reg_q998_init;
        else
          reg_q998 <= reg_q998_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q171_in <= (reg_q169 AND symb_decoder(16#6c#)) OR
 					(reg_q169 AND symb_decoder(16#4c#));
reg_q171_init <= '0' ;
	p_reg_q171: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q171 <= reg_q171_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q171 <= reg_q171_init;
        else
          reg_q171 <= reg_q171_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2561_in <= (reg_q2559 AND symb_decoder(16#45#)) OR
 					(reg_q2559 AND symb_decoder(16#65#));
reg_q2561_init <= '0' ;
	p_reg_q2561: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2561 <= reg_q2561_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2561 <= reg_q2561_init;
        else
          reg_q2561 <= reg_q2561_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1586_in <= (reg_q1584 AND symb_decoder(16#53#)) OR
 					(reg_q1584 AND symb_decoder(16#73#));
reg_q1586_init <= '0' ;
	p_reg_q1586: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1586 <= reg_q1586_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1586 <= reg_q1586_init;
        else
          reg_q1586 <= reg_q1586_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2320_in <= (reg_q2318 AND symb_decoder(16#21#));
reg_q2320_init <= '0' ;
	p_reg_q2320: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2320 <= reg_q2320_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2320 <= reg_q2320_init;
        else
          reg_q2320 <= reg_q2320_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q42_in <= (reg_q40 AND symb_decoder(16#2e#));
reg_q42_init <= '0' ;
	p_reg_q42: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q42 <= reg_q42_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q42 <= reg_q42_init;
        else
          reg_q42 <= reg_q42_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q44_in <= (reg_q42 AND symb_decoder(16#2e#));
reg_q44_init <= '0' ;
	p_reg_q44: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q44 <= reg_q44_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q44 <= reg_q44_init;
        else
          reg_q44 <= reg_q44_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1518_in <= (reg_q1516 AND symb_decoder(16#6e#)) OR
 					(reg_q1516 AND symb_decoder(16#4e#));
reg_q1518_init <= '0' ;
	p_reg_q1518: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1518 <= reg_q1518_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1518 <= reg_q1518_init;
        else
          reg_q1518 <= reg_q1518_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2626_in <= (reg_q2624 AND symb_decoder(16#41#)) OR
 					(reg_q2624 AND symb_decoder(16#61#));
reg_q2626_init <= '0' ;
	p_reg_q2626: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2626 <= reg_q2626_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2626 <= reg_q2626_init;
        else
          reg_q2626 <= reg_q2626_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2589_in <= (reg_q2587 AND symb_decoder(16#55#)) OR
 					(reg_q2587 AND symb_decoder(16#75#));
reg_q2589_init <= '0' ;
	p_reg_q2589: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2589 <= reg_q2589_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2589 <= reg_q2589_init;
        else
          reg_q2589 <= reg_q2589_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2591_in <= (reg_q2589 AND symb_decoder(16#52#)) OR
 					(reg_q2589 AND symb_decoder(16#72#));
reg_q2591_init <= '0' ;
	p_reg_q2591: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2591 <= reg_q2591_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2591 <= reg_q2591_init;
        else
          reg_q2591 <= reg_q2591_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1870_in <= (reg_q1868 AND symb_decoder(16#50#)) OR
 					(reg_q1868 AND symb_decoder(16#70#));
reg_q1870_init <= '0' ;
	p_reg_q1870: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1870 <= reg_q1870_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1870 <= reg_q1870_init;
        else
          reg_q1870 <= reg_q1870_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1157_in <= (reg_q1155 AND symb_decoder(16#0d#));
reg_q1157_init <= '0' ;
	p_reg_q1157: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1157 <= reg_q1157_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1157 <= reg_q1157_init;
        else
          reg_q1157 <= reg_q1157_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q776_in <= (reg_q774 AND symb_decoder(16#3a#));
reg_q776_init <= '0' ;
	p_reg_q776: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q776 <= reg_q776_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q776 <= reg_q776_init;
        else
          reg_q776 <= reg_q776_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2186_in <= (reg_q2184 AND symb_decoder(16#6f#)) OR
 					(reg_q2184 AND symb_decoder(16#4f#));
reg_q2186_init <= '0' ;
	p_reg_q2186: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2186 <= reg_q2186_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2186 <= reg_q2186_init;
        else
          reg_q2186 <= reg_q2186_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q480_in <= (reg_q478 AND symb_decoder(16#2e#));
reg_q480_init <= '0' ;
	p_reg_q480: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q480 <= reg_q480_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q480 <= reg_q480_init;
        else
          reg_q480 <= reg_q480_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q97_in <= (reg_q95 AND symb_decoder(16#31#));
reg_q97_init <= '0' ;
	p_reg_q97: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q97 <= reg_q97_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q97 <= reg_q97_init;
        else
          reg_q97 <= reg_q97_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1080_in <= (reg_q1078 AND symb_decoder(16#65#)) OR
 					(reg_q1078 AND symb_decoder(16#45#));
reg_q1080_init <= '0' ;
	p_reg_q1080: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1080 <= reg_q1080_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1080 <= reg_q1080_init;
        else
          reg_q1080 <= reg_q1080_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1121_in <= (reg_q1119 AND symb_decoder(16#65#)) OR
 					(reg_q1119 AND symb_decoder(16#45#));
reg_q1121_init <= '0' ;
	p_reg_q1121: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1121 <= reg_q1121_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1121 <= reg_q1121_init;
        else
          reg_q1121 <= reg_q1121_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1486_in <= (reg_q1484 AND symb_decoder(16#5c#));
reg_q1486_init <= '0' ;
	p_reg_q1486: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1486 <= reg_q1486_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1486 <= reg_q1486_init;
        else
          reg_q1486 <= reg_q1486_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2082_in <= (reg_q2080 AND symb_decoder(16#76#));
reg_q2082_init <= '0' ;
	p_reg_q2082: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2082 <= reg_q2082_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2082 <= reg_q2082_init;
        else
          reg_q2082 <= reg_q2082_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q492_in <= (reg_q490 AND symb_decoder(16#30#));
reg_q492_init <= '0' ;
	p_reg_q492: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q492 <= reg_q492_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q492 <= reg_q492_init;
        else
          reg_q492 <= reg_q492_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q544_in <= (reg_q542 AND symb_decoder(16#5b#));
reg_q544_init <= '0' ;
	p_reg_q544: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q544 <= reg_q544_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q544 <= reg_q544_init;
        else
          reg_q544 <= reg_q544_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2099_in <= (reg_q2097 AND symb_decoder(16#69#)) OR
 					(reg_q2097 AND symb_decoder(16#49#));
reg_q2099_init <= '0' ;
	p_reg_q2099: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2099 <= reg_q2099_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2099 <= reg_q2099_init;
        else
          reg_q2099 <= reg_q2099_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q216_in <= (reg_q214 AND symb_decoder(16#52#)) OR
 					(reg_q214 AND symb_decoder(16#72#));
reg_q216_init <= '0' ;
	p_reg_q216: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q216 <= reg_q216_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q216 <= reg_q216_init;
        else
          reg_q216 <= reg_q216_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1639_in <= (reg_q1637 AND symb_decoder(16#0d#));
reg_q1639_init <= '0' ;
	p_reg_q1639: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1639 <= reg_q1639_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1639 <= reg_q1639_init;
        else
          reg_q1639 <= reg_q1639_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2393_in <= (reg_q2391 AND symb_decoder(16#63#)) OR
 					(reg_q2391 AND symb_decoder(16#43#));
reg_q2393_init <= '0' ;
	p_reg_q2393: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2393 <= reg_q2393_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2393 <= reg_q2393_init;
        else
          reg_q2393 <= reg_q2393_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q542_in <= (reg_q540 AND symb_decoder(16#30#));
reg_q542_init <= '0' ;
	p_reg_q542: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q542 <= reg_q542_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q542 <= reg_q542_init;
        else
          reg_q542 <= reg_q542_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2504_in <= (reg_q2502 AND symb_decoder(16#50#));
reg_q2504_init <= '0' ;
	p_reg_q2504: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2504 <= reg_q2504_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2504 <= reg_q2504_init;
        else
          reg_q2504 <= reg_q2504_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1066_in <= (reg_q1064 AND symb_decoder(16#65#)) OR
 					(reg_q1064 AND symb_decoder(16#45#));
reg_q1066_init <= '0' ;
	p_reg_q1066: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1066 <= reg_q1066_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1066 <= reg_q1066_init;
        else
          reg_q1066 <= reg_q1066_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q180_in <= (reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q179 AND symb_decoder(16#31#));
reg_q180_init <= '0' ;
	p_reg_q180: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q180 <= reg_q180_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q180 <= reg_q180_init;
        else
          reg_q180 <= reg_q180_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q574_in <= (reg_q572 AND symb_decoder(16#25#));
reg_q574_init <= '0' ;
	p_reg_q574: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q574 <= reg_q574_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q574 <= reg_q574_init;
        else
          reg_q574 <= reg_q574_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q272_in <= (reg_q270 AND symb_decoder(16#31#));
reg_q272_init <= '0' ;
	p_reg_q272: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q272 <= reg_q272_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q272 <= reg_q272_init;
        else
          reg_q272 <= reg_q272_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1010_in <= (reg_q1008 AND symb_decoder(16#0a#));
reg_q1010_init <= '0' ;
	p_reg_q1010: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1010 <= reg_q1010_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1010 <= reg_q1010_init;
        else
          reg_q1010 <= reg_q1010_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q508_in <= (reg_q506 AND symb_decoder(16#25#));
reg_q508_init <= '0' ;
	p_reg_q508: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q508 <= reg_q508_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q508 <= reg_q508_init;
        else
          reg_q508 <= reg_q508_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q259_in <= (reg_q257 AND symb_decoder(16#ff#));
reg_q259_init <= '0' ;
	p_reg_q259: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q259 <= reg_q259_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q259 <= reg_q259_init;
        else
          reg_q259 <= reg_q259_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q554_in <= (reg_q552 AND symb_decoder(16#5f#));
reg_q554_init <= '0' ;
	p_reg_q554: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q554 <= reg_q554_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q554 <= reg_q554_init;
        else
          reg_q554 <= reg_q554_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2495_in <= (reg_q2493 AND symb_decoder(16#32#));
reg_q2495_init <= '0' ;
	p_reg_q2495: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2495 <= reg_q2495_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2495 <= reg_q2495_init;
        else
          reg_q2495 <= reg_q2495_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2184_in <= (reg_q2182 AND symb_decoder(16#49#)) OR
 					(reg_q2182 AND symb_decoder(16#69#));
reg_q2184_init <= '0' ;
	p_reg_q2184: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2184 <= reg_q2184_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2184 <= reg_q2184_init;
        else
          reg_q2184 <= reg_q2184_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2068_in <= (reg_q2066 AND symb_decoder(16#46#));
reg_q2068_init <= '0' ;
	p_reg_q2068: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2068 <= reg_q2068_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2068 <= reg_q2068_init;
        else
          reg_q2068 <= reg_q2068_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q572_in <= (reg_q570 AND symb_decoder(16#31#));
reg_q572_init <= '0' ;
	p_reg_q572: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q572 <= reg_q572_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q572 <= reg_q572_init;
        else
          reg_q572 <= reg_q572_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2004_in <= (reg_q2002 AND symb_decoder(16#66#)) OR
 					(reg_q2002 AND symb_decoder(16#46#));
reg_q2004_init <= '0' ;
	p_reg_q2004: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2004 <= reg_q2004_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2004 <= reg_q2004_init;
        else
          reg_q2004 <= reg_q2004_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q30_in <= (reg_q28 AND symb_decoder(16#43#)) OR
 					(reg_q28 AND symb_decoder(16#63#));
reg_q30_init <= '0' ;
	p_reg_q30: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q30 <= reg_q30_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q30 <= reg_q30_init;
        else
          reg_q30 <= reg_q30_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2478_in <= (reg_q2476 AND symb_decoder(16#31#));
reg_q2478_init <= '0' ;
	p_reg_q2478: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2478 <= reg_q2478_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2478 <= reg_q2478_init;
        else
          reg_q2478 <= reg_q2478_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q482_in <= (reg_q480 AND symb_decoder(16#32#));
reg_q482_init <= '0' ;
	p_reg_q482: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q482 <= reg_q482_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q482 <= reg_q482_init;
        else
          reg_q482 <= reg_q482_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q484_in <= (reg_q482 AND symb_decoder(16#2e#));
reg_q484_init <= '0' ;
	p_reg_q484: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q484 <= reg_q484_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q484 <= reg_q484_init;
        else
          reg_q484 <= reg_q484_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q490_in <= (reg_q488 AND symb_decoder(16#32#));
reg_q490_init <= '0' ;
	p_reg_q490: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q490 <= reg_q490_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q490 <= reg_q490_init;
        else
          reg_q490 <= reg_q490_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2449_in <= (reg_q2447 AND symb_decoder(16#23#));
reg_q2449_init <= '0' ;
	p_reg_q2449: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2449 <= reg_q2449_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2449 <= reg_q2449_init;
        else
          reg_q2449 <= reg_q2449_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2547_in <= (reg_q2545 AND symb_decoder(16#65#)) OR
 					(reg_q2545 AND symb_decoder(16#45#));
reg_q2547_init <= '0' ;
	p_reg_q2547: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2547 <= reg_q2547_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2547 <= reg_q2547_init;
        else
          reg_q2547 <= reg_q2547_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q953_in <= (reg_q951 AND symb_decoder(16#00#));
reg_q953_init <= '0' ;
	p_reg_q953: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q953 <= reg_q953_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q953 <= reg_q953_init;
        else
          reg_q953 <= reg_q953_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2060_in <= (reg_q2058 AND symb_decoder(16#65#));
reg_q2060_init <= '0' ;
	p_reg_q2060: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2060 <= reg_q2060_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2060 <= reg_q2060_init;
        else
          reg_q2060 <= reg_q2060_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q783_in <= (reg_q781 AND symb_decoder(16#4d#)) OR
 					(reg_q781 AND symb_decoder(16#6d#));
reg_q783_init <= '0' ;
	p_reg_q783: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q783 <= reg_q783_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q783 <= reg_q783_init;
        else
          reg_q783 <= reg_q783_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q893_in <= (reg_q889 AND symb_decoder(16#5c#)) OR
 					(reg_q896 AND symb_decoder(16#5c#));
reg_q893_init <= '0' ;
	p_reg_q893: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q893 <= reg_q893_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q893 <= reg_q893_init;
        else
          reg_q893 <= reg_q893_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q886_in <= (reg_q893 AND symb_decoder(16#5d#));
reg_q886_init <= '0' ;
	p_reg_q886: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q886 <= reg_q886_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q886 <= reg_q886_init;
        else
          reg_q886 <= reg_q886_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2062_in <= (reg_q2060 AND symb_decoder(16#66#));
reg_q2062_init <= '0' ;
	p_reg_q2062: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2062 <= reg_q2062_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2062 <= reg_q2062_init;
        else
          reg_q2062 <= reg_q2062_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2381_in <= (reg_q2379 AND symb_decoder(16#0a#));
reg_q2381_init <= '0' ;
	p_reg_q2381: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2381 <= reg_q2381_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2381 <= reg_q2381_init;
        else
          reg_q2381 <= reg_q2381_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q648_in <= (reg_q646 AND symb_decoder(16#32#));
reg_q648_init <= '0' ;
	p_reg_q648: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q648 <= reg_q648_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q648 <= reg_q648_init;
        else
          reg_q648 <= reg_q648_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q811_in <= (reg_q809 AND symb_decoder(16#5e#));
reg_q811_init <= '0' ;
	p_reg_q811: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q811 <= reg_q811_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q811 <= reg_q811_init;
        else
          reg_q811 <= reg_q811_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1641_in <= (reg_q1639 AND symb_decoder(16#0a#));
reg_q1641_init <= '0' ;
	p_reg_q1641: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1641 <= reg_q1641_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1641 <= reg_q1641_init;
        else
          reg_q1641 <= reg_q1641_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q677_in <= (reg_q675 AND symb_decoder(16#5c#));
reg_q677_init <= '0' ;
	p_reg_q677: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q677 <= reg_q677_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q677 <= reg_q677_init;
        else
          reg_q677 <= reg_q677_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q662_in <= (reg_q660 AND symb_decoder(16#31#));
reg_q662_init <= '0' ;
	p_reg_q662: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q662 <= reg_q662_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q662 <= reg_q662_init;
        else
          reg_q662 <= reg_q662_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q846_in <= (reg_q844 AND symb_decoder(16#5e#));
reg_q846_init <= '0' ;
	p_reg_q846: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q846 <= reg_q846_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q846 <= reg_q846_init;
        else
          reg_q846 <= reg_q846_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2690_in <= (reg_q2688 AND symb_decoder(16#5c#));
reg_q2690_init <= '0' ;
	p_reg_q2690: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2690 <= reg_q2690_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2690 <= reg_q2690_init;
        else
          reg_q2690 <= reg_q2690_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2088_in <= (reg_q2086 AND symb_decoder(16#3a#));
reg_q2088_init <= '0' ;
	p_reg_q2088: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2088 <= reg_q2088_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2088 <= reg_q2088_init;
        else
          reg_q2088 <= reg_q2088_in;
        end if;
      end if;
    end if;
  end process;

	FINAL <= reg_q1541 OR reg_q2530 OR reg_q2320 OR reg_q1221 OR reg_q300 OR reg_q1600 OR reg_q1952 OR reg_q175 OR reg_q88 OR reg_q886 OR reg_q2121 OR reg_q811 OR reg_q1193 OR reg_q1010 OR reg_q2465 OR reg_q953 OR reg_q2206 OR reg_q2613 OR reg_q1882 OR reg_q2516 OR reg_q1824 OR reg_q2482 OR reg_q1108 OR reg_q554 OR reg_q2088 OR reg_q662 OR reg_q776 OR reg_q1995 OR reg_q1518 OR reg_q1449 OR reg_q700 OR reg_q1641 OR reg_q2692 OR reg_q1047 OR reg_q2693 OR reg_q411 OR reg_q259 OR reg_q677 OR reg_q1357 OR reg_q2381 OR reg_q887 OR reg_q44 OR reg_q2499 OR reg_q222 OR reg_q1294 OR reg_q711 OR reg_q2050 OR reg_q2249 OR reg_q884 OR reg_q846 OR reg_q1740 OR reg_q450;

	end architecture;
	