
	library ieee;
use ieee.std_logic_1164.all;

architecture http_backdoor of pattern_match is

--#################################################
-- start section fullgraph: 0

  -- state q2695
  signal reg_q2695        : std_logic;
  signal reg_q2695_in     : std_logic;
  		

  -- state q1452
  signal reg_q1452        : std_logic;
  signal reg_q1452_in     : std_logic;
  		
  signal reg_fullgraph0       : std_logic_vector(1 downto 0);
  signal reg_fullgraph0_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph0_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph0_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph0
  --#################################################			
		

  -- state q1826
  signal reg_q1826        : std_logic;
  signal reg_q1826_in     : std_logic;
  signal reg_q1826_init   : std_logic;
		
--#################################################
-- start section fullgraph: 2

  -- state q1139
  signal reg_q1139        : std_logic;
  signal reg_q1139_in     : std_logic;
  		

  -- state q828
  signal reg_q828        : std_logic;
  signal reg_q828_in     : std_logic;
  		

  -- state q848
  signal reg_q848        : std_logic;
  signal reg_q848_in     : std_logic;
  		

  -- state q2579
  signal reg_q2579        : std_logic;
  signal reg_q2579_in     : std_logic;
  		

  -- state q955
  signal reg_q955        : std_logic;
  signal reg_q955_in     : std_logic;
  		

  -- state q933
  signal reg_q933        : std_logic;
  signal reg_q933_in     : std_logic;
  		

  -- state q251
  signal reg_q251        : std_logic;
  signal reg_q251_in     : std_logic;
  		

  -- state q253
  signal reg_q253        : std_logic;
  signal reg_q253_in     : std_logic;
  		

  -- state q1331
  signal reg_q1331        : std_logic;
  signal reg_q1331_in     : std_logic;
  		

  -- state q1333
  signal reg_q1333        : std_logic;
  signal reg_q1333_in     : std_logic;
  		

  -- state q1997
  signal reg_q1997        : std_logic;
  signal reg_q1997_in     : std_logic;
  		

  -- state q2302
  signal reg_q2302        : std_logic;
  signal reg_q2302_in     : std_logic;
  		

  -- state q361
  signal reg_q361        : std_logic;
  signal reg_q361_in     : std_logic;
  		

  -- state q363
  signal reg_q363        : std_logic;
  signal reg_q363_in     : std_logic;
  		

  -- state q1104
  signal reg_q1104        : std_logic;
  signal reg_q1104_in     : std_logic;
  		

  -- state q1106
  signal reg_q1106        : std_logic;
  signal reg_q1106_in     : std_logic;
  		

  -- state q1668
  signal reg_q1668        : std_logic;
  signal reg_q1668_in     : std_logic;
  		

  -- state q1670
  signal reg_q1670        : std_logic;
  signal reg_q1670_in     : std_logic;
  		

  -- state q2351
  signal reg_q2351        : std_logic;
  signal reg_q2351_in     : std_logic;
  		

  -- state q420
  signal reg_q420        : std_logic;
  signal reg_q420_in     : std_logic;
  		

  -- state q422
  signal reg_q422        : std_logic;
  signal reg_q422_in     : std_logic;
  		

  -- state q1147
  signal reg_q1147        : std_logic;
  signal reg_q1147_in     : std_logic;
  		

  -- state q982
  signal reg_q982        : std_logic;
  signal reg_q982_in     : std_logic;
  		

  -- state q984
  signal reg_q984        : std_logic;
  signal reg_q984_in     : std_logic;
  		

  -- state q1299
  signal reg_q1299        : std_logic;
  signal reg_q1299_in     : std_logic;
  		

  -- state q2603
  signal reg_q2603        : std_logic;
  signal reg_q2603_in     : std_logic;
  		

  -- state q2605
  signal reg_q2605        : std_logic;
  signal reg_q2605_in     : std_logic;
  		

  -- state q2172
  signal reg_q2172        : std_logic;
  signal reg_q2172_in     : std_logic;
  		

  -- state q2274
  signal reg_q2274        : std_logic;
  signal reg_q2274_in     : std_logic;
  		

  -- state q2276
  signal reg_q2276        : std_logic;
  signal reg_q2276_in     : std_logic;
  		

  -- state q1035
  signal reg_q1035        : std_logic;
  signal reg_q1035_in     : std_logic;
  		

  -- state q1037
  signal reg_q1037        : std_logic;
  signal reg_q1037_in     : std_logic;
  		

  -- state q671
  signal reg_q671        : std_logic;
  signal reg_q671_in     : std_logic;
  		

  -- state q673
  signal reg_q673        : std_logic;
  signal reg_q673_in     : std_logic;
  		

  -- state q1478
  signal reg_q1478        : std_logic;
  signal reg_q1478_in     : std_logic;
  		

  -- state q1480
  signal reg_q1480        : std_logic;
  signal reg_q1480_in     : std_logic;
  		

  -- state q2018
  signal reg_q2018        : std_logic;
  signal reg_q2018_in     : std_logic;
  		

  -- state q2020
  signal reg_q2020        : std_logic;
  signal reg_q2020_in     : std_logic;
  		

  -- state q1527
  signal reg_q1527        : std_logic;
  signal reg_q1527_in     : std_logic;
  		

  -- state q1529
  signal reg_q1529        : std_logic;
  signal reg_q1529_in     : std_logic;
  		

  -- state q1301
  signal reg_q1301        : std_logic;
  signal reg_q1301_in     : std_logic;
  		

  -- state q1660
  signal reg_q1660        : std_logic;
  signal reg_q1660_in     : std_logic;
  		

  -- state q1662
  signal reg_q1662        : std_logic;
  signal reg_q1662_in     : std_logic;
  		

  -- state q1441
  signal reg_q1441        : std_logic;
  signal reg_q1441_in     : std_logic;
  		

  -- state q1443
  signal reg_q1443        : std_logic;
  signal reg_q1443_in     : std_logic;
  		

  -- state q2353
  signal reg_q2353        : std_logic;
  signal reg_q2353_in     : std_logic;
  		

  -- state q2278
  signal reg_q2278        : std_logic;
  signal reg_q2278_in     : std_logic;
  		

  -- state q1027
  signal reg_q1027        : std_logic;
  signal reg_q1027_in     : std_logic;
  		

  -- state q1029
  signal reg_q1029        : std_logic;
  signal reg_q1029_in     : std_logic;
  		

  -- state q1084
  signal reg_q1084        : std_logic;
  signal reg_q1084_in     : std_logic;
  		

  -- state q1086
  signal reg_q1086        : std_logic;
  signal reg_q1086_in     : std_logic;
  		

  -- state q2514
  signal reg_q2514        : std_logic;
  signal reg_q2514_in     : std_logic;
  		

  -- state q2516
  signal reg_q2516        : std_logic;
  signal reg_q2516_in     : std_logic;
  		

  -- state q1724
  signal reg_q1724        : std_logic;
  signal reg_q1724_in     : std_logic;
  		

  -- state q1726
  signal reg_q1726        : std_logic;
  signal reg_q1726_in     : std_logic;
  		

  -- state q1335
  signal reg_q1335        : std_logic;
  signal reg_q1335_in     : std_logic;
  		

  -- state q2109
  signal reg_q2109        : std_logic;
  signal reg_q2109_in     : std_logic;
  		

  -- state q2111
  signal reg_q2111        : std_logic;
  signal reg_q2111_in     : std_logic;
  		

  -- state q1355
  signal reg_q1355        : std_logic;
  signal reg_q1355_in     : std_logic;
  		

  -- state q1357
  signal reg_q1357        : std_logic;
  signal reg_q1357_in     : std_logic;
  		

  -- state q2004
  signal reg_q2004        : std_logic;
  signal reg_q2004_in     : std_logic;
  		

  -- state q1191
  signal reg_q1191        : std_logic;
  signal reg_q1191_in     : std_logic;
  		

  -- state q1193
  signal reg_q1193        : std_logic;
  signal reg_q1193_in     : std_logic;
  		

  -- state q1580
  signal reg_q1580        : std_logic;
  signal reg_q1580_in     : std_logic;
  		

  -- state q824
  signal reg_q824        : std_logic;
  signal reg_q824_in     : std_logic;
  		

  -- state q826
  signal reg_q826        : std_logic;
  signal reg_q826_in     : std_logic;
  		

  -- state q690
  signal reg_q690        : std_logic;
  signal reg_q690_in     : std_logic;
  		

  -- state q692
  signal reg_q692        : std_logic;
  signal reg_q692_in     : std_logic;
  		

  -- state q709
  signal reg_q709        : std_logic;
  signal reg_q709_in     : std_logic;
  		

  -- state q711
  signal reg_q711        : std_logic;
  signal reg_q711_in     : std_logic;
  		

  -- state q373
  signal reg_q373        : std_logic;
  signal reg_q373_in     : std_logic;
  		

  -- state q375
  signal reg_q375        : std_logic;
  signal reg_q375_in     : std_logic;
  		

  -- state q247
  signal reg_q247        : std_logic;
  signal reg_q247_in     : std_logic;
  		

  -- state q249
  signal reg_q249        : std_logic;
  signal reg_q249_in     : std_logic;
  		

  -- state q2038
  signal reg_q2038        : std_logic;
  signal reg_q2038_in     : std_logic;
  		

  -- state q2040
  signal reg_q2040        : std_logic;
  signal reg_q2040_in     : std_logic;
  		

  -- state q1975
  signal reg_q1975        : std_logic;
  signal reg_q1975_in     : std_logic;
  		

  -- state q1248
  signal reg_q1248        : std_logic;
  signal reg_q1248_in     : std_logic;
  		

  -- state q2369
  signal reg_q2369        : std_logic;
  signal reg_q2369_in     : std_logic;
  		

  -- state q1094
  signal reg_q1094        : std_logic;
  signal reg_q1094_in     : std_logic;
  		

  -- state q1096
  signal reg_q1096        : std_logic;
  signal reg_q1096_in     : std_logic;
  		

  -- state q1108
  signal reg_q1108        : std_logic;
  signal reg_q1108_in     : std_logic;
  		

  -- state q56
  signal reg_q56        : std_logic;
  signal reg_q56_in     : std_logic;
  		

  -- state q58
  signal reg_q58        : std_logic;
  signal reg_q58_in     : std_logic;
  		

  -- state q101
  signal reg_q101        : std_logic;
  signal reg_q101_in     : std_logic;
  		

  -- state q103
  signal reg_q103        : std_logic;
  signal reg_q103_in     : std_logic;
  		

  -- state q2480
  signal reg_q2480        : std_logic;
  signal reg_q2480_in     : std_logic;
  		

  -- state q2482
  signal reg_q2482        : std_logic;
  signal reg_q2482_in     : std_logic;
  		

  -- state q1482
  signal reg_q1482        : std_logic;
  signal reg_q1482_in     : std_logic;
  		

  -- state q367
  signal reg_q367        : std_logic;
  signal reg_q367_in     : std_logic;
  		

  -- state q369
  signal reg_q369        : std_logic;
  signal reg_q369_in     : std_logic;
  		

  -- state q700
  signal reg_q700        : std_logic;
  signal reg_q700_in     : std_logic;
  		

  -- state q196
  signal reg_q196        : std_logic;
  signal reg_q196_in     : std_logic;
  		

  -- state q198
  signal reg_q198        : std_logic;
  signal reg_q198_in     : std_logic;
  		

  -- state q418
  signal reg_q418        : std_logic;
  signal reg_q418_in     : std_logic;
  		

  -- state q1688
  signal reg_q1688        : std_logic;
  signal reg_q1688_in     : std_logic;
  		

  -- state q1690
  signal reg_q1690        : std_logic;
  signal reg_q1690_in     : std_logic;
  		

  -- state q357
  signal reg_q357        : std_logic;
  signal reg_q357_in     : std_logic;
  		

  -- state q359
  signal reg_q359        : std_logic;
  signal reg_q359_in     : std_logic;
  		

  -- state q2101
  signal reg_q2101        : std_logic;
  signal reg_q2101_in     : std_logic;
  		

  -- state q2103
  signal reg_q2103        : std_logic;
  signal reg_q2103_in     : std_logic;
  		

  -- state q2375
  signal reg_q2375        : std_logic;
  signal reg_q2375_in     : std_logic;
  		

  -- state q2377
  signal reg_q2377        : std_logic;
  signal reg_q2377_in     : std_logic;
  		

  -- state q2361
  signal reg_q2361        : std_logic;
  signal reg_q2361_in     : std_logic;
  		

  -- state q2363
  signal reg_q2363        : std_logic;
  signal reg_q2363_in     : std_logic;
  		

  -- state q121
  signal reg_q121        : std_logic;
  signal reg_q121_in     : std_logic;
  		

  -- state q123
  signal reg_q123        : std_logic;
  signal reg_q123_in     : std_logic;
  		

  -- state q2613
  signal reg_q2613        : std_logic;
  signal reg_q2613_in     : std_logic;
  		

  -- state q818
  signal reg_q818        : std_logic;
  signal reg_q818_in     : std_logic;
  		

  -- state q2593
  signal reg_q2593        : std_logic;
  signal reg_q2593_in     : std_logic;
  		

  -- state q2595
  signal reg_q2595        : std_logic;
  signal reg_q2595_in     : std_logic;
  		

  -- state q426
  signal reg_q426        : std_logic;
  signal reg_q426_in     : std_logic;
  		

  -- state q428
  signal reg_q428        : std_logic;
  signal reg_q428_in     : std_logic;
  		

  -- state q2337
  signal reg_q2337        : std_logic;
  signal reg_q2337_in     : std_logic;
  		

  -- state q127
  signal reg_q127        : std_logic;
  signal reg_q127_in     : std_logic;
  		

  -- state q1337
  signal reg_q1337        : std_logic;
  signal reg_q1337_in     : std_logic;
  		

  -- state q2341
  signal reg_q2341        : std_logic;
  signal reg_q2341_in     : std_logic;
  		

  -- state q2343
  signal reg_q2343        : std_logic;
  signal reg_q2343_in     : std_logic;
  		

  -- state q966
  signal reg_q966        : std_logic;
  signal reg_q966_in     : std_logic;
  		

  -- state q968
  signal reg_q968        : std_logic;
  signal reg_q968_in     : std_logic;
  		

  -- state q1676
  signal reg_q1676        : std_logic;
  signal reg_q1676_in     : std_logic;
  		

  -- state q1678
  signal reg_q1678        : std_logic;
  signal reg_q1678_in     : std_logic;
  		

  -- state q379
  signal reg_q379        : std_logic;
  signal reg_q379_in     : std_logic;
  		

  -- state q381
  signal reg_q381        : std_logic;
  signal reg_q381_in     : std_logic;
  		

  -- state q2577
  signal reg_q2577        : std_logic;
  signal reg_q2577_in     : std_logic;
  		

  -- state q2688
  signal reg_q2688        : std_logic;
  signal reg_q2688_in     : std_logic;
  		

  -- state q2690
  signal reg_q2690        : std_logic;
  signal reg_q2690_in     : std_logic;
  		

  -- state q1531
  signal reg_q1531        : std_logic;
  signal reg_q1531_in     : std_logic;
  		

  -- state q1674
  signal reg_q1674        : std_logic;
  signal reg_q1674_in     : std_logic;
  		

  -- state q756
  signal reg_q756        : std_logic;
  signal reg_q756_in     : std_logic;
  		

  -- state q1305
  signal reg_q1305        : std_logic;
  signal reg_q1305_in     : std_logic;
  		

  -- state q1307
  signal reg_q1307        : std_logic;
  signal reg_q1307_in     : std_logic;
  		

  -- state q1425
  signal reg_q1425        : std_logic;
  signal reg_q1425_in     : std_logic;
  		

  -- state q1427
  signal reg_q1427        : std_logic;
  signal reg_q1427_in     : std_logic;
  		

  -- state q194
  signal reg_q194        : std_logic;
  signal reg_q194_in     : std_logic;
  		

  -- state q115
  signal reg_q115        : std_logic;
  signal reg_q115_in     : std_logic;
  		

  -- state q117
  signal reg_q117        : std_logic;
  signal reg_q117_in     : std_logic;
  		

  -- state q1250
  signal reg_q1250        : std_logic;
  signal reg_q1250_in     : std_logic;
  		

  -- state q1252
  signal reg_q1252        : std_logic;
  signal reg_q1252_in     : std_logic;
  		

  -- state q2620
  signal reg_q2620        : std_logic;
  signal reg_q2620_in     : std_logic;
  		

  -- state q2622
  signal reg_q2622        : std_logic;
  signal reg_q2622_in     : std_logic;
  		

  -- state q2042
  signal reg_q2042        : std_logic;
  signal reg_q2042_in     : std_logic;
  		

  -- state q1421
  signal reg_q1421        : std_logic;
  signal reg_q1421_in     : std_logic;
  		

  -- state q1423
  signal reg_q1423        : std_logic;
  signal reg_q1423_in     : std_logic;
  		

  -- state q1680
  signal reg_q1680        : std_logic;
  signal reg_q1680_in     : std_logic;
  		

  -- state q1682
  signal reg_q1682        : std_logic;
  signal reg_q1682_in     : std_logic;
  		

  -- state q74
  signal reg_q74        : std_logic;
  signal reg_q74_in     : std_logic;
  		

  -- state q76
  signal reg_q76        : std_logic;
  signal reg_q76_in     : std_logic;
  		

  -- state q113
  signal reg_q113        : std_logic;
  signal reg_q113_in     : std_logic;
  		

  -- state q1187
  signal reg_q1187        : std_logic;
  signal reg_q1187_in     : std_logic;
  		

  -- state q1189
  signal reg_q1189        : std_logic;
  signal reg_q1189_in     : std_logic;
  		

  -- state q1714
  signal reg_q1714        : std_logic;
  signal reg_q1714_in     : std_logic;
  		

  -- state q1716
  signal reg_q1716        : std_logic;
  signal reg_q1716_in     : std_logic;
  		

  -- state q341
  signal reg_q341        : std_logic;
  signal reg_q341_in     : std_logic;
  		

  -- state q343
  signal reg_q343        : std_logic;
  signal reg_q343_in     : std_logic;
  		

  -- state q2117
  signal reg_q2117        : std_logic;
  signal reg_q2117_in     : std_logic;
  		

  -- state q2119
  signal reg_q2119        : std_logic;
  signal reg_q2119_in     : std_logic;
  		

  -- state q1574
  signal reg_q1574        : std_logic;
  signal reg_q1574_in     : std_logic;
  		

  -- state q1576
  signal reg_q1576        : std_logic;
  signal reg_q1576_in     : std_logic;
  		

  -- state q2215
  signal reg_q2215        : std_logic;
  signal reg_q2215_in     : std_logic;
  		

  -- state q2217
  signal reg_q2217        : std_logic;
  signal reg_q2217_in     : std_logic;
  		

  -- state q2609
  signal reg_q2609        : std_logic;
  signal reg_q2609_in     : std_logic;
  		

  -- state q2611
  signal reg_q2611        : std_logic;
  signal reg_q2611_in     : std_logic;
  		

  -- state q2168
  signal reg_q2168        : std_logic;
  signal reg_q2168_in     : std_logic;
  		

  -- state q2170
  signal reg_q2170        : std_logic;
  signal reg_q2170_in     : std_logic;
  		

  -- state q994
  signal reg_q994        : std_logic;
  signal reg_q994_in     : std_logic;
  		

  -- state q996
  signal reg_q996        : std_logic;
  signal reg_q996_in     : std_logic;
  		

  -- state q237
  signal reg_q237        : std_logic;
  signal reg_q237_in     : std_logic;
  		

  -- state q257
  signal reg_q257        : std_logic;
  signal reg_q257_in     : std_logic;
  		

  -- state q2535
  signal reg_q2535        : std_logic;
  signal reg_q2535_in     : std_logic;
  		

  -- state q2537
  signal reg_q2537        : std_logic;
  signal reg_q2537_in     : std_logic;
  		

  -- state q2284
  signal reg_q2284        : std_logic;
  signal reg_q2284_in     : std_logic;
  		

  -- state q2286
  signal reg_q2286        : std_logic;
  signal reg_q2286_in     : std_logic;
  		

  -- state q682
  signal reg_q682        : std_logic;
  signal reg_q682_in     : std_logic;
  		

  -- state q998
  signal reg_q998        : std_logic;
  signal reg_q998_in     : std_logic;
  		

  -- state q1000
  signal reg_q1000        : std_logic;
  signal reg_q1000_in     : std_logic;
  		

  -- state q1698
  signal reg_q1698        : std_logic;
  signal reg_q1698_in     : std_logic;
  		

  -- state q1700
  signal reg_q1700        : std_logic;
  signal reg_q1700_in     : std_logic;
  		

  -- state q2243
  signal reg_q2243        : std_logic;
  signal reg_q2243_in     : std_logic;
  		

  -- state q2245
  signal reg_q2245        : std_logic;
  signal reg_q2245_in     : std_logic;
  		

  -- state q1578
  signal reg_q1578        : std_logic;
  signal reg_q1578_in     : std_logic;
  		

  -- state q1145
  signal reg_q1145        : std_logic;
  signal reg_q1145_in     : std_logic;
  		

  -- state q1736
  signal reg_q1736        : std_logic;
  signal reg_q1736_in     : std_logic;
  		

  -- state q1738
  signal reg_q1738        : std_logic;
  signal reg_q1738_in     : std_logic;
  		

  -- state q2670
  signal reg_q2670        : std_logic;
  signal reg_q2670_in     : std_logic;
  		

  -- state q2672
  signal reg_q2672        : std_logic;
  signal reg_q2672_in     : std_logic;
  		

  -- state q288
  signal reg_q288        : std_logic;
  signal reg_q288_in     : std_logic;
  		

  -- state q290
  signal reg_q290        : std_logic;
  signal reg_q290_in     : std_logic;
  		

  -- state q125
  signal reg_q125        : std_logic;
  signal reg_q125_in     : std_logic;
  		

  -- state q1002
  signal reg_q1002        : std_logic;
  signal reg_q1002_in     : std_logic;
  		

  -- state q980
  signal reg_q980        : std_logic;
  signal reg_q980_in     : std_logic;
  		

  -- state q1702
  signal reg_q1702        : std_logic;
  signal reg_q1702_in     : std_logic;
  		

  -- state q371
  signal reg_q371        : std_logic;
  signal reg_q371_in     : std_logic;
  		

  -- state q919
  signal reg_q919        : std_logic;
  signal reg_q919_in     : std_logic;
  		

  -- state q921
  signal reg_q921        : std_logic;
  signal reg_q921_in     : std_logic;
  		

  -- state q1582
  signal reg_q1582        : std_logic;
  signal reg_q1582_in     : std_logic;
  		

  -- state q931
  signal reg_q931        : std_logic;
  signal reg_q931_in     : std_logic;
  		

  -- state q1315
  signal reg_q1315        : std_logic;
  signal reg_q1315_in     : std_logic;
  		

  -- state q1317
  signal reg_q1317        : std_logic;
  signal reg_q1317_in     : std_logic;
  		

  -- state q1102
  signal reg_q1102        : std_logic;
  signal reg_q1102_in     : std_logic;
  		

  -- state q2692
  signal reg_q2692        : std_logic;
  signal reg_q2692_in     : std_logic;
  		

  -- state q2371
  signal reg_q2371        : std_logic;
  signal reg_q2371_in     : std_logic;
  		

  -- state q2373
  signal reg_q2373        : std_logic;
  signal reg_q2373_in     : std_logic;
  		

  -- state q2589
  signal reg_q2589        : std_logic;
  signal reg_q2589_in     : std_logic;
  		

  -- state q2591
  signal reg_q2591        : std_logic;
  signal reg_q2591_in     : std_logic;
  		

  -- state q2030
  signal reg_q2030        : std_logic;
  signal reg_q2030_in     : std_logic;
  		

  -- state q1339
  signal reg_q1339        : std_logic;
  signal reg_q1339_in     : std_logic;
  		

  -- state q1341
  signal reg_q1341        : std_logic;
  signal reg_q1341_in     : std_logic;
  		

  -- state q167
  signal reg_q167        : std_logic;
  signal reg_q167_in     : std_logic;
  		

  -- state q169
  signal reg_q169        : std_logic;
  signal reg_q169_in     : std_logic;
  		

  -- state q450
  signal reg_q450        : std_logic;
  signal reg_q450_in     : std_logic;
  		

  -- state q2221
  signal reg_q2221        : std_logic;
  signal reg_q2221_in     : std_logic;
  		

  -- state q2223
  signal reg_q2223        : std_logic;
  signal reg_q2223_in     : std_logic;
  		

  -- state q2634
  signal reg_q2634        : std_logic;
  signal reg_q2634_in     : std_logic;
  		

  -- state q2636
  signal reg_q2636        : std_logic;
  signal reg_q2636_in     : std_logic;
  		

  -- state q2272
  signal reg_q2272        : std_logic;
  signal reg_q2272_in     : std_logic;
  		

  -- state q2115
  signal reg_q2115        : std_logic;
  signal reg_q2115_in     : std_logic;
  		

  -- state q333
  signal reg_q333        : std_logic;
  signal reg_q333_in     : std_logic;
  		

  -- state q335
  signal reg_q335        : std_logic;
  signal reg_q335_in     : std_logic;
  		

  -- state q1460
  signal reg_q1460        : std_logic;
  signal reg_q1460_in     : std_logic;
  		

  -- state q1462
  signal reg_q1462        : std_logic;
  signal reg_q1462_in     : std_logic;
  		

  -- state q2333
  signal reg_q2333        : std_logic;
  signal reg_q2333_in     : std_logic;
  		

  -- state q2335
  signal reg_q2335        : std_logic;
  signal reg_q2335_in     : std_logic;
  		

  -- state q2227
  signal reg_q2227        : std_logic;
  signal reg_q2227_in     : std_logic;
  		

  -- state q2229
  signal reg_q2229        : std_logic;
  signal reg_q2229_in     : std_logic;
  		

  -- state q1466
  signal reg_q1466        : std_logic;
  signal reg_q1466_in     : std_logic;
  		

  -- state q1468
  signal reg_q1468        : std_logic;
  signal reg_q1468_in     : std_logic;
  		

  -- state q1072
  signal reg_q1072        : std_logic;
  signal reg_q1072_in     : std_logic;
  		

  -- state q1074
  signal reg_q1074        : std_logic;
  signal reg_q1074_in     : std_logic;
  		

  -- state q2474
  signal reg_q2474        : std_logic;
  signal reg_q2474_in     : std_logic;
  		

  -- state q2476
  signal reg_q2476        : std_logic;
  signal reg_q2476_in     : std_logic;
  		

  -- state q1560
  signal reg_q1560        : std_logic;
  signal reg_q1560_in     : std_logic;
  		

  -- state q1562
  signal reg_q1562        : std_logic;
  signal reg_q1562_in     : std_logic;
  		

  -- state q686
  signal reg_q686        : std_logic;
  signal reg_q686_in     : std_logic;
  		

  -- state q688
  signal reg_q688        : std_logic;
  signal reg_q688_in     : std_logic;
  		

  -- state q1734
  signal reg_q1734        : std_logic;
  signal reg_q1734_in     : std_logic;
  		

  -- state q1704
  signal reg_q1704        : std_logic;
  signal reg_q1704_in     : std_logic;
  		

  -- state q305
  signal reg_q305        : std_logic;
  signal reg_q305_in     : std_logic;
  		

  -- state q2028
  signal reg_q2028        : std_logic;
  signal reg_q2028_in     : std_logic;
  		

  -- state q235
  signal reg_q235        : std_logic;
  signal reg_q235_in     : std_logic;
  		

  -- state q1143
  signal reg_q1143        : std_logic;
  signal reg_q1143_in     : std_logic;
  		

  -- state q1541
  signal reg_q1541        : std_logic;
  signal reg_q1541_in     : std_logic;
  		

  -- state q1546
  signal reg_q1546        : std_logic;
  signal reg_q1546_in     : std_logic;
  		

  -- state q1548
  signal reg_q1548        : std_logic;
  signal reg_q1548_in     : std_logic;
  		

  -- state q2022
  signal reg_q2022        : std_logic;
  signal reg_q2022_in     : std_logic;
  		

  -- state q2024
  signal reg_q2024        : std_logic;
  signal reg_q2024_in     : std_logic;
  		

  -- state q1730
  signal reg_q1730        : std_logic;
  signal reg_q1730_in     : std_logic;
  		

  -- state q1732
  signal reg_q1732        : std_logic;
  signal reg_q1732_in     : std_logic;
  		

  -- state q2225
  signal reg_q2225        : std_logic;
  signal reg_q2225_in     : std_logic;
  		

  -- state q1470
  signal reg_q1470        : std_logic;
  signal reg_q1470_in     : std_logic;
  		

  -- state q1472
  signal reg_q1472        : std_logic;
  signal reg_q1472_in     : std_logic;
  		

  -- state q111
  signal reg_q111        : std_logic;
  signal reg_q111_in     : std_logic;
  		

  -- state q133
  signal reg_q133        : std_logic;
  signal reg_q133_in     : std_logic;
  		

  -- state q135
  signal reg_q135        : std_logic;
  signal reg_q135_in     : std_logic;
  		

  -- state q2292
  signal reg_q2292        : std_logic;
  signal reg_q2292_in     : std_logic;
  		

  -- state q2294
  signal reg_q2294        : std_logic;
  signal reg_q2294_in     : std_logic;
  		

  -- state q1080
  signal reg_q1080        : std_logic;
  signal reg_q1080_in     : std_logic;
  		

  -- state q1082
  signal reg_q1082        : std_logic;
  signal reg_q1082_in     : std_logic;
  		

  -- state q2247
  signal reg_q2247        : std_logic;
  signal reg_q2247_in     : std_logic;
  		

  -- state q2249
  signal reg_q2249        : std_logic;
  signal reg_q2249_in     : std_logic;
  		

  -- state q245
  signal reg_q245        : std_logic;
  signal reg_q245_in     : std_logic;
  		

  -- state q742
  signal reg_q742        : std_logic;
  signal reg_q742_in     : std_logic;
  		

  -- state q744
  signal reg_q744        : std_logic;
  signal reg_q744_in     : std_logic;
  		

  -- state q1090
  signal reg_q1090        : std_logic;
  signal reg_q1090_in     : std_logic;
  		

  -- state q129
  signal reg_q129        : std_logic;
  signal reg_q129_in     : std_logic;
  		

  -- state q1135
  signal reg_q1135        : std_logic;
  signal reg_q1135_in     : std_logic;
  		

  -- state q1137
  signal reg_q1137        : std_logic;
  signal reg_q1137_in     : std_logic;
  		

  -- state q1431
  signal reg_q1431        : std_logic;
  signal reg_q1431_in     : std_logic;
  		

  -- state q1433
  signal reg_q1433        : std_logic;
  signal reg_q1433_in     : std_logic;
  		

  -- state q2308
  signal reg_q2308        : std_logic;
  signal reg_q2308_in     : std_logic;
  		

  -- state q2310
  signal reg_q2310        : std_logic;
  signal reg_q2310_in     : std_logic;
  		

  -- state q2597
  signal reg_q2597        : std_logic;
  signal reg_q2597_in     : std_logic;
  		

  -- state q1708
  signal reg_q1708        : std_logic;
  signal reg_q1708_in     : std_logic;
  		

  -- state q2258
  signal reg_q2258        : std_logic;
  signal reg_q2258_in     : std_logic;
  		

  -- state q2260
  signal reg_q2260        : std_logic;
  signal reg_q2260_in     : std_logic;
  		

  -- state q978
  signal reg_q978        : std_logic;
  signal reg_q978_in     : std_logic;
  		

  -- state q988
  signal reg_q988        : std_logic;
  signal reg_q988_in     : std_logic;
  		

  -- state q990
  signal reg_q990        : std_logic;
  signal reg_q990_in     : std_logic;
  		

  -- state q2565
  signal reg_q2565        : std_logic;
  signal reg_q2565_in     : std_logic;
  		

  -- state q2567
  signal reg_q2567        : std_logic;
  signal reg_q2567_in     : std_logic;
  		

  -- state q1325
  signal reg_q1325        : std_logic;
  signal reg_q1325_in     : std_logic;
  		

  -- state q1327
  signal reg_q1327        : std_logic;
  signal reg_q1327_in     : std_logic;
  		

  -- state q149
  signal reg_q149        : std_logic;
  signal reg_q149_in     : std_logic;
  		

  -- state q1088
  signal reg_q1088        : std_logic;
  signal reg_q1088_in     : std_logic;
  		

  -- state q137
  signal reg_q137        : std_logic;
  signal reg_q137_in     : std_logic;
  		

  -- state q675
  signal reg_q675        : std_logic;
  signal reg_q675_in     : std_logic;
  		

  -- state q2136
  signal reg_q2136        : std_logic;
  signal reg_q2136_in     : std_logic;
  		

  -- state q2138
  signal reg_q2138        : std_logic;
  signal reg_q2138_in     : std_logic;
  		

  -- state q119
  signal reg_q119        : std_logic;
  signal reg_q119_in     : std_logic;
  		

  -- state q255
  signal reg_q255        : std_logic;
  signal reg_q255_in     : std_logic;
  		

  -- state q915
  signal reg_q915        : std_logic;
  signal reg_q915_in     : std_logic;
  		

  -- state q1008
  signal reg_q1008        : std_logic;
  signal reg_q1008_in     : std_logic;
  		

  -- state q1010
  signal reg_q1010        : std_logic;
  signal reg_q1010_in     : std_logic;
  		

  -- state q1672
  signal reg_q1672        : std_logic;
  signal reg_q1672_in     : std_logic;
  		

  -- state q2642
  signal reg_q2642        : std_logic;
  signal reg_q2642_in     : std_logic;
  		

  -- state q2644
  signal reg_q2644        : std_logic;
  signal reg_q2644_in     : std_logic;
  		

  -- state q2599
  signal reg_q2599        : std_logic;
  signal reg_q2599_in     : std_logic;
  		

  -- state q2601
  signal reg_q2601        : std_logic;
  signal reg_q2601_in     : std_logic;
  		

  -- state q1637
  signal reg_q1637        : std_logic;
  signal reg_q1637_in     : std_logic;
  		

  -- state q1639
  signal reg_q1639        : std_logic;
  signal reg_q1639_in     : std_logic;
  		

  -- state q107
  signal reg_q107        : std_logic;
  signal reg_q107_in     : std_logic;
  		

  -- state q109
  signal reg_q109        : std_logic;
  signal reg_q109_in     : std_logic;
  		

  -- state q783
  signal reg_q783        : std_logic;
  signal reg_q783_in     : std_logic;
  		

  -- state q785
  signal reg_q785        : std_logic;
  signal reg_q785_in     : std_logic;
  		

  -- state q1092
  signal reg_q1092        : std_logic;
  signal reg_q1092_in     : std_logic;
  		

  -- state q1347
  signal reg_q1347        : std_logic;
  signal reg_q1347_in     : std_logic;
  		

  -- state q1349
  signal reg_q1349        : std_logic;
  signal reg_q1349_in     : std_logic;
  		

  -- state q1115
  signal reg_q1115        : std_logic;
  signal reg_q1115_in     : std_logic;
  		

  -- state q1117
  signal reg_q1117        : std_logic;
  signal reg_q1117_in     : std_logic;
  		

  -- state q448
  signal reg_q448        : std_logic;
  signal reg_q448_in     : std_logic;
  		

  -- state q192
  signal reg_q192        : std_logic;
  signal reg_q192_in     : std_logic;
  		

  -- state q395
  signal reg_q395        : std_logic;
  signal reg_q395_in     : std_logic;
  		

  -- state q397
  signal reg_q397        : std_logic;
  signal reg_q397_in     : std_logic;
  		

  -- state q84
  signal reg_q84        : std_logic;
  signal reg_q84_in     : std_logic;
  		

  -- state q86
  signal reg_q86        : std_logic;
  signal reg_q86_in     : std_logic;
  		

  -- state q365
  signal reg_q365        : std_logic;
  signal reg_q365_in     : std_logic;
  		

  -- state q698
  signal reg_q698        : std_logic;
  signal reg_q698_in     : std_logic;
  		

  -- state q1437
  signal reg_q1437        : std_logic;
  signal reg_q1437_in     : std_logic;
  		

  -- state q964
  signal reg_q964        : std_logic;
  signal reg_q964_in     : std_logic;
  		

  -- state q748
  signal reg_q748        : std_logic;
  signal reg_q748_in     : std_logic;
  		

  -- state q750
  signal reg_q750        : std_logic;
  signal reg_q750_in     : std_logic;
  		

  -- state q1435
  signal reg_q1435        : std_logic;
  signal reg_q1435_in     : std_logic;
  		

  -- state q1692
  signal reg_q1692        : std_logic;
  signal reg_q1692_in     : std_logic;
  		

  -- state q1262
  signal reg_q1262        : std_logic;
  signal reg_q1262_in     : std_logic;
  		

  -- state q1264
  signal reg_q1264        : std_logic;
  signal reg_q1264_in     : std_logic;
  		

  -- state q2686
  signal reg_q2686        : std_logic;
  signal reg_q2686_in     : std_logic;
  		

  -- state q2349
  signal reg_q2349        : std_logic;
  signal reg_q2349_in     : std_logic;
  		

  -- state q1023
  signal reg_q1023        : std_logic;
  signal reg_q1023_in     : std_logic;
  		

  -- state q1025
  signal reg_q1025        : std_logic;
  signal reg_q1025_in     : std_logic;
  		

  -- state q1133
  signal reg_q1133        : std_logic;
  signal reg_q1133_in     : std_logic;
  		

  -- state q2575
  signal reg_q2575        : std_logic;
  signal reg_q2575_in     : std_logic;
  		

  -- state q1272
  signal reg_q1272        : std_logic;
  signal reg_q1272_in     : std_logic;
  		

  -- state q1274
  signal reg_q1274        : std_logic;
  signal reg_q1274_in     : std_logic;
  		

  -- state q1504
  signal reg_q1504        : std_logic;
  signal reg_q1504_in     : std_logic;
  		

  -- state q1506
  signal reg_q1506        : std_logic;
  signal reg_q1506_in     : std_logic;
  		

  -- state q2497
  signal reg_q2497        : std_logic;
  signal reg_q2497_in     : std_logic;
  		

  -- state q2499
  signal reg_q2499        : std_logic;
  signal reg_q2499_in     : std_logic;
  		

  -- state q923
  signal reg_q923        : std_logic;
  signal reg_q923_in     : std_logic;
  		

  -- state q925
  signal reg_q925        : std_logic;
  signal reg_q925_in     : std_logic;
  		

  -- state q1635
  signal reg_q1635        : std_logic;
  signal reg_q1635_in     : std_logic;
  		

  -- state q323
  signal reg_q323        : std_logic;
  signal reg_q323_in     : std_logic;
  		

  -- state q325
  signal reg_q325        : std_logic;
  signal reg_q325_in     : std_logic;
  		

  -- state q292
  signal reg_q292        : std_logic;
  signal reg_q292_in     : std_logic;
  		

  -- state q294
  signal reg_q294        : std_logic;
  signal reg_q294_in     : std_logic;
  		

  -- state q1664
  signal reg_q1664        : std_logic;
  signal reg_q1664_in     : std_logic;
  		

  -- state q1666
  signal reg_q1666        : std_logic;
  signal reg_q1666_in     : std_logic;
  		

  -- state q377
  signal reg_q377        : std_logic;
  signal reg_q377_in     : std_logic;
  		

  -- state q1652
  signal reg_q1652        : std_logic;
  signal reg_q1652_in     : std_logic;
  		

  -- state q1728
  signal reg_q1728        : std_logic;
  signal reg_q1728_in     : std_logic;
  		

  -- state q1151
  signal reg_q1151        : std_logic;
  signal reg_q1151_in     : std_logic;
  		

  -- state q1153
  signal reg_q1153        : std_logic;
  signal reg_q1153_in     : std_logic;
  		

  -- state q1971
  signal reg_q1971        : std_logic;
  signal reg_q1971_in     : std_logic;
  		

  -- state q1973
  signal reg_q1973        : std_logic;
  signal reg_q1973_in     : std_logic;
  		

  -- state q1552
  signal reg_q1552        : std_logic;
  signal reg_q1552_in     : std_logic;
  		

  -- state q1179
  signal reg_q1179        : std_logic;
  signal reg_q1179_in     : std_logic;
  		

  -- state q1181
  signal reg_q1181        : std_logic;
  signal reg_q1181_in     : std_logic;
  		

  -- state q913
  signal reg_q913        : std_logic;
  signal reg_q913_in     : std_logic;
  		

  -- state q2304
  signal reg_q2304        : std_logic;
  signal reg_q2304_in     : std_logic;
  		

  -- state q2306
  signal reg_q2306        : std_logic;
  signal reg_q2306_in     : std_logic;
  		

  -- state q1319
  signal reg_q1319        : std_logic;
  signal reg_q1319_in     : std_logic;
  		

  -- state q986
  signal reg_q986        : std_logic;
  signal reg_q986_in     : std_logic;
  		

  -- state q82
  signal reg_q82        : std_logic;
  signal reg_q82_in     : std_logic;
  		

  -- state q280
  signal reg_q280        : std_logic;
  signal reg_q280_in     : std_logic;
  		

  -- state q282
  signal reg_q282        : std_logic;
  signal reg_q282_in     : std_logic;
  		

  -- state q2158
  signal reg_q2158        : std_logic;
  signal reg_q2158_in     : std_logic;
  		

  -- state q2160
  signal reg_q2160        : std_logic;
  signal reg_q2160_in     : std_logic;
  		

  -- state q1484
  signal reg_q1484        : std_logic;
  signal reg_q1484_in     : std_logic;
  		

  -- state q2674
  signal reg_q2674        : std_logic;
  signal reg_q2674_in     : std_logic;
  		

  -- state q2676
  signal reg_q2676        : std_logic;
  signal reg_q2676_in     : std_logic;
  		

  -- state q440
  signal reg_q440        : std_logic;
  signal reg_q440_in     : std_logic;
  		

  -- state q442
  signal reg_q442        : std_logic;
  signal reg_q442_in     : std_logic;
  		

  -- state q403
  signal reg_q403        : std_logic;
  signal reg_q403_in     : std_logic;
  		

  -- state q405
  signal reg_q405        : std_logic;
  signal reg_q405_in     : std_logic;
  		

  -- state q1246
  signal reg_q1246        : std_logic;
  signal reg_q1246_in     : std_logic;
  		

  -- state q752
  signal reg_q752        : std_logic;
  signal reg_q752_in     : std_logic;
  		

  -- state q1445
  signal reg_q1445        : std_logic;
  signal reg_q1445_in     : std_logic;
  		

  -- state q2288
  signal reg_q2288        : std_logic;
  signal reg_q2288_in     : std_logic;
  		

  -- state q1490
  signal reg_q1490        : std_logic;
  signal reg_q1490_in     : std_logic;
  		

  -- state q2130
  signal reg_q2130        : std_logic;
  signal reg_q2130_in     : std_logic;
  		

  -- state q2280
  signal reg_q2280        : std_logic;
  signal reg_q2280_in     : std_logic;
  		

  -- state q2282
  signal reg_q2282        : std_logic;
  signal reg_q2282_in     : std_logic;
  		

  -- state q1535
  signal reg_q1535        : std_logic;
  signal reg_q1535_in     : std_logic;
  		

  -- state q1537
  signal reg_q1537        : std_logic;
  signal reg_q1537_in     : std_logic;
  		

  -- state q313
  signal reg_q313        : std_logic;
  signal reg_q313_in     : std_logic;
  		

  -- state q315
  signal reg_q315        : std_logic;
  signal reg_q315_in     : std_logic;
  		

  -- state q1556
  signal reg_q1556        : std_logic;
  signal reg_q1556_in     : std_logic;
  		

  -- state q1558
  signal reg_q1558        : std_logic;
  signal reg_q1558_in     : std_logic;
  		

  -- state q1439
  signal reg_q1439        : std_logic;
  signal reg_q1439_in     : std_logic;
  		

  -- state q2357
  signal reg_q2357        : std_logic;
  signal reg_q2357_in     : std_logic;
  		

  -- state q2359
  signal reg_q2359        : std_logic;
  signal reg_q2359_in     : std_logic;
  		

  -- state q2105
  signal reg_q2105        : std_logic;
  signal reg_q2105_in     : std_logic;
  		

  -- state q2640
  signal reg_q2640        : std_logic;
  signal reg_q2640_in     : std_logic;
  		

  -- state q241
  signal reg_q241        : std_logic;
  signal reg_q241_in     : std_logic;
  		

  -- state q1313
  signal reg_q1313        : std_logic;
  signal reg_q1313_in     : std_logic;
  		

  -- state q1256
  signal reg_q1256        : std_logic;
  signal reg_q1256_in     : std_logic;
  		

  -- state q1033
  signal reg_q1033        : std_logic;
  signal reg_q1033_in     : std_logic;
  		

  -- state q2624
  signal reg_q2624        : std_logic;
  signal reg_q2624_in     : std_logic;
  		

  -- state q974
  signal reg_q974        : std_logic;
  signal reg_q974_in     : std_logic;
  		

  -- state q976
  signal reg_q976        : std_logic;
  signal reg_q976_in     : std_logic;
  		

  -- state q992
  signal reg_q992        : std_logic;
  signal reg_q992_in     : std_logic;
  		

  -- state q298
  signal reg_q298        : std_logic;
  signal reg_q298_in     : std_logic;
  		

  -- state q300
  signal reg_q300        : std_logic;
  signal reg_q300_in     : std_logic;
  		

  -- state q696
  signal reg_q696        : std_logic;
  signal reg_q696_in     : std_logic;
  		

  -- state q1539
  signal reg_q1539        : std_logic;
  signal reg_q1539_in     : std_logic;
  		

  -- state q161
  signal reg_q161        : std_logic;
  signal reg_q161_in     : std_logic;
  		

  -- state q163
  signal reg_q163        : std_logic;
  signal reg_q163_in     : std_logic;
  		

  -- state q2547
  signal reg_q2547        : std_logic;
  signal reg_q2547_in     : std_logic;
  		

  -- state q2549
  signal reg_q2549        : std_logic;
  signal reg_q2549_in     : std_logic;
  		

  -- state q1070
  signal reg_q1070        : std_logic;
  signal reg_q1070_in     : std_logic;
  		

  -- state q438
  signal reg_q438        : std_logic;
  signal reg_q438_in     : std_logic;
  		

  -- state q1710
  signal reg_q1710        : std_logic;
  signal reg_q1710_in     : std_logic;
  		

  -- state q1712
  signal reg_q1712        : std_logic;
  signal reg_q1712_in     : std_logic;
  		

  -- state q407
  signal reg_q407        : std_logic;
  signal reg_q407_in     : std_logic;
  		

  -- state q409
  signal reg_q409        : std_logic;
  signal reg_q409_in     : std_logic;
  		

  -- state q2470
  signal reg_q2470        : std_logic;
  signal reg_q2470_in     : std_logic;
  		

  -- state q2472
  signal reg_q2472        : std_logic;
  signal reg_q2472_in     : std_logic;
  		

  -- state q200
  signal reg_q200        : std_logic;
  signal reg_q200_in     : std_logic;
  		

  -- state q88
  signal reg_q88        : std_logic;
  signal reg_q88_in     : std_logic;
  		

  -- state q1230
  signal reg_q1230        : std_logic;
  signal reg_q1230_in     : std_logic;
  		

  -- state q1232
  signal reg_q1232        : std_logic;
  signal reg_q1232_in     : std_logic;
  		

  -- state q2646
  signal reg_q2646        : std_logic;
  signal reg_q2646_in     : std_logic;
  		

  -- state q2648
  signal reg_q2648        : std_logic;
  signal reg_q2648_in     : std_logic;
  		

  -- state q1254
  signal reg_q1254        : std_logic;
  signal reg_q1254_in     : std_logic;
  		

  -- state q1474
  signal reg_q1474        : std_logic;
  signal reg_q1474_in     : std_logic;
  		

  -- state q66
  signal reg_q66        : std_logic;
  signal reg_q66_in     : std_logic;
  		

  -- state q68
  signal reg_q68        : std_logic;
  signal reg_q68_in     : std_logic;
  		

  -- state q2300
  signal reg_q2300        : std_logic;
  signal reg_q2300_in     : std_logic;
  		

  -- state q2268
  signal reg_q2268        : std_logic;
  signal reg_q2268_in     : std_logic;
  		

  -- state q2270
  signal reg_q2270        : std_logic;
  signal reg_q2270_in     : std_logic;
  		

  -- state q2032
  signal reg_q2032        : std_logic;
  signal reg_q2032_in     : std_logic;
  		

  -- state q2034
  signal reg_q2034        : std_logic;
  signal reg_q2034_in     : std_logic;
  		

  -- state q430
  signal reg_q430        : std_logic;
  signal reg_q430_in     : std_logic;
  		

  -- state q766
  signal reg_q766        : std_logic;
  signal reg_q766_in     : std_logic;
  		

  -- state q768
  signal reg_q768        : std_logic;
  signal reg_q768_in     : std_logic;
  		

  -- state q2662
  signal reg_q2662        : std_logic;
  signal reg_q2662_in     : std_logic;
  		

  -- state q2664
  signal reg_q2664        : std_logic;
  signal reg_q2664_in     : std_logic;
  		

  -- state q139
  signal reg_q139        : std_logic;
  signal reg_q139_in     : std_logic;
  		

  -- state q1141
  signal reg_q1141        : std_logic;
  signal reg_q1141_in     : std_logic;
  		

  -- state q2010
  signal reg_q2010        : std_logic;
  signal reg_q2010_in     : std_logic;
  		

  -- state q2012
  signal reg_q2012        : std_logic;
  signal reg_q2012_in     : std_logic;
  		

  -- state q1068
  signal reg_q1068        : std_logic;
  signal reg_q1068_in     : std_logic;
  		

  -- state q2557
  signal reg_q2557        : std_logic;
  signal reg_q2557_in     : std_logic;
  		

  -- state q2559
  signal reg_q2559        : std_logic;
  signal reg_q2559_in     : std_logic;
  		

  -- state q1617
  signal reg_q1617        : std_logic;
  signal reg_q1617_in     : std_logic;
  		

  -- state q1619
  signal reg_q1619        : std_logic;
  signal reg_q1619_in     : std_logic;
  		

  -- state q1258
  signal reg_q1258        : std_logic;
  signal reg_q1258_in     : std_logic;
  		

  -- state q1260
  signal reg_q1260        : std_logic;
  signal reg_q1260_in     : std_logic;
  		

  -- state q734
  signal reg_q734        : std_logic;
  signal reg_q734_in     : std_logic;
  		

  -- state q1447
  signal reg_q1447        : std_logic;
  signal reg_q1447_in     : std_logic;
  		

  -- state q2014
  signal reg_q2014        : std_logic;
  signal reg_q2014_in     : std_logic;
  		

  -- state q2502
  signal reg_q2502        : std_logic;
  signal reg_q2502_in     : std_logic;
  		

  -- state q2296
  signal reg_q2296        : std_logic;
  signal reg_q2296_in     : std_logic;
  		

  -- state q2298
  signal reg_q2298        : std_logic;
  signal reg_q2298_in     : std_logic;
  		

  -- state q1159
  signal reg_q1159        : std_logic;
  signal reg_q1159_in     : std_logic;
  		

  -- state q444
  signal reg_q444        : std_logic;
  signal reg_q444_in     : std_logic;
  		

  -- state q446
  signal reg_q446        : std_logic;
  signal reg_q446_in     : std_logic;
  		

  -- state q1183
  signal reg_q1183        : std_logic;
  signal reg_q1183_in     : std_logic;
  		

  -- state q1185
  signal reg_q1185        : std_logic;
  signal reg_q1185_in     : std_logic;
  		

  -- state q962
  signal reg_q962        : std_logic;
  signal reg_q962_in     : std_logic;
  		

  -- state q2573
  signal reg_q2573        : std_logic;
  signal reg_q2573_in     : std_logic;
  		

  -- state q1123
  signal reg_q1123        : std_logic;
  signal reg_q1123_in     : std_logic;
  		

  -- state q1125
  signal reg_q1125        : std_logic;
  signal reg_q1125_in     : std_logic;
  		

  -- state q1613
  signal reg_q1613        : std_logic;
  signal reg_q1613_in     : std_logic;
  		

  -- state q2339
  signal reg_q2339        : std_logic;
  signal reg_q2339_in     : std_logic;
  		

  -- state q667
  signal reg_q667        : std_logic;
  signal reg_q667_in     : std_logic;
  		

  -- state q60
  signal reg_q60        : std_logic;
  signal reg_q60_in     : std_logic;
  		

  -- state q399
  signal reg_q399        : std_logic;
  signal reg_q399_in     : std_logic;
  		

  -- state q2650
  signal reg_q2650        : std_logic;
  signal reg_q2650_in     : std_logic;
  		

  -- state q1076
  signal reg_q1076        : std_logic;
  signal reg_q1076_in     : std_logic;
  		

  -- state q1078
  signal reg_q1078        : std_logic;
  signal reg_q1078_in     : std_logic;
  		

  -- state q284
  signal reg_q284        : std_logic;
  signal reg_q284_in     : std_logic;
  		

  -- state q2095
  signal reg_q2095        : std_logic;
  signal reg_q2095_in     : std_logic;
  		

  -- state q171
  signal reg_q171        : std_logic;
  signal reg_q171_in     : std_logic;
  		

  -- state q239
  signal reg_q239        : std_logic;
  signal reg_q239_in     : std_logic;
  		

  -- state q278
  signal reg_q278        : std_logic;
  signal reg_q278_in     : std_logic;
  		

  -- state q105
  signal reg_q105        : std_logic;
  signal reg_q105_in     : std_logic;
  		

  -- state q2148
  signal reg_q2148        : std_logic;
  signal reg_q2148_in     : std_logic;
  		

  -- state q1343
  signal reg_q1343        : std_logic;
  signal reg_q1343_in     : std_logic;
  		

  -- state q1625
  signal reg_q1625        : std_logic;
  signal reg_q1625_in     : std_logic;
  		

  -- state q1627
  signal reg_q1627        : std_logic;
  signal reg_q1627_in     : std_logic;
  		

  -- state q349
  signal reg_q349        : std_logic;
  signal reg_q349_in     : std_logic;
  		

  -- state q351
  signal reg_q351        : std_logic;
  signal reg_q351_in     : std_logic;
  		

  -- state q1648
  signal reg_q1648        : std_logic;
  signal reg_q1648_in     : std_logic;
  		

  -- state q307
  signal reg_q307        : std_logic;
  signal reg_q307_in     : std_logic;
  		

  -- state q2290
  signal reg_q2290        : std_logic;
  signal reg_q2290_in     : std_logic;
  		

  -- state q1533
  signal reg_q1533        : std_logic;
  signal reg_q1533_in     : std_logic;
  		

  -- state q2237
  signal reg_q2237        : std_logic;
  signal reg_q2237_in     : std_logic;
  		

  -- state q2239
  signal reg_q2239        : std_logic;
  signal reg_q2239_in     : std_logic;
  		

  -- state q1242
  signal reg_q1242        : std_logic;
  signal reg_q1242_in     : std_logic;
  		

  -- state q1244
  signal reg_q1244        : std_logic;
  signal reg_q1244_in     : std_logic;
  		

  -- state q1282
  signal reg_q1282        : std_logic;
  signal reg_q1282_in     : std_logic;
  		

  -- state q1284
  signal reg_q1284        : std_logic;
  signal reg_q1284_in     : std_logic;
  		

  -- state q1570
  signal reg_q1570        : std_logic;
  signal reg_q1570_in     : std_logic;
  		

  -- state q1572
  signal reg_q1572        : std_logic;
  signal reg_q1572_in     : std_logic;
  		

  -- state q1706
  signal reg_q1706        : std_logic;
  signal reg_q1706_in     : std_logic;
  		

  -- state q436
  signal reg_q436        : std_logic;
  signal reg_q436_in     : std_logic;
  		

  -- state q220
  signal reg_q220        : std_logic;
  signal reg_q220_in     : std_logic;
  		

  -- state q222
  signal reg_q222        : std_logic;
  signal reg_q222_in     : std_logic;
  		

  -- state q210
  signal reg_q210        : std_logic;
  signal reg_q210_in     : std_logic;
  		

  -- state q212
  signal reg_q212        : std_logic;
  signal reg_q212_in     : std_logic;
  		

  -- state q78
  signal reg_q78        : std_logic;
  signal reg_q78_in     : std_logic;
  		

  -- state q80
  signal reg_q80        : std_logic;
  signal reg_q80_in     : std_logic;
  		

  -- state q684
  signal reg_q684        : std_logic;
  signal reg_q684_in     : std_logic;
  		

  -- state q1039
  signal reg_q1039        : std_logic;
  signal reg_q1039_in     : std_logic;
  		

  -- state q1041
  signal reg_q1041        : std_logic;
  signal reg_q1041_in     : std_logic;
  		

  -- state q2241
  signal reg_q2241        : std_logic;
  signal reg_q2241_in     : std_logic;
  		

  -- state q2233
  signal reg_q2233        : std_logic;
  signal reg_q2233_in     : std_logic;
  		

  -- state q2235
  signal reg_q2235        : std_logic;
  signal reg_q2235_in     : std_logic;
  		

  -- state q972
  signal reg_q972        : std_logic;
  signal reg_q972_in     : std_logic;
  		

  -- state q2219
  signal reg_q2219        : std_logic;
  signal reg_q2219_in     : std_logic;
  		

  -- state q1492
  signal reg_q1492        : std_logic;
  signal reg_q1492_in     : std_logic;
  		

  -- state q1554
  signal reg_q1554        : std_logic;
  signal reg_q1554_in     : std_logic;
  		

  -- state q2495
  signal reg_q2495        : std_logic;
  signal reg_q2495_in     : std_logic;
  		

  -- state q2231
  signal reg_q2231        : std_logic;
  signal reg_q2231_in     : std_logic;
  		

  -- state q724
  signal reg_q724        : std_logic;
  signal reg_q724_in     : std_logic;
  		

  -- state q726
  signal reg_q726        : std_logic;
  signal reg_q726_in     : std_logic;
  		

  -- state q2113
  signal reg_q2113        : std_logic;
  signal reg_q2113_in     : std_logic;
  		

  -- state q2144
  signal reg_q2144        : std_logic;
  signal reg_q2144_in     : std_logic;
  		

  -- state q2146
  signal reg_q2146        : std_logic;
  signal reg_q2146_in     : std_logic;
  		

  -- state q1228
  signal reg_q1228        : std_logic;
  signal reg_q1228_in     : std_logic;
  		

  -- state q1650
  signal reg_q1650        : std_logic;
  signal reg_q1650_in     : std_logic;
  		

  -- state q147
  signal reg_q147        : std_logic;
  signal reg_q147_in     : std_logic;
  		

  -- state q296
  signal reg_q296        : std_logic;
  signal reg_q296_in     : std_logic;
  		

  -- state q1611
  signal reg_q1611        : std_logic;
  signal reg_q1611_in     : std_logic;
  		

  -- state q1169
  signal reg_q1169        : std_logic;
  signal reg_q1169_in     : std_logic;
  		

  -- state q1171
  signal reg_q1171        : std_logic;
  signal reg_q1171_in     : std_logic;
  		

  -- state q1017
  signal reg_q1017        : std_logic;
  signal reg_q1017_in     : std_logic;
  		

  -- state q1019
  signal reg_q1019        : std_logic;
  signal reg_q1019_in     : std_logic;
  		

  -- state q2571
  signal reg_q2571        : std_logic;
  signal reg_q2571_in     : std_logic;
  		

  -- state q1615
  signal reg_q1615        : std_logic;
  signal reg_q1615_in     : std_logic;
  		

  -- state q2561
  signal reg_q2561        : std_logic;
  signal reg_q2561_in     : std_logic;
  		

  -- state q1353
  signal reg_q1353        : std_logic;
  signal reg_q1353_in     : std_logic;
  		

  -- state q1127
  signal reg_q1127        : std_logic;
  signal reg_q1127_in     : std_logic;
  		

  -- state q1129
  signal reg_q1129        : std_logic;
  signal reg_q1129_in     : std_logic;
  		

  -- state q1351
  signal reg_q1351        : std_logic;
  signal reg_q1351_in     : std_logic;
  		

  -- state q385
  signal reg_q385        : std_logic;
  signal reg_q385_in     : std_logic;
  		

  -- state q387
  signal reg_q387        : std_logic;
  signal reg_q387_in     : std_logic;
  		

  -- state q432
  signal reg_q432        : std_logic;
  signal reg_q432_in     : std_logic;
  		

  -- state q2318
  signal reg_q2318        : std_logic;
  signal reg_q2318_in     : std_logic;
  		

  -- state q2320
  signal reg_q2320        : std_logic;
  signal reg_q2320_in     : std_logic;
  		

  -- state q2682
  signal reg_q2682        : std_logic;
  signal reg_q2682_in     : std_logic;
  		

  -- state q2684
  signal reg_q2684        : std_logic;
  signal reg_q2684_in     : std_logic;
  		

  -- state q1514
  signal reg_q1514        : std_logic;
  signal reg_q1514_in     : std_logic;
  		

  -- state q1516
  signal reg_q1516        : std_logic;
  signal reg_q1516_in     : std_logic;
  		

  -- state q2107
  signal reg_q2107        : std_logic;
  signal reg_q2107_in     : std_logic;
  		

  -- state q728
  signal reg_q728        : std_logic;
  signal reg_q728_in     : std_logic;
  		

  -- state q2329
  signal reg_q2329        : std_logic;
  signal reg_q2329_in     : std_logic;
  		

  -- state q2331
  signal reg_q2331        : std_logic;
  signal reg_q2331_in     : std_logic;
  		

  -- state q1157
  signal reg_q1157        : std_logic;
  signal reg_q1157_in     : std_logic;
  		

  -- state q2654
  signal reg_q2654        : std_logic;
  signal reg_q2654_in     : std_logic;
  		

  -- state q2656
  signal reg_q2656        : std_logic;
  signal reg_q2656_in     : std_logic;
  		

  -- state q2607
  signal reg_q2607        : std_logic;
  signal reg_q2607_in     : std_logic;
  		

  -- state q1345
  signal reg_q1345        : std_logic;
  signal reg_q1345_in     : std_logic;
  		

  -- state q347
  signal reg_q347        : std_logic;
  signal reg_q347_in     : std_logic;
  		

  -- state q1488
  signal reg_q1488        : std_logic;
  signal reg_q1488_in     : std_logic;
  		

  -- state q1286
  signal reg_q1286        : std_logic;
  signal reg_q1286_in     : std_logic;
  		

  -- state q321
  signal reg_q321        : std_logic;
  signal reg_q321_in     : std_logic;
  		

  -- state q1508
  signal reg_q1508        : std_logic;
  signal reg_q1508_in     : std_logic;
  		

  -- state q1510
  signal reg_q1510        : std_logic;
  signal reg_q1510_in     : std_logic;
  		

  -- state q2099
  signal reg_q2099        : std_logic;
  signal reg_q2099_in     : std_logic;
  		

  -- state q70
  signal reg_q70        : std_logic;
  signal reg_q70_in     : std_logic;
  		

  -- state q970
  signal reg_q970        : std_logic;
  signal reg_q970_in     : std_logic;
  		

  -- state q760
  signal reg_q760        : std_logic;
  signal reg_q760_in     : std_logic;
  		

  -- state q762
  signal reg_q762        : std_logic;
  signal reg_q762_in     : std_logic;
  		

  -- state q707
  signal reg_q707        : std_logic;
  signal reg_q707_in     : std_logic;
  		

  -- state q1234
  signal reg_q1234        : std_logic;
  signal reg_q1234_in     : std_logic;
  		

  -- state q1173
  signal reg_q1173        : std_logic;
  signal reg_q1173_in     : std_logic;
  		

  -- state q1175
  signal reg_q1175        : std_logic;
  signal reg_q1175_in     : std_logic;
  		

  -- state q2512
  signal reg_q2512        : std_logic;
  signal reg_q2512_in     : std_logic;
  		

  -- state q2652
  signal reg_q2652        : std_logic;
  signal reg_q2652_in     : std_logic;
  		

  -- state q1584
  signal reg_q1584        : std_logic;
  signal reg_q1584_in     : std_logic;
  		

  -- state q1006
  signal reg_q1006        : std_logic;
  signal reg_q1006_in     : std_logic;
  		

  -- state q1486
  signal reg_q1486        : std_logic;
  signal reg_q1486_in     : std_logic;
  		

  -- state q331
  signal reg_q331        : std_logic;
  signal reg_q331_in     : std_logic;
  		

  -- state q1270
  signal reg_q1270        : std_logic;
  signal reg_q1270_in     : std_logic;
  		

  -- state q141
  signal reg_q141        : std_logic;
  signal reg_q141_in     : std_logic;
  		

  -- state q143
  signal reg_q143        : std_logic;
  signal reg_q143_in     : std_logic;
  		

  -- state q353
  signal reg_q353        : std_logic;
  signal reg_q353_in     : std_logic;
  		

  -- state q355
  signal reg_q355        : std_logic;
  signal reg_q355_in     : std_logic;
  		

  -- state q2668
  signal reg_q2668        : std_logic;
  signal reg_q2668_in     : std_logic;
  		

  -- state q72
  signal reg_q72        : std_logic;
  signal reg_q72_in     : std_logic;
  		

  -- state q165
  signal reg_q165        : std_logic;
  signal reg_q165_in     : std_logic;
  		

  -- state q1454
  signal reg_q1454        : std_logic;
  signal reg_q1454_in     : std_logic;
  		

  -- state q1456
  signal reg_q1456        : std_logic;
  signal reg_q1456_in     : std_logic;
  		

  -- state q1607
  signal reg_q1607        : std_logic;
  signal reg_q1607_in     : std_logic;
  		

  -- state q1131
  signal reg_q1131        : std_logic;
  signal reg_q1131_in     : std_logic;
  		

  -- state q907
  signal reg_q907        : std_logic;
  signal reg_q907_in     : std_logic;
  		

  -- state q2254
  signal reg_q2254        : std_logic;
  signal reg_q2254_in     : std_logic;
  		

  -- state q2256
  signal reg_q2256        : std_logic;
  signal reg_q2256_in     : std_logic;
  		

  -- state q1629
  signal reg_q1629        : std_logic;
  signal reg_q1629_in     : std_logic;
  		

  -- state q1631
  signal reg_q1631        : std_logic;
  signal reg_q1631_in     : std_logic;
  		

  -- state q157
  signal reg_q157        : std_logic;
  signal reg_q157_in     : std_logic;
  		

  -- state q159
  signal reg_q159        : std_logic;
  signal reg_q159_in     : std_logic;
  		

  -- state q1590
  signal reg_q1590        : std_logic;
  signal reg_q1590_in     : std_logic;
  		

  -- state q1592
  signal reg_q1592        : std_logic;
  signal reg_q1592_in     : std_logic;
  		

  -- state q1564
  signal reg_q1564        : std_logic;
  signal reg_q1564_in     : std_logic;
  		

  -- state q1566
  signal reg_q1566        : std_logic;
  signal reg_q1566_in     : std_logic;
  		

  -- state q1720
  signal reg_q1720        : std_logic;
  signal reg_q1720_in     : std_logic;
  		

  -- state q1722
  signal reg_q1722        : std_logic;
  signal reg_q1722_in     : std_logic;
  		

  -- state q2006
  signal reg_q2006        : std_logic;
  signal reg_q2006_in     : std_logic;
  		

  -- state q1965
  signal reg_q1965        : std_logic;
  signal reg_q1965_in     : std_logic;
  		

  -- state q1967
  signal reg_q1967        : std_logic;
  signal reg_q1967_in     : std_logic;
  		

  -- state q272
  signal reg_q272        : std_logic;
  signal reg_q272_in     : std_logic;
  		

  -- state q274
  signal reg_q274        : std_logic;
  signal reg_q274_in     : std_logic;
  		

  -- state q2264
  signal reg_q2264        : std_logic;
  signal reg_q2264_in     : std_logic;
  		

  -- state q2266
  signal reg_q2266        : std_logic;
  signal reg_q2266_in     : std_logic;
  		

  -- state q204
  signal reg_q204        : std_logic;
  signal reg_q204_in     : std_logic;
  		

  -- state q206
  signal reg_q206        : std_logic;
  signal reg_q206_in     : std_logic;
  		

  -- state q1311
  signal reg_q1311        : std_logic;
  signal reg_q1311_in     : std_logic;
  		

  -- state q909
  signal reg_q909        : std_logic;
  signal reg_q909_in     : std_logic;
  		

  -- state q911
  signal reg_q911        : std_logic;
  signal reg_q911_in     : std_logic;
  		

  -- state q2164
  signal reg_q2164        : std_logic;
  signal reg_q2164_in     : std_logic;
  		

  -- state q2166
  signal reg_q2166        : std_logic;
  signal reg_q2166_in     : std_logic;
  		

  -- state q1098
  signal reg_q1098        : std_logic;
  signal reg_q1098_in     : std_logic;
  		

  -- state q2563
  signal reg_q2563        : std_logic;
  signal reg_q2563_in     : std_logic;
  		

  -- state q2121
  signal reg_q2121        : std_logic;
  signal reg_q2121_in     : std_logic;
  		

  -- state q151
  signal reg_q151        : std_logic;
  signal reg_q151_in     : std_logic;
  		

  -- state q1121
  signal reg_q1121        : std_logic;
  signal reg_q1121_in     : std_logic;
  		

  -- state q243
  signal reg_q243        : std_logic;
  signal reg_q243_in     : std_logic;
  		

  -- state q1043
  signal reg_q1043        : std_logic;
  signal reg_q1043_in     : std_logic;
  		

  -- state q1045
  signal reg_q1045        : std_logic;
  signal reg_q1045_in     : std_logic;
  		

  -- state q276
  signal reg_q276        : std_logic;
  signal reg_q276_in     : std_logic;
  		

  -- state q1047
  signal reg_q1047        : std_logic;
  signal reg_q1047_in     : std_logic;
  		

  -- state q2367
  signal reg_q2367        : std_logic;
  signal reg_q2367_in     : std_logic;
  		

  -- state q1066
  signal reg_q1066        : std_logic;
  signal reg_q1066_in     : std_logic;
  		

  -- state q1496
  signal reg_q1496        : std_logic;
  signal reg_q1496_in     : std_logic;
  		

  -- state q1498
  signal reg_q1498        : std_logic;
  signal reg_q1498_in     : std_logic;
  		

  -- state q1696
  signal reg_q1696        : std_logic;
  signal reg_q1696_in     : std_logic;
  		

  -- state q1494
  signal reg_q1494        : std_logic;
  signal reg_q1494_in     : std_logic;
  		

  -- state q2036
  signal reg_q2036        : std_logic;
  signal reg_q2036_in     : std_logic;
  		

  -- state q1684
  signal reg_q1684        : std_logic;
  signal reg_q1684_in     : std_logic;
  		

  -- state q337
  signal reg_q337        : std_logic;
  signal reg_q337_in     : std_logic;
  		

  -- state q339
  signal reg_q339        : std_logic;
  signal reg_q339_in     : std_logic;
  		

  -- state q1959
  signal reg_q1959        : std_logic;
  signal reg_q1959_in     : std_logic;
  		

  -- state q1961
  signal reg_q1961        : std_logic;
  signal reg_q1961_in     : std_logic;
  		

  -- state q1518
  signal reg_q1518        : std_logic;
  signal reg_q1518_in     : std_logic;
  		

  -- state q1656
  signal reg_q1656        : std_logic;
  signal reg_q1656_in     : std_logic;
  		

  -- state q1658
  signal reg_q1658        : std_logic;
  signal reg_q1658_in     : std_logic;
  		

  -- state q2314
  signal reg_q2314        : std_logic;
  signal reg_q2314_in     : std_logic;
  		

  -- state q2316
  signal reg_q2316        : std_logic;
  signal reg_q2316_in     : std_logic;
  		

  -- state q2638
  signal reg_q2638        : std_logic;
  signal reg_q2638_in     : std_logic;
  		

  -- state q2142
  signal reg_q2142        : std_logic;
  signal reg_q2142_in     : std_logic;
  		

  -- state q2660
  signal reg_q2660        : std_logic;
  signal reg_q2660_in     : std_logic;
  		

  -- state q1568
  signal reg_q1568        : std_logic;
  signal reg_q1568_in     : std_logic;
  		

  -- state q1062
  signal reg_q1062        : std_logic;
  signal reg_q1062_in     : std_logic;
  		

  -- state q1064
  signal reg_q1064        : std_logic;
  signal reg_q1064_in     : std_logic;
  		

  -- state q1686
  signal reg_q1686        : std_logic;
  signal reg_q1686_in     : std_logic;
  		

  -- state q1240
  signal reg_q1240        : std_logic;
  signal reg_q1240_in     : std_logic;
  		

  -- state q764
  signal reg_q764        : std_logic;
  signal reg_q764_in     : std_logic;
  		

  -- state q1119
  signal reg_q1119        : std_logic;
  signal reg_q1119_in     : std_logic;
  		

  -- state q1476
  signal reg_q1476        : std_logic;
  signal reg_q1476_in     : std_logic;
  		

  -- state q62
  signal reg_q62        : std_logic;
  signal reg_q62_in     : std_logic;
  		

  -- state q2678
  signal reg_q2678        : std_logic;
  signal reg_q2678_in     : std_logic;
  		

  -- state q327
  signal reg_q327        : std_logic;
  signal reg_q327_in     : std_logic;
  		

  -- state q329
  signal reg_q329        : std_logic;
  signal reg_q329_in     : std_logic;
  		

  -- state q1718
  signal reg_q1718        : std_logic;
  signal reg_q1718_in     : std_logic;
  		

  -- state q1054
  signal reg_q1054        : std_logic;
  signal reg_q1054_in     : std_logic;
  		

  -- state q1056
  signal reg_q1056        : std_logic;
  signal reg_q1056_in     : std_logic;
  		

  -- state q1512
  signal reg_q1512        : std_logic;
  signal reg_q1512_in     : std_logic;
  		

  -- state q2262
  signal reg_q2262        : std_logic;
  signal reg_q2262_in     : std_logic;
  		

  -- state q1167
  signal reg_q1167        : std_logic;
  signal reg_q1167_in     : std_logic;
  		

  -- state q2379
  signal reg_q2379        : std_logic;
  signal reg_q2379_in     : std_logic;
  		

  -- state q2016
  signal reg_q2016        : std_logic;
  signal reg_q2016_in     : std_logic;
  		

  -- state q64
  signal reg_q64        : std_logic;
  signal reg_q64_in     : std_logic;
  		

  -- state q1623
  signal reg_q1623        : std_logic;
  signal reg_q1623_in     : std_logic;
  		

  -- state q145
  signal reg_q145        : std_logic;
  signal reg_q145_in     : std_logic;
  		

  -- state q1594
  signal reg_q1594        : std_logic;
  signal reg_q1594_in     : std_logic;
  		

  -- state q1596
  signal reg_q1596        : std_logic;
  signal reg_q1596_in     : std_logic;
  		

  -- state q2626
  signal reg_q2626        : std_logic;
  signal reg_q2626_in     : std_logic;
  		

  -- state q2365
  signal reg_q2365        : std_logic;
  signal reg_q2365_in     : std_logic;
  		

  -- state q1609
  signal reg_q1609        : std_logic;
  signal reg_q1609_in     : std_logic;
  		

  -- state q1058
  signal reg_q1058        : std_logic;
  signal reg_q1058_in     : std_logic;
  		

  -- state q1060
  signal reg_q1060        : std_logic;
  signal reg_q1060_in     : std_logic;
  		

  -- state q208
  signal reg_q208        : std_logic;
  signal reg_q208_in     : std_logic;
  		

  -- state q1621
  signal reg_q1621        : std_logic;
  signal reg_q1621_in     : std_logic;
  		

  -- state q694
  signal reg_q694        : std_logic;
  signal reg_q694_in     : std_logic;
  		

  -- state q214
  signal reg_q214        : std_logic;
  signal reg_q214_in     : std_logic;
  		

  -- state q2555
  signal reg_q2555        : std_logic;
  signal reg_q2555_in     : std_logic;
  		

  -- state q2152
  signal reg_q2152        : std_logic;
  signal reg_q2152_in     : std_logic;
  		

  -- state q2154
  signal reg_q2154        : std_logic;
  signal reg_q2154_in     : std_logic;
  		

  -- state q2312
  signal reg_q2312        : std_logic;
  signal reg_q2312_in     : std_logic;
  		

  -- state q311
  signal reg_q311        : std_logic;
  signal reg_q311_in     : std_logic;
  		

  -- state q1500
  signal reg_q1500        : std_logic;
  signal reg_q1500_in     : std_logic;
  		

  -- state q317
  signal reg_q317        : std_logic;
  signal reg_q317_in     : std_logic;
  		

  -- state q2680
  signal reg_q2680        : std_logic;
  signal reg_q2680_in     : std_logic;
  		

  -- state q1266
  signal reg_q1266        : std_logic;
  signal reg_q1266_in     : std_logic;
  		

  -- state q1268
  signal reg_q1268        : std_logic;
  signal reg_q1268_in     : std_logic;
  		

  -- state q2628
  signal reg_q2628        : std_logic;
  signal reg_q2628_in     : std_logic;
  		

  -- state q2630
  signal reg_q2630        : std_logic;
  signal reg_q2630_in     : std_logic;
  		

  -- state q1429
  signal reg_q1429        : std_logic;
  signal reg_q1429_in     : std_logic;
  		

  -- state q1236
  signal reg_q1236        : std_logic;
  signal reg_q1236_in     : std_logic;
  		

  -- state q1238
  signal reg_q1238        : std_logic;
  signal reg_q1238_in     : std_logic;
  		

  -- state q2478
  signal reg_q2478        : std_logic;
  signal reg_q2478_in     : std_logic;
  		

  -- state q722
  signal reg_q722        : std_logic;
  signal reg_q722_in     : std_logic;
  		

  -- state q391
  signal reg_q391        : std_logic;
  signal reg_q391_in     : std_logic;
  		

  -- state q393
  signal reg_q393        : std_logic;
  signal reg_q393_in     : std_logic;
  		

  -- state q1280
  signal reg_q1280        : std_logic;
  signal reg_q1280_in     : std_logic;
  		

  -- state q2569
  signal reg_q2569        : std_logic;
  signal reg_q2569_in     : std_logic;
  		

  -- state q202
  signal reg_q202        : std_logic;
  signal reg_q202_in     : std_logic;
  		

  -- state q268
  signal reg_q268        : std_logic;
  signal reg_q268_in     : std_logic;
  		

  -- state q270
  signal reg_q270        : std_logic;
  signal reg_q270_in     : std_logic;
  		

  -- state q173
  signal reg_q173        : std_logic;
  signal reg_q173_in     : std_logic;
  		

  -- state q175
  signal reg_q175        : std_logic;
  signal reg_q175_in     : std_logic;
  		

  -- state q669
  signal reg_q669        : std_logic;
  signal reg_q669_in     : std_logic;
  		

  -- state q1502
  signal reg_q1502        : std_logic;
  signal reg_q1502_in     : std_logic;
  		

  -- state q738
  signal reg_q738        : std_logic;
  signal reg_q738_in     : std_logic;
  		

  -- state q54
  signal reg_q54        : std_logic;
  signal reg_q54_in     : std_logic;
  		

  -- state q1963
  signal reg_q1963        : std_logic;
  signal reg_q1963_in     : std_logic;
  		

  -- state q2381
  signal reg_q2381        : std_logic;
  signal reg_q2381_in     : std_logic;
  		

  -- state q2345
  signal reg_q2345        : std_logic;
  signal reg_q2345_in     : std_logic;
  		

  -- state q2008
  signal reg_q2008        : std_logic;
  signal reg_q2008_in     : std_logic;
  		

  -- state q730
  signal reg_q730        : std_logic;
  signal reg_q730_in     : std_logic;
  		

  -- state q1321
  signal reg_q1321        : std_logic;
  signal reg_q1321_in     : std_logic;
  		

  -- state q1323
  signal reg_q1323        : std_logic;
  signal reg_q1323_in     : std_logic;
  		

  -- state q1309
  signal reg_q1309        : std_logic;
  signal reg_q1309_in     : std_logic;
  		

  -- state q99
  signal reg_q99        : std_logic;
  signal reg_q99_in     : std_logic;
  		

  -- state q1586
  signal reg_q1586        : std_logic;
  signal reg_q1586_in     : std_logic;
  		

  -- state q2156
  signal reg_q2156        : std_logic;
  signal reg_q2156_in     : std_logic;
  		

  -- state q319
  signal reg_q319        : std_logic;
  signal reg_q319_in     : std_logic;
  		

  -- state q2026
  signal reg_q2026        : std_logic;
  signal reg_q2026_in     : std_logic;
  		

  -- state q401
  signal reg_q401        : std_logic;
  signal reg_q401_in     : std_logic;
  		

  -- state q2666
  signal reg_q2666        : std_logic;
  signal reg_q2666_in     : std_logic;
  		

  -- state q286
  signal reg_q286        : std_logic;
  signal reg_q286_in     : std_logic;
  		

  -- state q2658
  signal reg_q2658        : std_logic;
  signal reg_q2658_in     : std_logic;
  		

  -- state q754
  signal reg_q754        : std_logic;
  signal reg_q754_in     : std_logic;
  		

  -- state q345
  signal reg_q345        : std_logic;
  signal reg_q345_in     : std_logic;
  		

  -- state q1021
  signal reg_q1021        : std_logic;
  signal reg_q1021_in     : std_logic;
  		

  -- state q2539
  signal reg_q2539        : std_logic;
  signal reg_q2539_in     : std_logic;
  		

  -- state q1163
  signal reg_q1163        : std_logic;
  signal reg_q1163_in     : std_logic;
  		

  -- state q1165
  signal reg_q1165        : std_logic;
  signal reg_q1165_in     : std_logic;
  		

  -- state q411
  signal reg_q411        : std_logic;
  signal reg_q411_in     : std_logic;
  		

  -- state q720
  signal reg_q720        : std_logic;
  signal reg_q720_in     : std_logic;
  		

  -- state q1292
  signal reg_q1292        : std_logic;
  signal reg_q1292_in     : std_logic;
  		

  -- state q1294
  signal reg_q1294        : std_logic;
  signal reg_q1294_in     : std_logic;
  		

  -- state q2553
  signal reg_q2553        : std_logic;
  signal reg_q2553_in     : std_logic;
  		

  -- state q1449
  signal reg_q1449        : std_logic;
  signal reg_q1449_in     : std_logic;
  		

  -- state q1100
  signal reg_q1100        : std_logic;
  signal reg_q1100_in     : std_logic;
  		

  -- state q424
  signal reg_q424        : std_logic;
  signal reg_q424_in     : std_logic;
  		

  -- state q1177
  signal reg_q1177        : std_logic;
  signal reg_q1177_in     : std_logic;
  		

  -- state q2355
  signal reg_q2355        : std_logic;
  signal reg_q2355_in     : std_logic;
  		

  -- state q732
  signal reg_q732        : std_logic;
  signal reg_q732_in     : std_logic;
  		

  -- state q434
  signal reg_q434        : std_logic;
  signal reg_q434_in     : std_logic;
  		

  -- state q2551
  signal reg_q2551        : std_logic;
  signal reg_q2551_in     : std_logic;
  		

  -- state q2044
  signal reg_q2044        : std_logic;
  signal reg_q2044_in     : std_logic;
  		

  -- state q2046
  signal reg_q2046        : std_logic;
  signal reg_q2046_in     : std_logic;
  		

  -- state q2541
  signal reg_q2541        : std_logic;
  signal reg_q2541_in     : std_logic;
  		

  -- state q1588
  signal reg_q1588        : std_logic;
  signal reg_q1588_in     : std_logic;
  		

  -- state q2693
  signal reg_q2693        : std_logic;
  signal reg_q2693_in     : std_logic;
  		

  -- state q2543
  signal reg_q2543        : std_logic;
  signal reg_q2543_in     : std_logic;
  		

  -- state q2545
  signal reg_q2545        : std_logic;
  signal reg_q2545_in     : std_logic;
  		

  -- state q2347
  signal reg_q2347        : std_logic;
  signal reg_q2347_in     : std_logic;
  		

  -- state q1740
  signal reg_q1740        : std_logic;
  signal reg_q1740_in     : std_logic;
  		

  -- state q1329
  signal reg_q1329        : std_logic;
  signal reg_q1329_in     : std_logic;
  		

  -- state q2632
  signal reg_q2632        : std_logic;
  signal reg_q2632_in     : std_logic;
  		

  -- state q1303
  signal reg_q1303        : std_logic;
  signal reg_q1303_in     : std_logic;
  		

  -- state q309
  signal reg_q309        : std_logic;
  signal reg_q309_in     : std_logic;
  		

  -- state q216
  signal reg_q216        : std_logic;
  signal reg_q216_in     : std_logic;
  		

  -- state q2134
  signal reg_q2134        : std_logic;
  signal reg_q2134_in     : std_logic;
  		

  -- state q770
  signal reg_q770        : std_logic;
  signal reg_q770_in     : std_logic;
  		

  -- state q155
  signal reg_q155        : std_logic;
  signal reg_q155_in     : std_logic;
  		

  -- state q2140
  signal reg_q2140        : std_logic;
  signal reg_q2140_in     : std_logic;
  		

  -- state q383
  signal reg_q383        : std_logic;
  signal reg_q383_in     : std_logic;
  		

  -- state q1633
  signal reg_q1633        : std_logic;
  signal reg_q1633_in     : std_logic;
  		

  -- state q772
  signal reg_q772        : std_logic;
  signal reg_q772_in     : std_logic;
  		

  -- state q1155
  signal reg_q1155        : std_logic;
  signal reg_q1155_in     : std_logic;
  		

  -- state q927
  signal reg_q927        : std_logic;
  signal reg_q927_in     : std_logic;
  		

  -- state q929
  signal reg_q929        : std_logic;
  signal reg_q929_in     : std_logic;
  		

  -- state q1969
  signal reg_q1969        : std_logic;
  signal reg_q1969_in     : std_logic;
  		

  -- state q1415
  signal reg_q1415        : std_logic;
  signal reg_q1415_in     : std_logic;
  		

  -- state q1417
  signal reg_q1417        : std_logic;
  signal reg_q1417_in     : std_logic;
  		

  -- state q153
  signal reg_q153        : std_logic;
  signal reg_q153_in     : std_logic;
  		

  -- state q1288
  signal reg_q1288        : std_logic;
  signal reg_q1288_in     : std_logic;
  		

  -- state q1276
  signal reg_q1276        : std_logic;
  signal reg_q1276_in     : std_logic;
  		

  -- state q2048
  signal reg_q2048        : std_logic;
  signal reg_q2048_in     : std_logic;
  		

  -- state q218
  signal reg_q218        : std_logic;
  signal reg_q218_in     : std_logic;
  		

  -- state q1149
  signal reg_q1149        : std_logic;
  signal reg_q1149_in     : std_logic;
  		

  -- state q259
  signal reg_q259        : std_logic;
  signal reg_q259_in     : std_logic;
  		

  -- state q2327
  signal reg_q2327        : std_logic;
  signal reg_q2327_in     : std_logic;
  		

  -- state q266
  signal reg_q266        : std_logic;
  signal reg_q266_in     : std_logic;
  		

  -- state q746
  signal reg_q746        : std_logic;
  signal reg_q746_in     : std_logic;
  		

  -- state q774
  signal reg_q774        : std_logic;
  signal reg_q774_in     : std_logic;
  		

  -- state q776
  signal reg_q776        : std_logic;
  signal reg_q776_in     : std_logic;
  		

  -- state q389
  signal reg_q389        : std_logic;
  signal reg_q389_in     : std_logic;
  		

  -- state q1598
  signal reg_q1598        : std_logic;
  signal reg_q1598_in     : std_logic;
  		

  -- state q1004
  signal reg_q1004        : std_logic;
  signal reg_q1004_in     : std_logic;
  		

  -- state q1419
  signal reg_q1419        : std_logic;
  signal reg_q1419_in     : std_logic;
  		

  -- state q1278
  signal reg_q1278        : std_logic;
  signal reg_q1278_in     : std_logic;
  		

  -- state q1654
  signal reg_q1654        : std_logic;
  signal reg_q1654_in     : std_logic;
  		

  -- state q1458
  signal reg_q1458        : std_logic;
  signal reg_q1458_in     : std_logic;
  		

  -- state q1641
  signal reg_q1641        : std_logic;
  signal reg_q1641_in     : std_logic;
  		

  -- state q1600
  signal reg_q1600        : std_logic;
  signal reg_q1600_in     : std_logic;
  		

  -- state q2097
  signal reg_q2097        : std_logic;
  signal reg_q2097_in     : std_logic;
  		

  -- state q1290
  signal reg_q1290        : std_logic;
  signal reg_q1290_in     : std_logic;
  		

  -- state q740
  signal reg_q740        : std_logic;
  signal reg_q740_in     : std_logic;
  		

  -- state q677
  signal reg_q677        : std_logic;
  signal reg_q677_in     : std_logic;
  		

  -- state q2050
  signal reg_q2050        : std_logic;
  signal reg_q2050_in     : std_logic;
  		
  signal reg_fullgraph2       : std_logic_vector(9 downto 0);
  signal reg_fullgraph2_in    : std_logic_vector(9 downto 0);
  signal reg_fullgraph2_init  : std_logic_vector(9 downto 0);
  signal reg_fullgraph2_sel   : std_logic_vector(1023 downto 0); 	
  -- end section fullgraph2
  --#################################################			
		

  -- state q178
  signal reg_q178        : std_logic;
  signal reg_q178_in     : std_logic;
  signal reg_q178_init   : std_logic;
		

  -- state q899
  signal reg_q899        : std_logic;
  signal reg_q899_in     : std_logic;
  signal reg_q899_init   : std_logic;
		

  -- state q225
  signal reg_q225        : std_logic;
  signal reg_q225_in     : std_logic;
  signal reg_q225_init   : std_logic;
		

  -- state q1297
  signal reg_q1297        : std_logic;
  signal reg_q1297_in     : std_logic;
  signal reg_q1297_init   : std_logic;
		
--#################################################
-- start section fullgraph: 7

  -- state q1876
  signal reg_q1876        : std_logic;
  signal reg_q1876_in     : std_logic;
  		

  -- state q1878
  signal reg_q1878        : std_logic;
  signal reg_q1878_in     : std_logic;
  		

  -- state q1792
  signal reg_q1792        : std_logic;
  signal reg_q1792_in     : std_logic;
  		

  -- state q1794
  signal reg_q1794        : std_logic;
  signal reg_q1794_in     : std_logic;
  		

  -- state q1852
  signal reg_q1852        : std_logic;
  signal reg_q1852_in     : std_logic;
  		

  -- state q1854
  signal reg_q1854        : std_logic;
  signal reg_q1854_in     : std_logic;
  		

  -- state q889
  signal reg_q889        : std_logic;
  signal reg_q889_in     : std_logic;
  		

  -- state q532
  signal reg_q532        : std_logic;
  signal reg_q532_in     : std_logic;
  		

  -- state q534
  signal reg_q534        : std_logic;
  signal reg_q534_in     : std_logic;
  		

  -- state q2419
  signal reg_q2419        : std_logic;
  signal reg_q2419_in     : std_logic;
  		

  -- state q2421
  signal reg_q2421        : std_logic;
  signal reg_q2421_in     : std_logic;
  		

  -- state q1770
  signal reg_q1770        : std_logic;
  signal reg_q1770_in     : std_logic;
  		

  -- state q616
  signal reg_q616        : std_logic;
  signal reg_q616_in     : std_logic;
  		

  -- state q526
  signal reg_q526        : std_logic;
  signal reg_q526_in     : std_logic;
  		

  -- state q945
  signal reg_q945        : std_logic;
  signal reg_q945_in     : std_logic;
  		

  -- state q947
  signal reg_q947        : std_logic;
  signal reg_q947_in     : std_logic;
  		

  -- state q791
  signal reg_q791        : std_logic;
  signal reg_q791_in     : std_logic;
  		

  -- state q856
  signal reg_q856        : std_logic;
  signal reg_q856_in     : std_logic;
  		

  -- state q858
  signal reg_q858        : std_logic;
  signal reg_q858_in     : std_logic;
  		

  -- state q1215
  signal reg_q1215        : std_logic;
  signal reg_q1215_in     : std_logic;
  		

  -- state q1217
  signal reg_q1217        : std_logic;
  signal reg_q1217_in     : std_logic;
  		

  -- state q937
  signal reg_q937        : std_logic;
  signal reg_q937_in     : std_logic;
  		

  -- state q939
  signal reg_q939        : std_logic;
  signal reg_q939_in     : std_logic;
  		

  -- state q1866
  signal reg_q1866        : std_logic;
  signal reg_q1866_in     : std_logic;
  		

  -- state q2002
  signal reg_q2002        : std_logic;
  signal reg_q2002_in     : std_logic;
  		

  -- state q520
  signal reg_q520        : std_logic;
  signal reg_q520_in     : std_logic;
  		

  -- state q522
  signal reg_q522        : std_logic;
  signal reg_q522_in     : std_logic;
  		

  -- state q2528
  signal reg_q2528        : std_logic;
  signal reg_q2528_in     : std_logic;
  		

  -- state q2530
  signal reg_q2530        : std_logic;
  signal reg_q2530_in     : std_logic;
  		

  -- state q2445
  signal reg_q2445        : std_logic;
  signal reg_q2445_in     : std_logic;
  		

  -- state q2447
  signal reg_q2447        : std_logic;
  signal reg_q2447_in     : std_logic;
  		

  -- state q1874
  signal reg_q1874        : std_logic;
  signal reg_q1874_in     : std_logic;
  		

  -- state q2078
  signal reg_q2078        : std_logic;
  signal reg_q2078_in     : std_logic;
  		

  -- state q2080
  signal reg_q2080        : std_logic;
  signal reg_q2080_in     : std_logic;
  		

  -- state q2178
  signal reg_q2178        : std_logic;
  signal reg_q2178_in     : std_logic;
  		

  -- state q2180
  signal reg_q2180        : std_logic;
  signal reg_q2180_in     : std_logic;
  		

  -- state q590
  signal reg_q590        : std_logic;
  signal reg_q590_in     : std_logic;
  		

  -- state q592
  signal reg_q592        : std_logic;
  signal reg_q592_in     : std_logic;
  		

  -- state q1387
  signal reg_q1387        : std_logic;
  signal reg_q1387_in     : std_logic;
  		

  -- state q1389
  signal reg_q1389        : std_logic;
  signal reg_q1389_in     : std_logic;
  		

  -- state q2405
  signal reg_q2405        : std_logic;
  signal reg_q2405_in     : std_logic;
  		

  -- state q2407
  signal reg_q2407        : std_logic;
  signal reg_q2407_in     : std_logic;
  		

  -- state q1920
  signal reg_q1920        : std_logic;
  signal reg_q1920_in     : std_logic;
  		

  -- state q1409
  signal reg_q1409        : std_logic;
  signal reg_q1409_in     : std_logic;
  		

  -- state q1411
  signal reg_q1411        : std_logic;
  signal reg_q1411_in     : std_logic;
  		

  -- state q2064
  signal reg_q2064        : std_logic;
  signal reg_q2064_in     : std_logic;
  		

  -- state q960
  signal reg_q960        : std_logic;
  signal reg_q960_in     : std_logic;
  		

  -- state q874
  signal reg_q874        : std_logic;
  signal reg_q874_in     : std_logic;
  		

  -- state q876
  signal reg_q876        : std_logic;
  signal reg_q876_in     : std_logic;
  		

  -- state q949
  signal reg_q949        : std_logic;
  signal reg_q949_in     : std_logic;
  		

  -- state q951
  signal reg_q951        : std_logic;
  signal reg_q951_in     : std_logic;
  		

  -- state q12
  signal reg_q12        : std_logic;
  signal reg_q12_in     : std_logic;
  		

  -- state q2409
  signal reg_q2409        : std_logic;
  signal reg_q2409_in     : std_logic;
  		

  -- state q882
  signal reg_q882        : std_logic;
  signal reg_q882_in     : std_logic;
  		

  -- state q2429
  signal reg_q2429        : std_logic;
  signal reg_q2429_in     : std_logic;
  		

  -- state q2526
  signal reg_q2526        : std_logic;
  signal reg_q2526_in     : std_logic;
  		

  -- state q2423
  signal reg_q2423        : std_logic;
  signal reg_q2423_in     : std_logic;
  		

  -- state q2425
  signal reg_q2425        : std_logic;
  signal reg_q2425_in     : std_logic;
  		

  -- state q2196
  signal reg_q2196        : std_logic;
  signal reg_q2196_in     : std_logic;
  		

  -- state q2198
  signal reg_q2198        : std_logic;
  signal reg_q2198_in     : std_logic;
  		

  -- state q854
  signal reg_q854        : std_logic;
  signal reg_q854_in     : std_logic;
  		

  -- state q612
  signal reg_q612        : std_logic;
  signal reg_q612_in     : std_logic;
  		

  -- state q614
  signal reg_q614        : std_logic;
  signal reg_q614_in     : std_logic;
  		

  -- state q34
  signal reg_q34        : std_logic;
  signal reg_q34_in     : std_logic;
  		

  -- state q36
  signal reg_q36        : std_logic;
  signal reg_q36_in     : std_logic;
  		

  -- state q2072
  signal reg_q2072        : std_logic;
  signal reg_q2072_in     : std_logic;
  		

  -- state q884
  signal reg_q884        : std_logic;
  signal reg_q884_in     : std_logic;
  		

  -- state q1207
  signal reg_q1207        : std_logic;
  signal reg_q1207_in     : std_logic;
  		

  -- state q1985
  signal reg_q1985        : std_logic;
  signal reg_q1985_in     : std_logic;
  		

  -- state q1401
  signal reg_q1401        : std_logic;
  signal reg_q1401_in     : std_logic;
  		

  -- state q1403
  signal reg_q1403        : std_logic;
  signal reg_q1403_in     : std_logic;
  		

  -- state q38
  signal reg_q38        : std_logic;
  signal reg_q38_in     : std_logic;
  		

  -- state q1916
  signal reg_q1916        : std_logic;
  signal reg_q1916_in     : std_logic;
  		

  -- state q1800
  signal reg_q1800        : std_logic;
  signal reg_q1800_in     : std_logic;
  		

  -- state q1226
  signal reg_q1226        : std_logic;
  signal reg_q1226_in     : std_logic;
  		

  -- state q2093
  signal reg_q2093        : std_logic;
  signal reg_q2093_in     : std_logic;
  		

  -- state q758
  signal reg_q758        : std_logic;
  signal reg_q758_in     : std_logic;
  		

  -- state q2182
  signal reg_q2182        : std_logic;
  signal reg_q2182_in     : std_logic;
  		

  -- state q2184
  signal reg_q2184        : std_logic;
  signal reg_q2184_in     : std_logic;
  		

  -- state q598
  signal reg_q598        : std_logic;
  signal reg_q598_in     : std_logic;
  		

  -- state q600
  signal reg_q600        : std_logic;
  signal reg_q600_in     : std_logic;
  		

  -- state q1981
  signal reg_q1981        : std_logic;
  signal reg_q1981_in     : std_logic;
  		

  -- state q2062
  signal reg_q2062        : std_logic;
  signal reg_q2062_in     : std_logic;
  		

  -- state q1393
  signal reg_q1393        : std_logic;
  signal reg_q1393_in     : std_logic;
  		

  -- state q474
  signal reg_q474        : std_logic;
  signal reg_q474_in     : std_logic;
  		

  -- state q476
  signal reg_q476        : std_logic;
  signal reg_q476_in     : std_logic;
  		

  -- state q2395
  signal reg_q2395        : std_logic;
  signal reg_q2395_in     : std_logic;
  		

  -- state q2397
  signal reg_q2397        : std_logic;
  signal reg_q2397_in     : std_logic;
  		

  -- state q1205
  signal reg_q1205        : std_logic;
  signal reg_q1205_in     : std_logic;
  		

  -- state q1924
  signal reg_q1924        : std_logic;
  signal reg_q1924_in     : std_logic;
  		

  -- state q2439
  signal reg_q2439        : std_logic;
  signal reg_q2439_in     : std_logic;
  		

  -- state q2441
  signal reg_q2441        : std_logic;
  signal reg_q2441_in     : std_logic;
  		

  -- state q630
  signal reg_q630        : std_logic;
  signal reg_q630_in     : std_logic;
  		

  -- state q1850
  signal reg_q1850        : std_logic;
  signal reg_q1850_in     : std_logic;
  		

  -- state q1888
  signal reg_q1888        : std_logic;
  signal reg_q1888_in     : std_logic;
  		

  -- state q1890
  signal reg_q1890        : std_logic;
  signal reg_q1890_in     : std_logic;
  		

  -- state q528
  signal reg_q528        : std_logic;
  signal reg_q528_in     : std_logic;
  		

  -- state q530
  signal reg_q530        : std_logic;
  signal reg_q530_in     : std_logic;
  		

  -- state q606
  signal reg_q606        : std_logic;
  signal reg_q606_in     : std_logic;
  		

  -- state q608
  signal reg_q608        : std_logic;
  signal reg_q608_in     : std_logic;
  		

  -- state q2431
  signal reg_q2431        : std_logic;
  signal reg_q2431_in     : std_logic;
  		

  -- state q2433
  signal reg_q2433        : std_logic;
  signal reg_q2433_in     : std_logic;
  		

  -- state q1987
  signal reg_q1987        : std_logic;
  signal reg_q1987_in     : std_logic;
  		

  -- state q1989
  signal reg_q1989        : std_logic;
  signal reg_q1989_in     : std_logic;
  		

  -- state q1832
  signal reg_q1832        : std_logic;
  signal reg_q1832_in     : std_logic;
  		

  -- state q1834
  signal reg_q1834        : std_logic;
  signal reg_q1834_in     : std_logic;
  		

  -- state q799
  signal reg_q799        : std_logic;
  signal reg_q799_in     : std_logic;
  		

  -- state q801
  signal reg_q801        : std_logic;
  signal reg_q801_in     : std_logic;
  		

  -- state q2415
  signal reg_q2415        : std_logic;
  signal reg_q2415_in     : std_logic;
  		

  -- state q1910
  signal reg_q1910        : std_logic;
  signal reg_q1910_in     : std_logic;
  		

  -- state q1912
  signal reg_q1912        : std_logic;
  signal reg_q1912_in     : std_logic;
  		

  -- state q578
  signal reg_q578        : std_logic;
  signal reg_q578_in     : std_logic;
  		

  -- state q580
  signal reg_q580        : std_logic;
  signal reg_q580_in     : std_logic;
  		

  -- state q1818
  signal reg_q1818        : std_logic;
  signal reg_q1818_in     : std_logic;
  		

  -- state q1820
  signal reg_q1820        : std_logic;
  signal reg_q1820_in     : std_logic;
  		

  -- state q1842
  signal reg_q1842        : std_logic;
  signal reg_q1842_in     : std_logic;
  		

  -- state q1844
  signal reg_q1844        : std_logic;
  signal reg_q1844_in     : std_logic;
  		

  -- state q18
  signal reg_q18        : std_logic;
  signal reg_q18_in     : std_logic;
  		

  -- state q1646
  signal reg_q1646        : std_logic;
  signal reg_q1646_in     : std_logic;
  		

  -- state q506
  signal reg_q506        : std_logic;
  signal reg_q506_in     : std_logic;
  		

  -- state q508
  signal reg_q508        : std_logic;
  signal reg_q508_in     : std_logic;
  		

  -- state q628
  signal reg_q628        : std_logic;
  signal reg_q628_in     : std_logic;
  		

  -- state q131
  signal reg_q131        : std_logic;
  signal reg_q131_in     : std_logic;
  		

  -- state q1381
  signal reg_q1381        : std_logic;
  signal reg_q1381_in     : std_logic;
  		

  -- state q1948
  signal reg_q1948        : std_logic;
  signal reg_q1948_in     : std_logic;
  		

  -- state q1950
  signal reg_q1950        : std_logic;
  signal reg_q1950_in     : std_logic;
  		

  -- state q1605
  signal reg_q1605        : std_logic;
  signal reg_q1605_in     : std_logic;
  		

  -- state q14
  signal reg_q14        : std_logic;
  signal reg_q14_in     : std_logic;
  		

  -- state q1979
  signal reg_q1979        : std_logic;
  signal reg_q1979_in     : std_logic;
  		

  -- state q795
  signal reg_q795        : std_logic;
  signal reg_q795_in     : std_logic;
  		

  -- state q797
  signal reg_q797        : std_logic;
  signal reg_q797_in     : std_logic;
  		

  -- state q510
  signal reg_q510        : std_logic;
  signal reg_q510_in     : std_logic;
  		

  -- state q1814
  signal reg_q1814        : std_logic;
  signal reg_q1814_in     : std_logic;
  		

  -- state q562
  signal reg_q562        : std_logic;
  signal reg_q562_in     : std_logic;
  		

  -- state q564
  signal reg_q564        : std_logic;
  signal reg_q564_in     : std_logic;
  		

  -- state q943
  signal reg_q943        : std_logic;
  signal reg_q943_in     : std_logic;
  		

  -- state q1942
  signal reg_q1942        : std_logic;
  signal reg_q1942_in     : std_logic;
  		

  -- state q1944
  signal reg_q1944        : std_logic;
  signal reg_q1944_in     : std_logic;
  		

  -- state q634
  signal reg_q634        : std_logic;
  signal reg_q634_in     : std_logic;
  		

  -- state q1213
  signal reg_q1213        : std_logic;
  signal reg_q1213_in     : std_logic;
  		

  -- state q1858
  signal reg_q1858        : std_logic;
  signal reg_q1858_in     : std_logic;
  		

  -- state q1860
  signal reg_q1860        : std_logic;
  signal reg_q1860_in     : std_logic;
  		

  -- state q1836
  signal reg_q1836        : std_logic;
  signal reg_q1836_in     : std_logic;
  		

  -- state q1525
  signal reg_q1525        : std_logic;
  signal reg_q1525_in     : std_logic;
  		

  -- state q878
  signal reg_q878        : std_logic;
  signal reg_q878_in     : std_logic;
  		

  -- state q1464
  signal reg_q1464        : std_logic;
  signal reg_q1464_in     : std_logic;
  		

  -- state q787
  signal reg_q787        : std_logic;
  signal reg_q787_in     : std_logic;
  		

  -- state q1862
  signal reg_q1862        : std_logic;
  signal reg_q1862_in     : std_logic;
  		

  -- state q1922
  signal reg_q1922        : std_logic;
  signal reg_q1922_in     : std_logic;
  		

  -- state q1550
  signal reg_q1550        : std_logic;
  signal reg_q1550_in     : std_logic;
  		

  -- state q1870
  signal reg_q1870        : std_logic;
  signal reg_q1870_in     : std_logic;
  		

  -- state q1991
  signal reg_q1991        : std_logic;
  signal reg_q1991_in     : std_logic;
  		

  -- state q1993
  signal reg_q1993        : std_logic;
  signal reg_q1993_in     : std_logic;
  		

  -- state q803
  signal reg_q803        : std_logic;
  signal reg_q803_in     : std_logic;
  		

  -- state q807
  signal reg_q807        : std_logic;
  signal reg_q807_in     : std_logic;
  		

  -- state q809
  signal reg_q809        : std_logic;
  signal reg_q809_in     : std_logic;
  		

  -- state q478
  signal reg_q478        : std_logic;
  signal reg_q478_in     : std_logic;
  		

  -- state q524
  signal reg_q524        : std_logic;
  signal reg_q524_in     : std_logic;
  		

  -- state q805
  signal reg_q805        : std_logic;
  signal reg_q805_in     : std_logic;
  		

  -- state q1219
  signal reg_q1219        : std_logic;
  signal reg_q1219_in     : std_logic;
  		

  -- state q1796
  signal reg_q1796        : std_logic;
  signal reg_q1796_in     : std_logic;
  		

  -- state q648
  signal reg_q648        : std_logic;
  signal reg_q648_in     : std_logic;
  		

  -- state q650
  signal reg_q650        : std_logic;
  signal reg_q650_in     : std_logic;
  		

  -- state q1822
  signal reg_q1822        : std_logic;
  signal reg_q1822_in     : std_logic;
  		

  -- state q1824
  signal reg_q1824        : std_logic;
  signal reg_q1824_in     : std_logic;
  		

  -- state q2192
  signal reg_q2192        : std_logic;
  signal reg_q2192_in     : std_logic;
  		

  -- state q1397
  signal reg_q1397        : std_logic;
  signal reg_q1397_in     : std_logic;
  		

  -- state q789
  signal reg_q789        : std_logic;
  signal reg_q789_in     : std_logic;
  		

  -- state q1830
  signal reg_q1830        : std_logic;
  signal reg_q1830_in     : std_logic;
  		

  -- state q1113
  signal reg_q1113        : std_logic;
  signal reg_q1113_in     : std_logic;
  		

  -- state q1983
  signal reg_q1983        : std_logic;
  signal reg_q1983_in     : std_logic;
  		

  -- state q1872
  signal reg_q1872        : std_logic;
  signal reg_q1872_in     : std_logic;
  		

  -- state q2186
  signal reg_q2186        : std_logic;
  signal reg_q2186_in     : std_logic;
  		

  -- state q2188
  signal reg_q2188        : std_logic;
  signal reg_q2188_in     : std_logic;
  		

  -- state q2162
  signal reg_q2162        : std_logic;
  signal reg_q2162_in     : std_logic;
  		

  -- state q1846
  signal reg_q1846        : std_logic;
  signal reg_q1846_in     : std_logic;
  		

  -- state q540
  signal reg_q540        : std_logic;
  signal reg_q540_in     : std_logic;
  		

  -- state q542
  signal reg_q542        : std_logic;
  signal reg_q542_in     : std_logic;
  		

  -- state q1798
  signal reg_q1798        : std_logic;
  signal reg_q1798_in     : std_logic;
  		

  -- state q1936
  signal reg_q1936        : std_logic;
  signal reg_q1936_in     : std_logic;
  		

  -- state q2200
  signal reg_q2200        : std_logic;
  signal reg_q2200_in     : std_logic;
  		

  -- state q941
  signal reg_q941        : std_logic;
  signal reg_q941_in     : std_logic;
  		

  -- state q572
  signal reg_q572        : std_logic;
  signal reg_q572_in     : std_logic;
  		

  -- state q574
  signal reg_q574        : std_logic;
  signal reg_q574_in     : std_logic;
  		

  -- state q862
  signal reg_q862        : std_logic;
  signal reg_q862_in     : std_logic;
  		

  -- state q1161
  signal reg_q1161        : std_logic;
  signal reg_q1161_in     : std_logic;
  		

  -- state q2524
  signal reg_q2524        : std_logic;
  signal reg_q2524_in     : std_logic;
  		

  -- state q638
  signal reg_q638        : std_logic;
  signal reg_q638_in     : std_logic;
  		

  -- state q640
  signal reg_q640        : std_logic;
  signal reg_q640_in     : std_logic;
  		

  -- state q594
  signal reg_q594        : std_logic;
  signal reg_q594_in     : std_logic;
  		

  -- state q32
  signal reg_q32        : std_logic;
  signal reg_q32_in     : std_logic;
  		

  -- state q872
  signal reg_q872        : std_logic;
  signal reg_q872_in     : std_logic;
  		

  -- state q2468
  signal reg_q2468        : std_logic;
  signal reg_q2468_in     : std_logic;
  		

  -- state q866
  signal reg_q866        : std_logic;
  signal reg_q866_in     : std_logic;
  		

  -- state q868
  signal reg_q868        : std_logic;
  signal reg_q868_in     : std_logic;
  		

  -- state q870
  signal reg_q870        : std_logic;
  signal reg_q870_in     : std_logic;
  		

  -- state q1399
  signal reg_q1399        : std_logic;
  signal reg_q1399_in     : std_logic;
  		

  -- state q1928
  signal reg_q1928        : std_logic;
  signal reg_q1928_in     : std_logic;
  		

  -- state q642
  signal reg_q642        : std_logic;
  signal reg_q642_in     : std_logic;
  		

  -- state q644
  signal reg_q644        : std_logic;
  signal reg_q644_in     : std_logic;
  		

  -- state q2487
  signal reg_q2487        : std_logic;
  signal reg_q2487_in     : std_logic;
  		

  -- state q2489
  signal reg_q2489        : std_logic;
  signal reg_q2489_in     : std_logic;
  		

  -- state q636
  signal reg_q636        : std_logic;
  signal reg_q636_in     : std_logic;
  		

  -- state q552
  signal reg_q552        : std_logic;
  signal reg_q552_in     : std_logic;
  		

  -- state q554
  signal reg_q554        : std_logic;
  signal reg_q554_in     : std_logic;
  		

  -- state q1365
  signal reg_q1365        : std_logic;
  signal reg_q1365_in     : std_logic;
  		

  -- state q1367
  signal reg_q1367        : std_logic;
  signal reg_q1367_in     : std_logic;
  		

  -- state q1812
  signal reg_q1812        : std_logic;
  signal reg_q1812_in     : std_logic;
  		

  -- state q1371
  signal reg_q1371        : std_logic;
  signal reg_q1371_in     : std_logic;
  		

  -- state q2399
  signal reg_q2399        : std_logic;
  signal reg_q2399_in     : std_logic;
  		

  -- state q2401
  signal reg_q2401        : std_logic;
  signal reg_q2401_in     : std_logic;
  		

  -- state q1908
  signal reg_q1908        : std_logic;
  signal reg_q1908_in     : std_logic;
  		

  -- state q584
  signal reg_q584        : std_logic;
  signal reg_q584_in     : std_logic;
  		

  -- state q586
  signal reg_q586        : std_logic;
  signal reg_q586_in     : std_logic;
  		

  -- state q576
  signal reg_q576        : std_logic;
  signal reg_q576_in     : std_logic;
  		

  -- state q20
  signal reg_q20        : std_logic;
  signal reg_q20_in     : std_logic;
  		

  -- state q2435
  signal reg_q2435        : std_logic;
  signal reg_q2435_in     : std_logic;
  		

  -- state q2437
  signal reg_q2437        : std_logic;
  signal reg_q2437_in     : std_logic;
  		

  -- state q2413
  signal reg_q2413        : std_logic;
  signal reg_q2413_in     : std_logic;
  		

  -- state q560
  signal reg_q560        : std_logic;
  signal reg_q560_in     : std_logic;
  		

  -- state q1804
  signal reg_q1804        : std_logic;
  signal reg_q1804_in     : std_logic;
  		

  -- state q1806
  signal reg_q1806        : std_logic;
  signal reg_q1806_in     : std_logic;
  		

  -- state q472
  signal reg_q472        : std_logic;
  signal reg_q472_in     : std_logic;
  		

  -- state q546
  signal reg_q546        : std_logic;
  signal reg_q546_in     : std_logic;
  		

  -- state q548
  signal reg_q548        : std_logic;
  signal reg_q548_in     : std_logic;
  		

  -- state q2493
  signal reg_q2493        : std_logic;
  signal reg_q2493_in     : std_logic;
  		

  -- state q582
  signal reg_q582        : std_logic;
  signal reg_q582_in     : std_logic;
  		

  -- state q492
  signal reg_q492        : std_logic;
  signal reg_q492_in     : std_logic;
  		

  -- state q494
  signal reg_q494        : std_logic;
  signal reg_q494_in     : std_logic;
  		

  -- state q602
  signal reg_q602        : std_logic;
  signal reg_q602_in     : std_logic;
  		

  -- state q2082
  signal reg_q2082        : std_logic;
  signal reg_q2082_in     : std_logic;
  		

  -- state q2084
  signal reg_q2084        : std_logic;
  signal reg_q2084_in     : std_logic;
  		

  -- state q2190
  signal reg_q2190        : std_logic;
  signal reg_q2190_in     : std_logic;
  		

  -- state q1838
  signal reg_q1838        : std_logic;
  signal reg_q1838_in     : std_logic;
  		

  -- state q1898
  signal reg_q1898        : std_logic;
  signal reg_q1898_in     : std_logic;
  		

  -- state q1900
  signal reg_q1900        : std_logic;
  signal reg_q1900_in     : std_logic;
  		

  -- state q8
  signal reg_q8        : std_logic;
  signal reg_q8_in     : std_logic;
  		

  -- state q496
  signal reg_q496        : std_logic;
  signal reg_q496_in     : std_logic;
  		

  -- state q498
  signal reg_q498        : std_logic;
  signal reg_q498_in     : std_logic;
  		

  -- state q462
  signal reg_q462        : std_logic;
  signal reg_q462_in     : std_logic;
  		

  -- state q464
  signal reg_q464        : std_logic;
  signal reg_q464_in     : std_logic;
  		

  -- state q568
  signal reg_q568        : std_logic;
  signal reg_q568_in     : std_logic;
  		

  -- state q1930
  signal reg_q1930        : std_logic;
  signal reg_q1930_in     : std_logic;
  		

  -- state q1932
  signal reg_q1932        : std_logic;
  signal reg_q1932_in     : std_logic;
  		

  -- state q512
  signal reg_q512        : std_logic;
  signal reg_q512_in     : std_logic;
  		

  -- state q1914
  signal reg_q1914        : std_logic;
  signal reg_q1914_in     : std_logic;
  		

  -- state q1379
  signal reg_q1379        : std_logic;
  signal reg_q1379_in     : std_logic;
  		

  -- state q1199
  signal reg_q1199        : std_logic;
  signal reg_q1199_in     : std_logic;
  		

  -- state q544
  signal reg_q544        : std_logic;
  signal reg_q544_in     : std_logic;
  		

  -- state q470
  signal reg_q470        : std_logic;
  signal reg_q470_in     : std_logic;
  		

  -- state q2508
  signal reg_q2508        : std_logic;
  signal reg_q2508_in     : std_logic;
  		

  -- state q480
  signal reg_q480        : std_logic;
  signal reg_q480_in     : std_logic;
  		

  -- state q482
  signal reg_q482        : std_logic;
  signal reg_q482_in     : std_logic;
  		

  -- state q500
  signal reg_q500        : std_logic;
  signal reg_q500_in     : std_logic;
  		

  -- state q1894
  signal reg_q1894        : std_logic;
  signal reg_q1894_in     : std_logic;
  		

  -- state q1896
  signal reg_q1896        : std_logic;
  signal reg_q1896_in     : std_logic;
  		

  -- state q820
  signal reg_q820        : std_logic;
  signal reg_q820_in     : std_logic;
  		

  -- state q905
  signal reg_q905        : std_logic;
  signal reg_q905_in     : std_logic;
  		

  -- state q24
  signal reg_q24        : std_logic;
  signal reg_q24_in     : std_logic;
  		

  -- state q1856
  signal reg_q1856        : std_logic;
  signal reg_q1856_in     : std_logic;
  		

  -- state q1203
  signal reg_q1203        : std_logic;
  signal reg_q1203_in     : std_logic;
  		

  -- state q1934
  signal reg_q1934        : std_logic;
  signal reg_q1934_in     : std_logic;
  		

  -- state q736
  signal reg_q736        : std_logic;
  signal reg_q736_in     : std_logic;
  		

  -- state q484
  signal reg_q484        : std_logic;
  signal reg_q484_in     : std_logic;
  		

  -- state q486
  signal reg_q486        : std_logic;
  signal reg_q486_in     : std_logic;
  		

  -- state q550
  signal reg_q550        : std_logic;
  signal reg_q550_in     : std_logic;
  		

  -- state q2086
  signal reg_q2086        : std_logic;
  signal reg_q2086_in     : std_logic;
  		

  -- state q2088
  signal reg_q2088        : std_logic;
  signal reg_q2088_in     : std_logic;
  		

  -- state q514
  signal reg_q514        : std_logic;
  signal reg_q514_in     : std_logic;
  		

  -- state q468
  signal reg_q468        : std_logic;
  signal reg_q468_in     : std_logic;
  		

  -- state q1902
  signal reg_q1902        : std_logic;
  signal reg_q1902_in     : std_logic;
  		

  -- state q28
  signal reg_q28        : std_logic;
  signal reg_q28_in     : std_logic;
  		

  -- state q30
  signal reg_q30        : std_logic;
  signal reg_q30_in     : std_logic;
  		

  -- state q917
  signal reg_q917        : std_logic;
  signal reg_q917_in     : std_logic;
  		

  -- state q2443
  signal reg_q2443        : std_logic;
  signal reg_q2443_in     : std_logic;
  		

  -- state q1808
  signal reg_q1808        : std_logic;
  signal reg_q1808_in     : std_logic;
  		

  -- state q1810
  signal reg_q1810        : std_logic;
  signal reg_q1810_in     : std_logic;
  		

  -- state q1369
  signal reg_q1369        : std_logic;
  signal reg_q1369_in     : std_logic;
  		

  -- state q588
  signal reg_q588        : std_logic;
  signal reg_q588_in     : std_logic;
  		

  -- state q1892
  signal reg_q1892        : std_logic;
  signal reg_q1892_in     : std_logic;
  		

  -- state q538
  signal reg_q538        : std_logic;
  signal reg_q538_in     : std_logic;
  		

  -- state q1391
  signal reg_q1391        : std_logic;
  signal reg_q1391_in     : std_logic;
  		

  -- state q502
  signal reg_q502        : std_logic;
  signal reg_q502_in     : std_logic;
  		

  -- state q504
  signal reg_q504        : std_logic;
  signal reg_q504_in     : std_logic;
  		

  -- state q466
  signal reg_q466        : std_logic;
  signal reg_q466_in     : std_logic;
  		

  -- state q2463
  signal reg_q2463        : std_logic;
  signal reg_q2463_in     : std_logic;
  		

  -- state q2391
  signal reg_q2391        : std_logic;
  signal reg_q2391_in     : std_logic;
  		

  -- state q2325
  signal reg_q2325        : std_logic;
  signal reg_q2325_in     : std_logic;
  		

  -- state q26
  signal reg_q26        : std_logic;
  signal reg_q26_in     : std_logic;
  		

  -- state q903
  signal reg_q903        : std_logic;
  signal reg_q903_in     : std_logic;
  		

  -- state q518
  signal reg_q518        : std_logic;
  signal reg_q518_in     : std_logic;
  		

  -- state q1840
  signal reg_q1840        : std_logic;
  signal reg_q1840_in     : std_logic;
  		

  -- state q624
  signal reg_q624        : std_logic;
  signal reg_q624_in     : std_logic;
  		

  -- state q626
  signal reg_q626        : std_logic;
  signal reg_q626_in     : std_logic;
  		

  -- state q516
  signal reg_q516        : std_logic;
  signal reg_q516_in     : std_logic;
  		

  -- state q1946
  signal reg_q1946        : std_logic;
  signal reg_q1946_in     : std_logic;
  		

  -- state q1864
  signal reg_q1864        : std_logic;
  signal reg_q1864_in     : std_logic;
  		

  -- state q1940
  signal reg_q1940        : std_logic;
  signal reg_q1940_in     : std_logic;
  		

  -- state q42
  signal reg_q42        : std_logic;
  signal reg_q42_in     : std_logic;
  		

  -- state q44
  signal reg_q44        : std_logic;
  signal reg_q44_in     : std_logic;
  		

  -- state q2202
  signal reg_q2202        : std_logic;
  signal reg_q2202_in     : std_logic;
  		

  -- state q2520
  signal reg_q2520        : std_logic;
  signal reg_q2520_in     : std_logic;
  		

  -- state q860
  signal reg_q860        : std_logic;
  signal reg_q860_in     : std_logic;
  		

  -- state q1031
  signal reg_q1031        : std_logic;
  signal reg_q1031_in     : std_logic;
  		

  -- state q2393
  signal reg_q2393        : std_logic;
  signal reg_q2393_in     : std_logic;
  		

  -- state q2204
  signal reg_q2204        : std_logic;
  signal reg_q2204_in     : std_logic;
  		

  -- state q2206
  signal reg_q2206        : std_logic;
  signal reg_q2206_in     : std_logic;
  		

  -- state q646
  signal reg_q646        : std_logic;
  signal reg_q646_in     : std_logic;
  		

  -- state q2403
  signal reg_q2403        : std_logic;
  signal reg_q2403_in     : std_logic;
  		

  -- state q1952
  signal reg_q1952        : std_logic;
  signal reg_q1952_in     : std_logic;
  		

  -- state q1405
  signal reg_q1405        : std_logic;
  signal reg_q1405_in     : std_logic;
  		

  -- state q1407
  signal reg_q1407        : std_logic;
  signal reg_q1407_in     : std_logic;
  		

  -- state q622
  signal reg_q622        : std_logic;
  signal reg_q622_in     : std_logic;
  		

  -- state q488
  signal reg_q488        : std_logic;
  signal reg_q488_in     : std_logic;
  		

  -- state q490
  signal reg_q490        : std_logic;
  signal reg_q490_in     : std_logic;
  		

  -- state q40
  signal reg_q40        : std_logic;
  signal reg_q40_in     : std_logic;
  		

  -- state q654
  signal reg_q654        : std_logic;
  signal reg_q654_in     : std_logic;
  		

  -- state q656
  signal reg_q656        : std_logic;
  signal reg_q656_in     : std_logic;
  		

  -- state q570
  signal reg_q570        : std_logic;
  signal reg_q570_in     : std_logic;
  		

  -- state q822
  signal reg_q822        : std_logic;
  signal reg_q822_in     : std_logic;
  		

  -- state q1363
  signal reg_q1363        : std_logic;
  signal reg_q1363_in     : std_logic;
  		

  -- state q2522
  signal reg_q2522        : std_logic;
  signal reg_q2522_in     : std_logic;
  		

  -- state q652
  signal reg_q652        : std_logic;
  signal reg_q652_in     : std_logic;
  		

  -- state q1413
  signal reg_q1413        : std_logic;
  signal reg_q1413_in     : std_logic;
  		

  -- state q610
  signal reg_q610        : std_logic;
  signal reg_q610_in     : std_logic;
  		

  -- state q536
  signal reg_q536        : std_logic;
  signal reg_q536_in     : std_logic;
  		

  -- state q2056
  signal reg_q2056        : std_logic;
  signal reg_q2056_in     : std_logic;
  		

  -- state q2058
  signal reg_q2058        : std_logic;
  signal reg_q2058_in     : std_logic;
  		

  -- state q660
  signal reg_q660        : std_logic;
  signal reg_q660_in     : std_logic;
  		

  -- state q662
  signal reg_q662        : std_logic;
  signal reg_q662_in     : std_logic;
  		

  -- state q2060
  signal reg_q2060        : std_logic;
  signal reg_q2060_in     : std_logic;
  		

  -- state q658
  signal reg_q658        : std_logic;
  signal reg_q658_in     : std_logic;
  		

  -- state q2076
  signal reg_q2076        : std_logic;
  signal reg_q2076_in     : std_logic;
  		
  signal reg_fullgraph7       : std_logic_vector(8 downto 0);
  signal reg_fullgraph7_in    : std_logic_vector(8 downto 0);
  signal reg_fullgraph7_init  : std_logic_vector(8 downto 0);
  signal reg_fullgraph7_sel   : std_logic_vector(511 downto 0); 	
  -- end section fullgraph7
  --#################################################			
		

  -- state q0
  signal reg_q0        : std_logic;
  signal reg_q0_in     : std_logic;
  signal reg_q0_init   : std_logic;
		

  -- state q850
  signal reg_q850        : std_logic;
  signal reg_q850_in     : std_logic;
  signal reg_q850_init   : std_logic;
		
--#################################################
-- start section fullgraph: 10

  -- state q2615
  signal reg_q2615        : std_logic;
  signal reg_q2615_in     : std_logic;
  		

  -- state q1112
  signal reg_q1112        : std_logic;
  signal reg_q1112_in     : std_logic;
  		

  -- state q953
  signal reg_q953        : std_logic;
  signal reg_q953_in     : std_logic;
  		

  -- state q2504
  signal reg_q2504        : std_logic;
  signal reg_q2504_in     : std_logic;
  		

  -- state q2506
  signal reg_q2506        : std_logic;
  signal reg_q2506_in     : std_logic;
  		

  -- state q2510
  signal reg_q2510        : std_logic;
  signal reg_q2510_in     : std_logic;
  		

  -- state q2491
  signal reg_q2491        : std_logic;
  signal reg_q2491_in     : std_logic;
  		

  -- state q2485
  signal reg_q2485        : std_logic;
  signal reg_q2485_in     : std_logic;
  		
  signal reg_fullgraph10       : std_logic_vector(3 downto 0);
  signal reg_fullgraph10_in    : std_logic_vector(3 downto 0);
  signal reg_fullgraph10_init  : std_logic_vector(3 downto 0);
  signal reg_fullgraph10_sel   : std_logic_vector(15 downto 0); 	
  -- end section fullgraph10
  --#################################################			
		

  -- state q1359
  signal reg_q1359        : std_logic;
  signal reg_q1359_in     : std_logic;
  signal reg_q1359_init   : std_logic;
		

  -- state q2618
  signal reg_q2618        : std_logic;
  signal reg_q2618_in     : std_logic;
  signal reg_q2618_init   : std_logic;
		

  -- state q1742
  signal reg_q1742        : std_logic;
  signal reg_q1742_in     : std_logic;
  signal reg_q1742_init   : std_logic;
		

  -- state q2383
  signal reg_q2383        : std_logic;
  signal reg_q2383_in     : std_logic;
  signal reg_q2383_init   : std_logic;
		

  -- state q2124
  signal reg_q2124        : std_logic;
  signal reg_q2124_in     : std_logic;
  signal reg_q2124_init   : std_logic;
		

  -- state q1111
  signal reg_q1111        : std_logic;
  signal reg_q1111_in     : std_logic;
  signal reg_q1111_init   : std_logic;
		

  -- state q556
  signal reg_q556        : std_logic;
  signal reg_q556_in     : std_logic;
  signal reg_q556_init   : std_logic;
		

  -- state q2091
  signal reg_q2091        : std_logic;
  signal reg_q2091_in     : std_logic;
  signal reg_q2091_init   : std_logic;
		

  -- state q452
  signal reg_q452        : std_logic;
  signal reg_q452_in     : std_logic;
  signal reg_q452_init   : std_logic;
		

  -- state q1195
  signal reg_q1195        : std_logic;
  signal reg_q1195_in     : std_logic;
  signal reg_q1195_init   : std_logic;
		

  -- state q1644
  signal reg_q1644        : std_logic;
  signal reg_q1644_in     : std_logic;
  signal reg_q1644_init   : std_logic;
		

  -- state q1603
  signal reg_q1603        : std_logic;
  signal reg_q1603_in     : std_logic;
  signal reg_q1603_init   : std_logic;
		

  -- state q2323
  signal reg_q2323        : std_logic;
  signal reg_q2323_in     : std_logic;
  signal reg_q2323_init   : std_logic;
		

  -- state q1013
  signal reg_q1013        : std_logic;
  signal reg_q1013_in     : std_logic;
  signal reg_q1013_init   : std_logic;
		

  -- state q46
  signal reg_q46        : std_logic;
  signal reg_q46_in     : std_logic;
  signal reg_q46_init   : std_logic;
		

  -- state q1050
  signal reg_q1050        : std_logic;
  signal reg_q1050_in     : std_logic;
  signal reg_q1050_init   : std_logic;
		

  -- state q680
  signal reg_q680        : std_logic;
  signal reg_q680_in     : std_logic;
  signal reg_q680_init   : std_logic;
		

  -- state q1521
  signal reg_q1521        : std_logic;
  signal reg_q1521_in     : std_logic;
  signal reg_q1521_init   : std_logic;
		

  -- state q1884
  signal reg_q1884        : std_logic;
  signal reg_q1884_in     : std_logic;
  signal reg_q1884_init   : std_logic;
		

  -- state q1955
  signal reg_q1955        : std_logic;
  signal reg_q1955_in     : std_logic;
  signal reg_q1955_init   : std_logic;
		

  -- state q262
  signal reg_q262        : std_logic;
  signal reg_q262_in     : std_logic;
  signal reg_q262_init   : std_logic;
		

  -- state q958
  signal reg_q958        : std_logic;
  signal reg_q958_in     : std_logic;
  signal reg_q958_init   : std_logic;
		

  -- state q816
  signal reg_q816        : std_logic;
  signal reg_q816_in     : std_logic;
  signal reg_q816_init   : std_logic;
		

  -- state q1224
  signal reg_q1224        : std_logic;
  signal reg_q1224_in     : std_logic;
  signal reg_q1224_init   : std_logic;
		

  -- state q896
  signal reg_q896        : std_logic;
  signal reg_q896_in     : std_logic;
  signal reg_q896_init   : std_logic;
		

  -- state q2000
  signal reg_q2000        : std_logic;
  signal reg_q2000_in     : std_logic;
  signal reg_q2000_init   : std_logic;
		

  -- state q2533
  signal reg_q2533        : std_logic;
  signal reg_q2533_in     : std_logic;
  signal reg_q2533_init   : std_logic;
		

  -- state q303
  signal reg_q303        : std_logic;
  signal reg_q303_in     : std_logic;
  signal reg_q303_init   : std_logic;
		

  -- state q665
  signal reg_q665        : std_logic;
  signal reg_q665_in     : std_logic;
  signal reg_q665_init   : std_logic;
		

  -- state q703
  signal reg_q703        : std_logic;
  signal reg_q703_in     : std_logic;
  signal reg_q703_init   : std_logic;
		

  -- state q414
  signal reg_q414        : std_logic;
  signal reg_q414_in     : std_logic;
  signal reg_q414_init   : std_logic;
		

  -- state q2252
  signal reg_q2252        : std_logic;
  signal reg_q2252_in     : std_logic;
  signal reg_q2252_init   : std_logic;
		
--#################################################
-- start section fullgraph: 43

  -- state q1772
  signal reg_q1772        : std_logic;
  signal reg_q1772_in     : std_logic;
  		

  -- state q618
  signal reg_q618        : std_logic;
  signal reg_q618_in     : std_logic;
  		

  -- state q48
  signal reg_q48        : std_logic;
  signal reg_q48_in     : std_logic;
  		

  -- state q227
  signal reg_q227        : std_logic;
  signal reg_q227_in     : std_logic;
  		

  -- state q229
  signal reg_q229        : std_logic;
  signal reg_q229_in     : std_logic;
  		

  -- state q233
  signal reg_q233        : std_logic;
  signal reg_q233_in     : std_logic;
  		

  -- state q182
  signal reg_q182        : std_logic;
  signal reg_q182_in     : std_logic;
  		

  -- state q184
  signal reg_q184        : std_logic;
  signal reg_q184_in     : std_logic;
  		

  -- state q231
  signal reg_q231        : std_logic;
  signal reg_q231_in     : std_logic;
  		

  -- state q1790
  signal reg_q1790        : std_logic;
  signal reg_q1790_in     : std_logic;
  		

  -- state q1385
  signal reg_q1385        : std_logic;
  signal reg_q1385_in     : std_logic;
  		

  -- state q1211
  signal reg_q1211        : std_logic;
  signal reg_q1211_in     : std_logic;
  		

  -- state q2451
  signal reg_q2451        : std_logic;
  signal reg_q2451_in     : std_logic;
  		

  -- state q2453
  signal reg_q2453        : std_logic;
  signal reg_q2453_in     : std_logic;
  		

  -- state q1015
  signal reg_q1015        : std_logic;
  signal reg_q1015_in     : std_logic;
  		

  -- state q2128
  signal reg_q2128        : std_logic;
  signal reg_q2128_in     : std_logic;
  		

  -- state q2213
  signal reg_q2213        : std_logic;
  signal reg_q2213_in     : std_logic;
  		

  -- state q264
  signal reg_q264        : std_logic;
  signal reg_q264_in     : std_logic;
  		

  -- state q705
  signal reg_q705        : std_logic;
  signal reg_q705_in     : std_logic;
  		

  -- state q2132
  signal reg_q2132        : std_logic;
  signal reg_q2132_in     : std_logic;
  		

  -- state q1957
  signal reg_q1957        : std_logic;
  signal reg_q1957_in     : std_logic;
  		

  -- state q2455
  signal reg_q2455        : std_logic;
  signal reg_q2455_in     : std_logic;
  		

  -- state q50
  signal reg_q50        : std_logic;
  signal reg_q50_in     : std_logic;
  		

  -- state q52
  signal reg_q52        : std_logic;
  signal reg_q52_in     : std_logic;
  		

  -- state q186
  signal reg_q186        : std_logic;
  signal reg_q186_in     : std_logic;
  		

  -- state q1906
  signal reg_q1906        : std_logic;
  signal reg_q1906_in     : std_logic;
  		

  -- state q188
  signal reg_q188        : std_logic;
  signal reg_q188_in     : std_logic;
  		

  -- state q190
  signal reg_q190        : std_logic;
  signal reg_q190_in     : std_logic;
  		

  -- state q2068
  signal reg_q2068        : std_logic;
  signal reg_q2068_in     : std_logic;
  		

  -- state q2449
  signal reg_q2449        : std_logic;
  signal reg_q2449_in     : std_logic;
  		

  -- state q1377
  signal reg_q1377        : std_logic;
  signal reg_q1377_in     : std_logic;
  		

  -- state q180
  signal reg_q180        : std_logic;
  signal reg_q180_in     : std_logic;
  		

  -- state q416
  signal reg_q416        : std_logic;
  signal reg_q416_in     : std_logic;
  		

  -- state q1694
  signal reg_q1694        : std_logic;
  signal reg_q1694_in     : std_logic;
  		

  -- state q718
  signal reg_q718        : std_logic;
  signal reg_q718_in     : std_logic;
  		

  -- state q2461
  signal reg_q2461        : std_logic;
  signal reg_q2461_in     : std_logic;
  		

  -- state q2070
  signal reg_q2070        : std_logic;
  signal reg_q2070_in     : std_logic;
  		

  -- state q2457
  signal reg_q2457        : std_logic;
  signal reg_q2457_in     : std_logic;
  		

  -- state q2459
  signal reg_q2459        : std_logic;
  signal reg_q2459_in     : std_logic;
  		

  -- state q2150
  signal reg_q2150        : std_logic;
  signal reg_q2150_in     : std_logic;
  		

  -- state q1375
  signal reg_q1375        : std_logic;
  signal reg_q1375_in     : std_logic;
  		

  -- state q97
  signal reg_q97        : std_logic;
  signal reg_q97_in     : std_logic;
  		

  -- state q2465
  signal reg_q2465        : std_logic;
  signal reg_q2465_in     : std_logic;
  		
  signal reg_fullgraph43       : std_logic_vector(5 downto 0);
  signal reg_fullgraph43_in    : std_logic_vector(5 downto 0);
  signal reg_fullgraph43_init  : std_logic_vector(5 downto 0);
  signal reg_fullgraph43_sel   : std_logic_vector(63 downto 0); 	
  -- end section fullgraph43
  --#################################################			
		

  -- state q2211
  signal reg_q2211        : std_logic;
  signal reg_q2211_in     : std_logic;
  signal reg_q2211_init   : std_logic;
		
--#################################################
-- start section fullgraph: 45

  -- state q813
  signal reg_q813        : std_logic;
  signal reg_q813_in     : std_logic;
  		

  -- state q1298
  signal reg_q1298        : std_logic;
  signal reg_q1298_in     : std_logic;
  		

  -- state q901
  signal reg_q901        : std_logic;
  signal reg_q901_in     : std_logic;
  		

  -- state q781
  signal reg_q781        : std_logic;
  signal reg_q781_in     : std_logic;
  		

  -- state q1052
  signal reg_q1052        : std_logic;
  signal reg_q1052_in     : std_logic;
  		

  -- state q2126
  signal reg_q2126        : std_logic;
  signal reg_q2126_in     : std_logic;
  		

  -- state q1523
  signal reg_q1523        : std_logic;
  signal reg_q1523_in     : std_logic;
  		

  -- state q2587
  signal reg_q2587        : std_logic;
  signal reg_q2587_in     : std_logic;
  		

  -- state q1995
  signal reg_q1995        : std_logic;
  signal reg_q1995_in     : std_logic;
  		
  signal reg_fullgraph45       : std_logic_vector(3 downto 0);
  signal reg_fullgraph45_in    : std_logic_vector(3 downto 0);
  signal reg_fullgraph45_init  : std_logic_vector(3 downto 0);
  signal reg_fullgraph45_sel   : std_logic_vector(15 downto 0); 	
  -- end section fullgraph45
  --#################################################			
		

  -- state q714
  signal reg_q714        : std_logic;
  signal reg_q714_in     : std_logic;
  signal reg_q714_init   : std_logic;
		

  -- state q1544
  signal reg_q1544        : std_logic;
  signal reg_q1544_in     : std_logic;
  signal reg_q1544_init   : std_logic;
		

  -- state q2208
  signal reg_q2208        : std_logic;
  signal reg_q2208_in     : std_logic;
  signal reg_q2208_init   : std_logic;
		
--#################################################
-- start section fullgraph: 49

  -- state q1209
  signal reg_q1209        : std_logic;
  signal reg_q1209_in     : std_logic;
  		

  -- state q832
  signal reg_q832        : std_logic;
  signal reg_q832_in     : std_logic;
  		

  -- state q1868
  signal reg_q1868        : std_logic;
  signal reg_q1868_in     : std_logic;
  		

  -- state q842
  signal reg_q842        : std_logic;
  signal reg_q842_in     : std_logic;
  		

  -- state q1918
  signal reg_q1918        : std_logic;
  signal reg_q1918_in     : std_logic;
  		

  -- state q2066
  signal reg_q2066        : std_logic;
  signal reg_q2066_in     : std_logic;
  		

  -- state q10
  signal reg_q10        : std_logic;
  signal reg_q10_in     : std_logic;
  		

  -- state q2411
  signal reg_q2411        : std_logic;
  signal reg_q2411_in     : std_logic;
  		

  -- state q880
  signal reg_q880        : std_logic;
  signal reg_q880_in     : std_logic;
  		

  -- state q2417
  signal reg_q2417        : std_logic;
  signal reg_q2417_in     : std_logic;
  		

  -- state q2427
  signal reg_q2427        : std_logic;
  signal reg_q2427_in     : std_logic;
  		

  -- state q1373
  signal reg_q1373        : std_logic;
  signal reg_q1373_in     : std_logic;
  		

  -- state q2074
  signal reg_q2074        : std_logic;
  signal reg_q2074_in     : std_logic;
  		

  -- state q2194
  signal reg_q2194        : std_logic;
  signal reg_q2194_in     : std_logic;
  		

  -- state q1802
  signal reg_q1802        : std_logic;
  signal reg_q1802_in     : std_logic;
  		

  -- state q1395
  signal reg_q1395        : std_logic;
  signal reg_q1395_in     : std_logic;
  		

  -- state q1926
  signal reg_q1926        : std_logic;
  signal reg_q1926_in     : std_logic;
  		

  -- state q632
  signal reg_q632        : std_logic;
  signal reg_q632_in     : std_logic;
  		

  -- state q887
  signal reg_q887        : std_logic;
  signal reg_q887_in     : std_logic;
  		

  -- state q1848
  signal reg_q1848        : std_logic;
  signal reg_q1848_in     : std_logic;
  		

  -- state q2176
  signal reg_q2176        : std_logic;
  signal reg_q2176_in     : std_logic;
  		

  -- state q16
  signal reg_q16        : std_logic;
  signal reg_q16_in     : std_logic;
  		

  -- state q1361
  signal reg_q1361        : std_logic;
  signal reg_q1361_in     : std_logic;
  		

  -- state q1938
  signal reg_q1938        : std_logic;
  signal reg_q1938_in     : std_logic;
  		

  -- state q1383
  signal reg_q1383        : std_logic;
  signal reg_q1383_in     : std_logic;
  		

  -- state q1880
  signal reg_q1880        : std_logic;
  signal reg_q1880_in     : std_logic;
  		

  -- state q1886
  signal reg_q1886        : std_logic;
  signal reg_q1886_in     : std_logic;
  		

  -- state q864
  signal reg_q864        : std_logic;
  signal reg_q864_in     : std_logic;
  		

  -- state q1816
  signal reg_q1816        : std_logic;
  signal reg_q1816_in     : std_logic;
  		

  -- state q893
  signal reg_q893        : std_logic;
  signal reg_q893_in     : std_logic;
  		

  -- state q604
  signal reg_q604        : std_logic;
  signal reg_q604_in     : std_logic;
  		

  -- state q1221
  signal reg_q1221        : std_logic;
  signal reg_q1221_in     : std_logic;
  		

  -- state q2385
  signal reg_q2385        : std_logic;
  signal reg_q2385_in     : std_logic;
  		

  -- state q596
  signal reg_q596        : std_logic;
  signal reg_q596_in     : std_logic;
  		

  -- state q716
  signal reg_q716        : std_logic;
  signal reg_q716_in     : std_logic;
  		

  -- state q1904
  signal reg_q1904        : std_logic;
  signal reg_q1904_in     : std_logic;
  		

  -- state q458
  signal reg_q458        : std_logic;
  signal reg_q458_in     : std_logic;
  		

  -- state q460
  signal reg_q460        : std_logic;
  signal reg_q460_in     : std_logic;
  		

  -- state q22
  signal reg_q22        : std_logic;
  signal reg_q22_in     : std_logic;
  		

  -- state q558
  signal reg_q558        : std_logic;
  signal reg_q558_in     : std_logic;
  		

  -- state q811
  signal reg_q811        : std_logic;
  signal reg_q811_in     : std_logic;
  		

  -- state q566
  signal reg_q566        : std_logic;
  signal reg_q566_in     : std_logic;
  		

  -- state q1201
  signal reg_q1201        : std_logic;
  signal reg_q1201_in     : std_logic;
  		

  -- state q886
  signal reg_q886        : std_logic;
  signal reg_q886_in     : std_logic;
  		

  -- state q2054
  signal reg_q2054        : std_logic;
  signal reg_q2054_in     : std_logic;
  		

  -- state q93
  signal reg_q93        : std_logic;
  signal reg_q93_in     : std_logic;
  		

  -- state q456
  signal reg_q456        : std_logic;
  signal reg_q456_in     : std_logic;
  		

  -- state q852
  signal reg_q852        : std_logic;
  signal reg_q852_in     : std_logic;
  		

  -- state q95
  signal reg_q95        : std_logic;
  signal reg_q95_in     : std_logic;
  		
  signal reg_fullgraph49       : std_logic_vector(5 downto 0);
  signal reg_fullgraph49_in    : std_logic_vector(5 downto 0);
  signal reg_fullgraph49_init  : std_logic_vector(5 downto 0);
  signal reg_fullgraph49_sel   : std_logic_vector(63 downto 0); 	
  -- end section fullgraph49
  --#################################################			
		

  -- state q2518
  signal reg_q2518        : std_logic;
  signal reg_q2518_in     : std_logic;
  signal reg_q2518_init   : std_logic;
		

  -- state q2052
  signal reg_q2052        : std_logic;
  signal reg_q2052_in     : std_logic;
  signal reg_q2052_init   : std_logic;
		

  -- state q779
  signal reg_q779        : std_logic;
  signal reg_q779_in     : std_logic;
  signal reg_q779_init   : std_logic;
		

  -- state q91
  signal reg_q91        : std_logic;
  signal reg_q91_in     : std_logic;
  signal reg_q91_init   : std_logic;
		
--#################################################
-- start section fullgraph: 54

  -- state q844
  signal reg_q844        : std_logic;
  signal reg_q844_in     : std_logic;
  		

  -- state q1645
  signal reg_q1645        : std_logic;
  signal reg_q1645_in     : std_logic;
  		

  -- state q834
  signal reg_q834        : std_logic;
  signal reg_q834_in     : std_logic;
  		

  -- state q1882
  signal reg_q1882        : std_logic;
  signal reg_q1882_in     : std_logic;
  		

  -- state q620
  signal reg_q620        : std_logic;
  signal reg_q620_in     : std_logic;
  		

  -- state q2387
  signal reg_q2387        : std_logic;
  signal reg_q2387_in     : std_logic;
  		

  -- state q454
  signal reg_q454        : std_logic;
  signal reg_q454_in     : std_logic;
  		

  -- state q1197
  signal reg_q1197        : std_logic;
  signal reg_q1197_in     : std_logic;
  		

  -- state q846
  signal reg_q846        : std_logic;
  signal reg_q846_in     : std_logic;
  		

  -- state q2389
  signal reg_q2389        : std_logic;
  signal reg_q2389_in     : std_logic;
  		
  signal reg_fullgraph54       : std_logic_vector(3 downto 0);
  signal reg_fullgraph54_in    : std_logic_vector(3 downto 0);
  signal reg_fullgraph54_init  : std_logic_vector(3 downto 0);
  signal reg_fullgraph54_sel   : std_logic_vector(15 downto 0); 	
  -- end section fullgraph54
  --#################################################			
		
--#################################################
-- start section fullgraph: 55

  -- state q1768
  signal reg_q1768        : std_logic;
  signal reg_q1768_in     : std_logic;
  		

  -- state q836
  signal reg_q836        : std_logic;
  signal reg_q836_in     : std_logic;
  		

  -- state q838
  signal reg_q838        : std_logic;
  signal reg_q838_in     : std_logic;
  		

  -- state q1828
  signal reg_q1828        : std_logic;
  signal reg_q1828_in     : std_logic;
  		
  signal reg_fullgraph55       : std_logic_vector(2 downto 0);
  signal reg_fullgraph55_in    : std_logic_vector(2 downto 0);
  signal reg_fullgraph55_init  : std_logic_vector(2 downto 0);
  signal reg_fullgraph55_sel   : std_logic_vector(7 downto 0); 	
  -- end section fullgraph55
  --#################################################			
		
--#################################################
-- start section fullgraph: 56

  -- state q817
  signal reg_q817        : std_logic;
  signal reg_q817_in     : std_logic;
  		

  -- state q840
  signal reg_q840        : std_logic;
  signal reg_q840_in     : std_logic;
  		
  signal reg_fullgraph56       : std_logic_vector(1 downto 0);
  signal reg_fullgraph56_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph56_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph56_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph56
  --#################################################			
		
--#################################################
-- start section fullgraph: 57

  -- state q1782
  signal reg_q1782        : std_logic;
  signal reg_q1782_in     : std_logic;
  		

  -- state q2
  signal reg_q2        : std_logic;
  signal reg_q2_in     : std_logic;
  		
  signal reg_fullgraph57       : std_logic_vector(1 downto 0);
  signal reg_fullgraph57_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph57_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph57_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph57
  --#################################################			
		
--#################################################
-- start section fullgraph: 58

  -- state q1784
  signal reg_q1784        : std_logic;
  signal reg_q1784_in     : std_logic;
  		

  -- state q4
  signal reg_q4        : std_logic;
  signal reg_q4_in     : std_logic;
  		
  signal reg_fullgraph58       : std_logic_vector(1 downto 0);
  signal reg_fullgraph58_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph58_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph58_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph58
  --#################################################			
		
--#################################################
-- start section fullgraph: 59

  -- state q2092
  signal reg_q2092        : std_logic;
  signal reg_q2092_in     : std_logic;
  		

  -- state q6
  signal reg_q6        : std_logic;
  signal reg_q6_in     : std_logic;
  		
  signal reg_fullgraph59       : std_logic_vector(1 downto 0);
  signal reg_fullgraph59_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph59_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph59_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph59
  --#################################################			
		

  -- state q1225
  signal reg_q1225        : std_logic;
  signal reg_q1225_in     : std_logic;
  signal reg_q1225_init   : std_logic;
		
--#################################################
-- start section fullgraph: 61

  -- state q2583
  signal reg_q2583        : std_logic;
  signal reg_q2583_in     : std_logic;
  		

  -- state q2585
  signal reg_q2585        : std_logic;
  signal reg_q2585_in     : std_logic;
  		
  signal reg_fullgraph61       : std_logic_vector(1 downto 0);
  signal reg_fullgraph61_in    : std_logic_vector(1 downto 0);
  signal reg_fullgraph61_init  : std_logic_vector(1 downto 0);
  signal reg_fullgraph61_sel   : std_logic_vector(3 downto 0); 	
  -- end section fullgraph61
  --#################################################			
		

  -- state q2001
  signal reg_q2001        : std_logic;
  signal reg_q2001_in     : std_logic;
  signal reg_q2001_init   : std_logic;
		

  -- state q681
  signal reg_q681        : std_logic;
  signal reg_q681_in     : std_logic;
  signal reg_q681_init   : std_logic;
		

  -- state q1754
  signal reg_q1754        : std_logic;
  signal reg_q1754_in     : std_logic;
  signal reg_q1754_init   : std_logic;
		

  -- state q1756
  signal reg_q1756        : std_logic;
  signal reg_q1756_in     : std_logic;
  signal reg_q1756_init   : std_logic;
		

  -- state q959
  signal reg_q959        : std_logic;
  signal reg_q959_in     : std_logic;
  signal reg_q959_init   : std_logic;
		

  -- state q900
  signal reg_q900        : std_logic;
  signal reg_q900_in     : std_logic;
  signal reg_q900_init   : std_logic;
		

  -- state q304
  signal reg_q304        : std_logic;
  signal reg_q304_in     : std_logic;
  signal reg_q304_init   : std_logic;
		

  -- state q1786
  signal reg_q1786        : std_logic;
  signal reg_q1786_in     : std_logic;
  signal reg_q1786_init   : std_logic;
		

  -- state q1788
  signal reg_q1788        : std_logic;
  signal reg_q1788_in     : std_logic;
  signal reg_q1788_init   : std_logic;
		

  -- state q1746
  signal reg_q1746        : std_logic;
  signal reg_q1746_in     : std_logic;
  signal reg_q1746_init   : std_logic;
		

  -- state q1748
  signal reg_q1748        : std_logic;
  signal reg_q1748_in     : std_logic;
  signal reg_q1748_init   : std_logic;
		

  -- state q1051
  signal reg_q1051        : std_logic;
  signal reg_q1051_in     : std_logic;
  signal reg_q1051_init   : std_logic;
		

  -- state q1764
  signal reg_q1764        : std_logic;
  signal reg_q1764_in     : std_logic;
  signal reg_q1764_init   : std_logic;
		

  -- state q1766
  signal reg_q1766        : std_logic;
  signal reg_q1766_in     : std_logic;
  signal reg_q1766_init   : std_logic;
		

  -- state q1453
  signal reg_q1453        : std_logic;
  signal reg_q1453_in     : std_logic;
  signal reg_q1453_init   : std_logic;
		

  -- state q1744
  signal reg_q1744        : std_logic;
  signal reg_q1744_in     : std_logic;
  signal reg_q1744_init   : std_logic;
		

  -- state q1774
  signal reg_q1774        : std_logic;
  signal reg_q1774_in     : std_logic;
  signal reg_q1774_init   : std_logic;
		

  -- state q1776
  signal reg_q1776        : std_logic;
  signal reg_q1776_in     : std_logic;
  signal reg_q1776_init   : std_logic;
		

  -- state q1014
  signal reg_q1014        : std_logic;
  signal reg_q1014_in     : std_logic;
  signal reg_q1014_init   : std_logic;
		

  -- state q1545
  signal reg_q1545        : std_logic;
  signal reg_q1545_in     : std_logic;
  signal reg_q1545_init   : std_logic;
		

  -- state q1780
  signal reg_q1780        : std_logic;
  signal reg_q1780_in     : std_logic;
  signal reg_q1780_init   : std_logic;
		

  -- state q2619
  signal reg_q2619        : std_logic;
  signal reg_q2619_in     : std_logic;
  signal reg_q2619_init   : std_logic;
		

  -- state q666
  signal reg_q666        : std_logic;
  signal reg_q666_in     : std_logic;
  signal reg_q666_init   : std_logic;
		

  -- state q2324
  signal reg_q2324        : std_logic;
  signal reg_q2324_in     : std_logic;
  signal reg_q2324_init   : std_logic;
		

  -- state q1752
  signal reg_q1752        : std_logic;
  signal reg_q1752_in     : std_logic;
  signal reg_q1752_init   : std_logic;
		

  -- state q704
  signal reg_q704        : std_logic;
  signal reg_q704_in     : std_logic;
  signal reg_q704_init   : std_logic;
		

  -- state q1522
  signal reg_q1522        : std_logic;
  signal reg_q1522_in     : std_logic;
  signal reg_q1522_init   : std_logic;
		

  -- state q1956
  signal reg_q1956        : std_logic;
  signal reg_q1956_in     : std_logic;
  signal reg_q1956_init   : std_logic;
		

  -- state q2534
  signal reg_q2534        : std_logic;
  signal reg_q2534_in     : std_logic;
  signal reg_q2534_init   : std_logic;
		

  -- state q780
  signal reg_q780        : std_logic;
  signal reg_q780_in     : std_logic;
  signal reg_q780_init   : std_logic;
		

  -- state q715
  signal reg_q715        : std_logic;
  signal reg_q715_in     : std_logic;
  signal reg_q715_init   : std_logic;
		

  -- state q1778
  signal reg_q1778        : std_logic;
  signal reg_q1778_in     : std_logic;
  signal reg_q1778_init   : std_logic;
		

  -- state q1604
  signal reg_q1604        : std_logic;
  signal reg_q1604_in     : std_logic;
  signal reg_q1604_init   : std_logic;
		

  -- state q2212
  signal reg_q2212        : std_logic;
  signal reg_q2212_in     : std_logic;
  signal reg_q2212_init   : std_logic;
		

  -- state q226
  signal reg_q226        : std_logic;
  signal reg_q226_in     : std_logic;
  signal reg_q226_init   : std_logic;
		

  -- state q2125
  signal reg_q2125        : std_logic;
  signal reg_q2125_in     : std_logic;
  signal reg_q2125_init   : std_logic;
		

  -- state q47
  signal reg_q47        : std_logic;
  signal reg_q47_in     : std_logic;
  signal reg_q47_init   : std_logic;
		

  -- state q1762
  signal reg_q1762        : std_logic;
  signal reg_q1762_in     : std_logic;
  signal reg_q1762_init   : std_logic;
		

  -- state q1760
  signal reg_q1760        : std_logic;
  signal reg_q1760_in     : std_logic;
  signal reg_q1760_init   : std_logic;
		

  -- state q415
  signal reg_q415        : std_logic;
  signal reg_q415_in     : std_logic;
  signal reg_q415_init   : std_logic;
		

  -- state q179
  signal reg_q179        : std_logic;
  signal reg_q179_in     : std_logic;
  signal reg_q179_init   : std_logic;
		

  -- state q1758
  signal reg_q1758        : std_logic;
  signal reg_q1758_in     : std_logic;
  signal reg_q1758_init   : std_logic;
		

  -- state q1750
  signal reg_q1750        : std_logic;
  signal reg_q1750_in     : std_logic;
  signal reg_q1750_init   : std_logic;
		

  -- state q2253
  signal reg_q2253        : std_logic;
  signal reg_q2253_in     : std_logic;
  signal reg_q2253_init   : std_logic;
		

  -- state q263
  signal reg_q263        : std_logic;
  signal reg_q263_in     : std_logic;
  signal reg_q263_init   : std_logic;
		

  -- state q92
  signal reg_q92        : std_logic;
  signal reg_q92_in     : std_logic;
  signal reg_q92_init   : std_logic;
		

  -- symbol decoder
  signal symb_decoder : std_logic_vector(2**DATA_WIDTH - 1 downto 0);

  -- intialization signal
  signal initialize   : std_logic;

	begin
	-- initialization
  	initialize <= INIT OR INPUT_EOF; 
	 
		symb_decoder(16#f5#) <= '1' when (INPUT = X"f5") else
                          '0';
		symb_decoder(16#b3#) <= '1' when (INPUT = X"b3") else
                          '0';
		symb_decoder(16#ea#) <= '1' when (INPUT = X"ea") else
                          '0';
		symb_decoder(16#d7#) <= '1' when (INPUT = X"d7") else
                          '0';
		symb_decoder(16#d5#) <= '1' when (INPUT = X"d5") else
                          '0';
		symb_decoder(16#a4#) <= '1' when (INPUT = X"a4") else
                          '0';
		symb_decoder(16#49#) <= '1' when (INPUT = X"49") else
                          '0';
		symb_decoder(16#85#) <= '1' when (INPUT = X"85") else
                          '0';
		symb_decoder(16#3a#) <= '1' when (INPUT = X"3a") else
                          '0';
		symb_decoder(16#2c#) <= '1' when (INPUT = X"2c") else
                          '0';
		symb_decoder(16#c1#) <= '1' when (INPUT = X"c1") else
                          '0';
		symb_decoder(16#ba#) <= '1' when (INPUT = X"ba") else
                          '0';
		symb_decoder(16#0f#) <= '1' when (INPUT = X"0f") else
                          '0';
		symb_decoder(16#df#) <= '1' when (INPUT = X"df") else
                          '0';
		symb_decoder(16#66#) <= '1' when (INPUT = X"66") else
                          '0';
		symb_decoder(16#e8#) <= '1' when (INPUT = X"e8") else
                          '0';
		symb_decoder(16#2d#) <= '1' when (INPUT = X"2d") else
                          '0';
		symb_decoder(16#bf#) <= '1' when (INPUT = X"bf") else
                          '0';
		symb_decoder(16#7a#) <= '1' when (INPUT = X"7a") else
                          '0';
		symb_decoder(16#31#) <= '1' when (INPUT = X"31") else
                          '0';
		symb_decoder(16#97#) <= '1' when (INPUT = X"97") else
                          '0';
		symb_decoder(16#93#) <= '1' when (INPUT = X"93") else
                          '0';
		symb_decoder(16#11#) <= '1' when (INPUT = X"11") else
                          '0';
		symb_decoder(16#1d#) <= '1' when (INPUT = X"1d") else
                          '0';
		symb_decoder(16#6f#) <= '1' when (INPUT = X"6f") else
                          '0';
		symb_decoder(16#f6#) <= '1' when (INPUT = X"f6") else
                          '0';
		symb_decoder(16#50#) <= '1' when (INPUT = X"50") else
                          '0';
		symb_decoder(16#de#) <= '1' when (INPUT = X"de") else
                          '0';
		symb_decoder(16#1f#) <= '1' when (INPUT = X"1f") else
                          '0';
		symb_decoder(16#6c#) <= '1' when (INPUT = X"6c") else
                          '0';
		symb_decoder(16#59#) <= '1' when (INPUT = X"59") else
                          '0';
		symb_decoder(16#39#) <= '1' when (INPUT = X"39") else
                          '0';
		symb_decoder(16#7d#) <= '1' when (INPUT = X"7d") else
                          '0';
		symb_decoder(16#d2#) <= '1' when (INPUT = X"d2") else
                          '0';
		symb_decoder(16#27#) <= '1' when (INPUT = X"27") else
                          '0';
		symb_decoder(16#2f#) <= '1' when (INPUT = X"2f") else
                          '0';
		symb_decoder(16#8d#) <= '1' when (INPUT = X"8d") else
                          '0';
		symb_decoder(16#a7#) <= '1' when (INPUT = X"a7") else
                          '0';
		symb_decoder(16#e2#) <= '1' when (INPUT = X"e2") else
                          '0';
		symb_decoder(16#c3#) <= '1' when (INPUT = X"c3") else
                          '0';
		symb_decoder(16#67#) <= '1' when (INPUT = X"67") else
                          '0';
		symb_decoder(16#38#) <= '1' when (INPUT = X"38") else
                          '0';
		symb_decoder(16#ad#) <= '1' when (INPUT = X"ad") else
                          '0';
		symb_decoder(16#cc#) <= '1' when (INPUT = X"cc") else
                          '0';
		symb_decoder(16#01#) <= '1' when (INPUT = X"01") else
                          '0';
		symb_decoder(16#ec#) <= '1' when (INPUT = X"ec") else
                          '0';
		symb_decoder(16#15#) <= '1' when (INPUT = X"15") else
                          '0';
		symb_decoder(16#c5#) <= '1' when (INPUT = X"c5") else
                          '0';
		symb_decoder(16#ef#) <= '1' when (INPUT = X"ef") else
                          '0';
		symb_decoder(16#e5#) <= '1' when (INPUT = X"e5") else
                          '0';
		symb_decoder(16#a9#) <= '1' when (INPUT = X"a9") else
                          '0';
		symb_decoder(16#6e#) <= '1' when (INPUT = X"6e") else
                          '0';
		symb_decoder(16#4a#) <= '1' when (INPUT = X"4a") else
                          '0';
		symb_decoder(16#9c#) <= '1' when (INPUT = X"9c") else
                          '0';
		symb_decoder(16#9f#) <= '1' when (INPUT = X"9f") else
                          '0';
		symb_decoder(16#54#) <= '1' when (INPUT = X"54") else
                          '0';
		symb_decoder(16#42#) <= '1' when (INPUT = X"42") else
                          '0';
		symb_decoder(16#cd#) <= '1' when (INPUT = X"cd") else
                          '0';
		symb_decoder(16#63#) <= '1' when (INPUT = X"63") else
                          '0';
		symb_decoder(16#dd#) <= '1' when (INPUT = X"dd") else
                          '0';
		symb_decoder(16#19#) <= '1' when (INPUT = X"19") else
                          '0';
		symb_decoder(16#d1#) <= '1' when (INPUT = X"d1") else
                          '0';
		symb_decoder(16#72#) <= '1' when (INPUT = X"72") else
                          '0';
		symb_decoder(16#7f#) <= '1' when (INPUT = X"7f") else
                          '0';
		symb_decoder(16#75#) <= '1' when (INPUT = X"75") else
                          '0';
		symb_decoder(16#08#) <= '1' when (INPUT = X"08") else
                          '0';
		symb_decoder(16#1c#) <= '1' when (INPUT = X"1c") else
                          '0';
		symb_decoder(16#6d#) <= '1' when (INPUT = X"6d") else
                          '0';
		symb_decoder(16#f8#) <= '1' when (INPUT = X"f8") else
                          '0';
		symb_decoder(16#16#) <= '1' when (INPUT = X"16") else
                          '0';
		symb_decoder(16#35#) <= '1' when (INPUT = X"35") else
                          '0';
		symb_decoder(16#e7#) <= '1' when (INPUT = X"e7") else
                          '0';
		symb_decoder(16#ce#) <= '1' when (INPUT = X"ce") else
                          '0';
		symb_decoder(16#b2#) <= '1' when (INPUT = X"b2") else
                          '0';
		symb_decoder(16#14#) <= '1' when (INPUT = X"14") else
                          '0';
		symb_decoder(16#6b#) <= '1' when (INPUT = X"6b") else
                          '0';
		symb_decoder(16#7c#) <= '1' when (INPUT = X"7c") else
                          '0';
		symb_decoder(16#e9#) <= '1' when (INPUT = X"e9") else
                          '0';
		symb_decoder(16#2b#) <= '1' when (INPUT = X"2b") else
                          '0';
		symb_decoder(16#d4#) <= '1' when (INPUT = X"d4") else
                          '0';
		symb_decoder(16#ab#) <= '1' when (INPUT = X"ab") else
                          '0';
		symb_decoder(16#5a#) <= '1' when (INPUT = X"5a") else
                          '0';
		symb_decoder(16#82#) <= '1' when (INPUT = X"82") else
                          '0';
		symb_decoder(16#5f#) <= '1' when (INPUT = X"5f") else
                          '0';
		symb_decoder(16#a5#) <= '1' when (INPUT = X"a5") else
                          '0';
		symb_decoder(16#83#) <= '1' when (INPUT = X"83") else
                          '0';
		symb_decoder(16#37#) <= '1' when (INPUT = X"37") else
                          '0';
		symb_decoder(16#84#) <= '1' when (INPUT = X"84") else
                          '0';
		symb_decoder(16#87#) <= '1' when (INPUT = X"87") else
                          '0';
		symb_decoder(16#fa#) <= '1' when (INPUT = X"fa") else
                          '0';
		symb_decoder(16#04#) <= '1' when (INPUT = X"04") else
                          '0';
		symb_decoder(16#9b#) <= '1' when (INPUT = X"9b") else
                          '0';
		symb_decoder(16#55#) <= '1' when (INPUT = X"55") else
                          '0';
		symb_decoder(16#1a#) <= '1' when (INPUT = X"1a") else
                          '0';
		symb_decoder(16#c8#) <= '1' when (INPUT = X"c8") else
                          '0';
		symb_decoder(16#58#) <= '1' when (INPUT = X"58") else
                          '0';
		symb_decoder(16#b9#) <= '1' when (INPUT = X"b9") else
                          '0';
		symb_decoder(16#db#) <= '1' when (INPUT = X"db") else
                          '0';
		symb_decoder(16#cf#) <= '1' when (INPUT = X"cf") else
                          '0';
		symb_decoder(16#0e#) <= '1' when (INPUT = X"0e") else
                          '0';
		symb_decoder(16#76#) <= '1' when (INPUT = X"76") else
                          '0';
		symb_decoder(16#06#) <= '1' when (INPUT = X"06") else
                          '0';
		symb_decoder(16#9e#) <= '1' when (INPUT = X"9e") else
                          '0';
		symb_decoder(16#9a#) <= '1' when (INPUT = X"9a") else
                          '0';
		symb_decoder(16#d6#) <= '1' when (INPUT = X"d6") else
                          '0';
		symb_decoder(16#62#) <= '1' when (INPUT = X"62") else
                          '0';
		symb_decoder(16#23#) <= '1' when (INPUT = X"23") else
                          '0';
		symb_decoder(16#43#) <= '1' when (INPUT = X"43") else
                          '0';
		symb_decoder(16#bd#) <= '1' when (INPUT = X"bd") else
                          '0';
		symb_decoder(16#8f#) <= '1' when (INPUT = X"8f") else
                          '0';
		symb_decoder(16#1e#) <= '1' when (INPUT = X"1e") else
                          '0';
		symb_decoder(16#61#) <= '1' when (INPUT = X"61") else
                          '0';
		symb_decoder(16#f2#) <= '1' when (INPUT = X"f2") else
                          '0';
		symb_decoder(16#5e#) <= '1' when (INPUT = X"5e") else
                          '0';
		symb_decoder(16#86#) <= '1' when (INPUT = X"86") else
                          '0';
		symb_decoder(16#a3#) <= '1' when (INPUT = X"a3") else
                          '0';
		symb_decoder(16#fd#) <= '1' when (INPUT = X"fd") else
                          '0';
		symb_decoder(16#ff#) <= '1' when (INPUT = X"ff") else
                          '0';
		symb_decoder(16#17#) <= '1' when (INPUT = X"17") else
                          '0';
		symb_decoder(16#2a#) <= '1' when (INPUT = X"2a") else
                          '0';
		symb_decoder(16#5b#) <= '1' when (INPUT = X"5b") else
                          '0';
		symb_decoder(16#28#) <= '1' when (INPUT = X"28") else
                          '0';
		symb_decoder(16#3f#) <= '1' when (INPUT = X"3f") else
                          '0';
		symb_decoder(16#89#) <= '1' when (INPUT = X"89") else
                          '0';
		symb_decoder(16#6a#) <= '1' when (INPUT = X"6a") else
                          '0';
		symb_decoder(16#0a#) <= '1' when (INPUT = X"0a") else
                          '0';
		symb_decoder(16#00#) <= '1' when (INPUT = X"00") else
                          '0';
		symb_decoder(16#c7#) <= '1' when (INPUT = X"c7") else
                          '0';
		symb_decoder(16#4c#) <= '1' when (INPUT = X"4c") else
                          '0';
		symb_decoder(16#03#) <= '1' when (INPUT = X"03") else
                          '0';
		symb_decoder(16#57#) <= '1' when (INPUT = X"57") else
                          '0';
		symb_decoder(16#d8#) <= '1' when (INPUT = X"d8") else
                          '0';
		symb_decoder(16#eb#) <= '1' when (INPUT = X"eb") else
                          '0';
		symb_decoder(16#a2#) <= '1' when (INPUT = X"a2") else
                          '0';
		symb_decoder(16#1b#) <= '1' when (INPUT = X"1b") else
                          '0';
		symb_decoder(16#b1#) <= '1' when (INPUT = X"b1") else
                          '0';
		symb_decoder(16#b0#) <= '1' when (INPUT = X"b0") else
                          '0';
		symb_decoder(16#12#) <= '1' when (INPUT = X"12") else
                          '0';
		symb_decoder(16#05#) <= '1' when (INPUT = X"05") else
                          '0';
		symb_decoder(16#7b#) <= '1' when (INPUT = X"7b") else
                          '0';
		symb_decoder(16#c6#) <= '1' when (INPUT = X"c6") else
                          '0';
		symb_decoder(16#53#) <= '1' when (INPUT = X"53") else
                          '0';
		symb_decoder(16#45#) <= '1' when (INPUT = X"45") else
                          '0';
		symb_decoder(16#91#) <= '1' when (INPUT = X"91") else
                          '0';
		symb_decoder(16#21#) <= '1' when (INPUT = X"21") else
                          '0';
		symb_decoder(16#7e#) <= '1' when (INPUT = X"7e") else
                          '0';
		symb_decoder(16#a1#) <= '1' when (INPUT = X"a1") else
                          '0';
		symb_decoder(16#c0#) <= '1' when (INPUT = X"c0") else
                          '0';
		symb_decoder(16#4f#) <= '1' when (INPUT = X"4f") else
                          '0';
		symb_decoder(16#48#) <= '1' when (INPUT = X"48") else
                          '0';
		symb_decoder(16#fc#) <= '1' when (INPUT = X"fc") else
                          '0';
		symb_decoder(16#44#) <= '1' when (INPUT = X"44") else
                          '0';
		symb_decoder(16#4b#) <= '1' when (INPUT = X"4b") else
                          '0';
		symb_decoder(16#d0#) <= '1' when (INPUT = X"d0") else
                          '0';
		symb_decoder(16#40#) <= '1' when (INPUT = X"40") else
                          '0';
		symb_decoder(16#34#) <= '1' when (INPUT = X"34") else
                          '0';
		symb_decoder(16#ca#) <= '1' when (INPUT = X"ca") else
                          '0';
		symb_decoder(16#81#) <= '1' when (INPUT = X"81") else
                          '0';
		symb_decoder(16#70#) <= '1' when (INPUT = X"70") else
                          '0';
		symb_decoder(16#b8#) <= '1' when (INPUT = X"b8") else
                          '0';
		symb_decoder(16#bb#) <= '1' when (INPUT = X"bb") else
                          '0';
		symb_decoder(16#a0#) <= '1' when (INPUT = X"a0") else
                          '0';
		symb_decoder(16#30#) <= '1' when (INPUT = X"30") else
                          '0';
		symb_decoder(16#60#) <= '1' when (INPUT = X"60") else
                          '0';
		symb_decoder(16#13#) <= '1' when (INPUT = X"13") else
                          '0';
		symb_decoder(16#e0#) <= '1' when (INPUT = X"e0") else
                          '0';
		symb_decoder(16#94#) <= '1' when (INPUT = X"94") else
                          '0';
		symb_decoder(16#e1#) <= '1' when (INPUT = X"e1") else
                          '0';
		symb_decoder(16#ed#) <= '1' when (INPUT = X"ed") else
                          '0';
		symb_decoder(16#41#) <= '1' when (INPUT = X"41") else
                          '0';
		symb_decoder(16#b4#) <= '1' when (INPUT = X"b4") else
                          '0';
		symb_decoder(16#be#) <= '1' when (INPUT = X"be") else
                          '0';
		symb_decoder(16#e3#) <= '1' when (INPUT = X"e3") else
                          '0';
		symb_decoder(16#25#) <= '1' when (INPUT = X"25") else
                          '0';
		symb_decoder(16#02#) <= '1' when (INPUT = X"02") else
                          '0';
		symb_decoder(16#22#) <= '1' when (INPUT = X"22") else
                          '0';
		symb_decoder(16#36#) <= '1' when (INPUT = X"36") else
                          '0';
		symb_decoder(16#52#) <= '1' when (INPUT = X"52") else
                          '0';
		symb_decoder(16#ae#) <= '1' when (INPUT = X"ae") else
                          '0';
		symb_decoder(16#09#) <= '1' when (INPUT = X"09") else
                          '0';
		symb_decoder(16#0d#) <= '1' when (INPUT = X"0d") else
                          '0';
		symb_decoder(16#c2#) <= '1' when (INPUT = X"c2") else
                          '0';
		symb_decoder(16#26#) <= '1' when (INPUT = X"26") else
                          '0';
		symb_decoder(16#c9#) <= '1' when (INPUT = X"c9") else
                          '0';
		symb_decoder(16#f9#) <= '1' when (INPUT = X"f9") else
                          '0';
		symb_decoder(16#8a#) <= '1' when (INPUT = X"8a") else
                          '0';
		symb_decoder(16#4d#) <= '1' when (INPUT = X"4d") else
                          '0';
		symb_decoder(16#3d#) <= '1' when (INPUT = X"3d") else
                          '0';
		symb_decoder(16#bc#) <= '1' when (INPUT = X"bc") else
                          '0';
		symb_decoder(16#dc#) <= '1' when (INPUT = X"dc") else
                          '0';
		symb_decoder(16#f7#) <= '1' when (INPUT = X"f7") else
                          '0';
		symb_decoder(16#8c#) <= '1' when (INPUT = X"8c") else
                          '0';
		symb_decoder(16#aa#) <= '1' when (INPUT = X"aa") else
                          '0';
		symb_decoder(16#f3#) <= '1' when (INPUT = X"f3") else
                          '0';
		symb_decoder(16#77#) <= '1' when (INPUT = X"77") else
                          '0';
		symb_decoder(16#ac#) <= '1' when (INPUT = X"ac") else
                          '0';
		symb_decoder(16#0c#) <= '1' when (INPUT = X"0c") else
                          '0';
		symb_decoder(16#95#) <= '1' when (INPUT = X"95") else
                          '0';
		symb_decoder(16#98#) <= '1' when (INPUT = X"98") else
                          '0';
		symb_decoder(16#b7#) <= '1' when (INPUT = X"b7") else
                          '0';
		symb_decoder(16#73#) <= '1' when (INPUT = X"73") else
                          '0';
		symb_decoder(16#51#) <= '1' when (INPUT = X"51") else
                          '0';
		symb_decoder(16#20#) <= '1' when (INPUT = X"20") else
                          '0';
		symb_decoder(16#e6#) <= '1' when (INPUT = X"e6") else
                          '0';
		symb_decoder(16#4e#) <= '1' when (INPUT = X"4e") else
                          '0';
		symb_decoder(16#e4#) <= '1' when (INPUT = X"e4") else
                          '0';
		symb_decoder(16#74#) <= '1' when (INPUT = X"74") else
                          '0';
		symb_decoder(16#71#) <= '1' when (INPUT = X"71") else
                          '0';
		symb_decoder(16#a6#) <= '1' when (INPUT = X"a6") else
                          '0';
		symb_decoder(16#f4#) <= '1' when (INPUT = X"f4") else
                          '0';
		symb_decoder(16#2e#) <= '1' when (INPUT = X"2e") else
                          '0';
		symb_decoder(16#5d#) <= '1' when (INPUT = X"5d") else
                          '0';
		symb_decoder(16#64#) <= '1' when (INPUT = X"64") else
                          '0';
		symb_decoder(16#78#) <= '1' when (INPUT = X"78") else
                          '0';
		symb_decoder(16#80#) <= '1' when (INPUT = X"80") else
                          '0';
		symb_decoder(16#fb#) <= '1' when (INPUT = X"fb") else
                          '0';
		symb_decoder(16#29#) <= '1' when (INPUT = X"29") else
                          '0';
		symb_decoder(16#b5#) <= '1' when (INPUT = X"b5") else
                          '0';
		symb_decoder(16#24#) <= '1' when (INPUT = X"24") else
                          '0';
		symb_decoder(16#88#) <= '1' when (INPUT = X"88") else
                          '0';
		symb_decoder(16#f1#) <= '1' when (INPUT = X"f1") else
                          '0';
		symb_decoder(16#fe#) <= '1' when (INPUT = X"fe") else
                          '0';
		symb_decoder(16#92#) <= '1' when (INPUT = X"92") else
                          '0';
		symb_decoder(16#68#) <= '1' when (INPUT = X"68") else
                          '0';
		symb_decoder(16#ee#) <= '1' when (INPUT = X"ee") else
                          '0';
		symb_decoder(16#46#) <= '1' when (INPUT = X"46") else
                          '0';
		symb_decoder(16#af#) <= '1' when (INPUT = X"af") else
                          '0';
		symb_decoder(16#33#) <= '1' when (INPUT = X"33") else
                          '0';
		symb_decoder(16#8e#) <= '1' when (INPUT = X"8e") else
                          '0';
		symb_decoder(16#8b#) <= '1' when (INPUT = X"8b") else
                          '0';
		symb_decoder(16#79#) <= '1' when (INPUT = X"79") else
                          '0';
		symb_decoder(16#07#) <= '1' when (INPUT = X"07") else
                          '0';
		symb_decoder(16#32#) <= '1' when (INPUT = X"32") else
                          '0';
		symb_decoder(16#5c#) <= '1' when (INPUT = X"5c") else
                          '0';
		symb_decoder(16#a8#) <= '1' when (INPUT = X"a8") else
                          '0';
		symb_decoder(16#56#) <= '1' when (INPUT = X"56") else
                          '0';
		symb_decoder(16#10#) <= '1' when (INPUT = X"10") else
                          '0';
		symb_decoder(16#3e#) <= '1' when (INPUT = X"3e") else
                          '0';
		symb_decoder(16#cb#) <= '1' when (INPUT = X"cb") else
                          '0';
		symb_decoder(16#b6#) <= '1' when (INPUT = X"b6") else
                          '0';
		symb_decoder(16#3c#) <= '1' when (INPUT = X"3c") else
                          '0';
		symb_decoder(16#90#) <= '1' when (INPUT = X"90") else
                          '0';
		symb_decoder(16#9d#) <= '1' when (INPUT = X"9d") else
                          '0';
		symb_decoder(16#3b#) <= '1' when (INPUT = X"3b") else
                          '0';
		symb_decoder(16#65#) <= '1' when (INPUT = X"65") else
                          '0';
		symb_decoder(16#99#) <= '1' when (INPUT = X"99") else
                          '0';
		symb_decoder(16#d9#) <= '1' when (INPUT = X"d9") else
                          '0';
		symb_decoder(16#0b#) <= '1' when (INPUT = X"0b") else
                          '0';
		symb_decoder(16#f0#) <= '1' when (INPUT = X"f0") else
                          '0';
		symb_decoder(16#18#) <= '1' when (INPUT = X"18") else
                          '0';
		symb_decoder(16#c4#) <= '1' when (INPUT = X"c4") else
                          '0';
		symb_decoder(16#69#) <= '1' when (INPUT = X"69") else
                          '0';
		symb_decoder(16#96#) <= '1' when (INPUT = X"96") else
                          '0';
		symb_decoder(16#d3#) <= '1' when (INPUT = X"d3") else
                          '0';
		symb_decoder(16#da#) <= '1' when (INPUT = X"da") else
                          '0';
		symb_decoder(16#47#) <= '1' when (INPUT = X"47") else
                          '0';

--######################################################
--fullgraph0

reg_q2695_in <= '0';
reg_q1452_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1452 AND symb_decoder(16#2f#)) OR
 					(reg_q1452 AND symb_decoder(16#85#)) OR
 					(reg_q1452 AND symb_decoder(16#e9#)) OR
 					(reg_q1452 AND symb_decoder(16#77#)) OR
 					(reg_q1452 AND symb_decoder(16#f4#)) OR
 					(reg_q1452 AND symb_decoder(16#7a#)) OR
 					(reg_q1452 AND symb_decoder(16#a9#)) OR
 					(reg_q1452 AND symb_decoder(16#45#)) OR
 					(reg_q1452 AND symb_decoder(16#9b#)) OR
 					(reg_q1452 AND symb_decoder(16#75#)) OR
 					(reg_q1452 AND symb_decoder(16#cf#)) OR
 					(reg_q1452 AND symb_decoder(16#88#)) OR
 					(reg_q1452 AND symb_decoder(16#a1#)) OR
 					(reg_q1452 AND symb_decoder(16#53#)) OR
 					(reg_q1452 AND symb_decoder(16#6a#)) OR
 					(reg_q1452 AND symb_decoder(16#74#)) OR
 					(reg_q1452 AND symb_decoder(16#ce#)) OR
 					(reg_q1452 AND symb_decoder(16#ee#)) OR
 					(reg_q1452 AND symb_decoder(16#79#)) OR
 					(reg_q1452 AND symb_decoder(16#e0#)) OR
 					(reg_q1452 AND symb_decoder(16#70#)) OR
 					(reg_q1452 AND symb_decoder(16#5e#)) OR
 					(reg_q1452 AND symb_decoder(16#fc#)) OR
 					(reg_q1452 AND symb_decoder(16#35#)) OR
 					(reg_q1452 AND symb_decoder(16#3e#)) OR
 					(reg_q1452 AND symb_decoder(16#7c#)) OR
 					(reg_q1452 AND symb_decoder(16#fa#)) OR
 					(reg_q1452 AND symb_decoder(16#d9#)) OR
 					(reg_q1452 AND symb_decoder(16#fd#)) OR
 					(reg_q1452 AND symb_decoder(16#f6#)) OR
 					(reg_q1452 AND symb_decoder(16#84#)) OR
 					(reg_q1452 AND symb_decoder(16#4f#)) OR
 					(reg_q1452 AND symb_decoder(16#9c#)) OR
 					(reg_q1452 AND symb_decoder(16#fb#)) OR
 					(reg_q1452 AND symb_decoder(16#b4#)) OR
 					(reg_q1452 AND symb_decoder(16#1a#)) OR
 					(reg_q1452 AND symb_decoder(16#63#)) OR
 					(reg_q1452 AND symb_decoder(16#03#)) OR
 					(reg_q1452 AND symb_decoder(16#9e#)) OR
 					(reg_q1452 AND symb_decoder(16#6d#)) OR
 					(reg_q1452 AND symb_decoder(16#ec#)) OR
 					(reg_q1452 AND symb_decoder(16#c4#)) OR
 					(reg_q1452 AND symb_decoder(16#6b#)) OR
 					(reg_q1452 AND symb_decoder(16#dd#)) OR
 					(reg_q1452 AND symb_decoder(16#14#)) OR
 					(reg_q1452 AND symb_decoder(16#39#)) OR
 					(reg_q1452 AND symb_decoder(16#cb#)) OR
 					(reg_q1452 AND symb_decoder(16#49#)) OR
 					(reg_q1452 AND symb_decoder(16#40#)) OR
 					(reg_q1452 AND symb_decoder(16#5b#)) OR
 					(reg_q1452 AND symb_decoder(16#cc#)) OR
 					(reg_q1452 AND symb_decoder(16#11#)) OR
 					(reg_q1452 AND symb_decoder(16#b2#)) OR
 					(reg_q1452 AND symb_decoder(16#87#)) OR
 					(reg_q1452 AND symb_decoder(16#1d#)) OR
 					(reg_q1452 AND symb_decoder(16#ad#)) OR
 					(reg_q1452 AND symb_decoder(16#df#)) OR
 					(reg_q1452 AND symb_decoder(16#50#)) OR
 					(reg_q1452 AND symb_decoder(16#c5#)) OR
 					(reg_q1452 AND symb_decoder(16#0a#)) OR
 					(reg_q1452 AND symb_decoder(16#f9#)) OR
 					(reg_q1452 AND symb_decoder(16#4b#)) OR
 					(reg_q1452 AND symb_decoder(16#2e#)) OR
 					(reg_q1452 AND symb_decoder(16#56#)) OR
 					(reg_q1452 AND symb_decoder(16#b3#)) OR
 					(reg_q1452 AND symb_decoder(16#3d#)) OR
 					(reg_q1452 AND symb_decoder(16#9f#)) OR
 					(reg_q1452 AND symb_decoder(16#08#)) OR
 					(reg_q1452 AND symb_decoder(16#07#)) OR
 					(reg_q1452 AND symb_decoder(16#3b#)) OR
 					(reg_q1452 AND symb_decoder(16#22#)) OR
 					(reg_q1452 AND symb_decoder(16#23#)) OR
 					(reg_q1452 AND symb_decoder(16#7b#)) OR
 					(reg_q1452 AND symb_decoder(16#9d#)) OR
 					(reg_q1452 AND symb_decoder(16#a8#)) OR
 					(reg_q1452 AND symb_decoder(16#65#)) OR
 					(reg_q1452 AND symb_decoder(16#bf#)) OR
 					(reg_q1452 AND symb_decoder(16#3f#)) OR
 					(reg_q1452 AND symb_decoder(16#32#)) OR
 					(reg_q1452 AND symb_decoder(16#8e#)) OR
 					(reg_q1452 AND symb_decoder(16#d0#)) OR
 					(reg_q1452 AND symb_decoder(16#c6#)) OR
 					(reg_q1452 AND symb_decoder(16#a0#)) OR
 					(reg_q1452 AND symb_decoder(16#4d#)) OR
 					(reg_q1452 AND symb_decoder(16#c1#)) OR
 					(reg_q1452 AND symb_decoder(16#04#)) OR
 					(reg_q1452 AND symb_decoder(16#62#)) OR
 					(reg_q1452 AND symb_decoder(16#a3#)) OR
 					(reg_q1452 AND symb_decoder(16#f7#)) OR
 					(reg_q1452 AND symb_decoder(16#be#)) OR
 					(reg_q1452 AND symb_decoder(16#e8#)) OR
 					(reg_q1452 AND symb_decoder(16#2c#)) OR
 					(reg_q1452 AND symb_decoder(16#b0#)) OR
 					(reg_q1452 AND symb_decoder(16#ba#)) OR
 					(reg_q1452 AND symb_decoder(16#4e#)) OR
 					(reg_q1452 AND symb_decoder(16#64#)) OR
 					(reg_q1452 AND symb_decoder(16#a6#)) OR
 					(reg_q1452 AND symb_decoder(16#68#)) OR
 					(reg_q1452 AND symb_decoder(16#a5#)) OR
 					(reg_q1452 AND symb_decoder(16#aa#)) OR
 					(reg_q1452 AND symb_decoder(16#43#)) OR
 					(reg_q1452 AND symb_decoder(16#b8#)) OR
 					(reg_q1452 AND symb_decoder(16#25#)) OR
 					(reg_q1452 AND symb_decoder(16#b7#)) OR
 					(reg_q1452 AND symb_decoder(16#28#)) OR
 					(reg_q1452 AND symb_decoder(16#98#)) OR
 					(reg_q1452 AND symb_decoder(16#cd#)) OR
 					(reg_q1452 AND symb_decoder(16#54#)) OR
 					(reg_q1452 AND symb_decoder(16#69#)) OR
 					(reg_q1452 AND symb_decoder(16#30#)) OR
 					(reg_q1452 AND symb_decoder(16#bd#)) OR
 					(reg_q1452 AND symb_decoder(16#e3#)) OR
 					(reg_q1452 AND symb_decoder(16#a7#)) OR
 					(reg_q1452 AND symb_decoder(16#19#)) OR
 					(reg_q1452 AND symb_decoder(16#7e#)) OR
 					(reg_q1452 AND symb_decoder(16#78#)) OR
 					(reg_q1452 AND symb_decoder(16#71#)) OR
 					(reg_q1452 AND symb_decoder(16#80#)) OR
 					(reg_q1452 AND symb_decoder(16#e7#)) OR
 					(reg_q1452 AND symb_decoder(16#f1#)) OR
 					(reg_q1452 AND symb_decoder(16#2b#)) OR
 					(reg_q1452 AND symb_decoder(16#76#)) OR
 					(reg_q1452 AND symb_decoder(16#5c#)) OR
 					(reg_q1452 AND symb_decoder(16#57#)) OR
 					(reg_q1452 AND symb_decoder(16#d5#)) OR
 					(reg_q1452 AND symb_decoder(16#44#)) OR
 					(reg_q1452 AND symb_decoder(16#3c#)) OR
 					(reg_q1452 AND symb_decoder(16#c7#)) OR
 					(reg_q1452 AND symb_decoder(16#61#)) OR
 					(reg_q1452 AND symb_decoder(16#97#)) OR
 					(reg_q1452 AND symb_decoder(16#d8#)) OR
 					(reg_q1452 AND symb_decoder(16#d1#)) OR
 					(reg_q1452 AND symb_decoder(16#1b#)) OR
 					(reg_q1452 AND symb_decoder(16#e6#)) OR
 					(reg_q1452 AND symb_decoder(16#af#)) OR
 					(reg_q1452 AND symb_decoder(16#f8#)) OR
 					(reg_q1452 AND symb_decoder(16#da#)) OR
 					(reg_q1452 AND symb_decoder(16#7f#)) OR
 					(reg_q1452 AND symb_decoder(16#1c#)) OR
 					(reg_q1452 AND symb_decoder(16#06#)) OR
 					(reg_q1452 AND symb_decoder(16#ae#)) OR
 					(reg_q1452 AND symb_decoder(16#58#)) OR
 					(reg_q1452 AND symb_decoder(16#47#)) OR
 					(reg_q1452 AND symb_decoder(16#17#)) OR
 					(reg_q1452 AND symb_decoder(16#8c#)) OR
 					(reg_q1452 AND symb_decoder(16#d6#)) OR
 					(reg_q1452 AND symb_decoder(16#09#)) OR
 					(reg_q1452 AND symb_decoder(16#2d#)) OR
 					(reg_q1452 AND symb_decoder(16#ac#)) OR
 					(reg_q1452 AND symb_decoder(16#29#)) OR
 					(reg_q1452 AND symb_decoder(16#3a#)) OR
 					(reg_q1452 AND symb_decoder(16#0d#)) OR
 					(reg_q1452 AND symb_decoder(16#8b#)) OR
 					(reg_q1452 AND symb_decoder(16#27#)) OR
 					(reg_q1452 AND symb_decoder(16#8f#)) OR
 					(reg_q1452 AND symb_decoder(16#c3#)) OR
 					(reg_q1452 AND symb_decoder(16#c9#)) OR
 					(reg_q1452 AND symb_decoder(16#83#)) OR
 					(reg_q1452 AND symb_decoder(16#e5#)) OR
 					(reg_q1452 AND symb_decoder(16#ab#)) OR
 					(reg_q1452 AND symb_decoder(16#37#)) OR
 					(reg_q1452 AND symb_decoder(16#6e#)) OR
 					(reg_q1452 AND symb_decoder(16#90#)) OR
 					(reg_q1452 AND symb_decoder(16#de#)) OR
 					(reg_q1452 AND symb_decoder(16#b5#)) OR
 					(reg_q1452 AND symb_decoder(16#24#)) OR
 					(reg_q1452 AND symb_decoder(16#5a#)) OR
 					(reg_q1452 AND symb_decoder(16#6c#)) OR
 					(reg_q1452 AND symb_decoder(16#f0#)) OR
 					(reg_q1452 AND symb_decoder(16#f5#)) OR
 					(reg_q1452 AND symb_decoder(16#36#)) OR
 					(reg_q1452 AND symb_decoder(16#e1#)) OR
 					(reg_q1452 AND symb_decoder(16#4a#)) OR
 					(reg_q1452 AND symb_decoder(16#e4#)) OR
 					(reg_q1452 AND symb_decoder(16#82#)) OR
 					(reg_q1452 AND symb_decoder(16#ca#)) OR
 					(reg_q1452 AND symb_decoder(16#96#)) OR
 					(reg_q1452 AND symb_decoder(16#b9#)) OR
 					(reg_q1452 AND symb_decoder(16#20#)) OR
 					(reg_q1452 AND symb_decoder(16#15#)) OR
 					(reg_q1452 AND symb_decoder(16#bb#)) OR
 					(reg_q1452 AND symb_decoder(16#5f#)) OR
 					(reg_q1452 AND symb_decoder(16#73#)) OR
 					(reg_q1452 AND symb_decoder(16#21#)) OR
 					(reg_q1452 AND symb_decoder(16#16#)) OR
 					(reg_q1452 AND symb_decoder(16#59#)) OR
 					(reg_q1452 AND symb_decoder(16#ef#)) OR
 					(reg_q1452 AND symb_decoder(16#ed#)) OR
 					(reg_q1452 AND symb_decoder(16#4c#)) OR
 					(reg_q1452 AND symb_decoder(16#c8#)) OR
 					(reg_q1452 AND symb_decoder(16#7d#)) OR
 					(reg_q1452 AND symb_decoder(16#0b#)) OR
 					(reg_q1452 AND symb_decoder(16#51#)) OR
 					(reg_q1452 AND symb_decoder(16#12#)) OR
 					(reg_q1452 AND symb_decoder(16#2a#)) OR
 					(reg_q1452 AND symb_decoder(16#0c#)) OR
 					(reg_q1452 AND symb_decoder(16#5d#)) OR
 					(reg_q1452 AND symb_decoder(16#42#)) OR
 					(reg_q1452 AND symb_decoder(16#95#)) OR
 					(reg_q1452 AND symb_decoder(16#c2#)) OR
 					(reg_q1452 AND symb_decoder(16#31#)) OR
 					(reg_q1452 AND symb_decoder(16#52#)) OR
 					(reg_q1452 AND symb_decoder(16#92#)) OR
 					(reg_q1452 AND symb_decoder(16#02#)) OR
 					(reg_q1452 AND symb_decoder(16#91#)) OR
 					(reg_q1452 AND symb_decoder(16#a2#)) OR
 					(reg_q1452 AND symb_decoder(16#d4#)) OR
 					(reg_q1452 AND symb_decoder(16#b6#)) OR
 					(reg_q1452 AND symb_decoder(16#41#)) OR
 					(reg_q1452 AND symb_decoder(16#93#)) OR
 					(reg_q1452 AND symb_decoder(16#6f#)) OR
 					(reg_q1452 AND symb_decoder(16#f3#)) OR
 					(reg_q1452 AND symb_decoder(16#89#)) OR
 					(reg_q1452 AND symb_decoder(16#bc#)) OR
 					(reg_q1452 AND symb_decoder(16#0f#)) OR
 					(reg_q1452 AND symb_decoder(16#67#)) OR
 					(reg_q1452 AND symb_decoder(16#13#)) OR
 					(reg_q1452 AND symb_decoder(16#26#)) OR
 					(reg_q1452 AND symb_decoder(16#d2#)) OR
 					(reg_q1452 AND symb_decoder(16#10#)) OR
 					(reg_q1452 AND symb_decoder(16#33#)) OR
 					(reg_q1452 AND symb_decoder(16#a4#)) OR
 					(reg_q1452 AND symb_decoder(16#72#)) OR
 					(reg_q1452 AND symb_decoder(16#c0#)) OR
 					(reg_q1452 AND symb_decoder(16#1f#)) OR
 					(reg_q1452 AND symb_decoder(16#34#)) OR
 					(reg_q1452 AND symb_decoder(16#ea#)) OR
 					(reg_q1452 AND symb_decoder(16#60#)) OR
 					(reg_q1452 AND symb_decoder(16#ff#)) OR
 					(reg_q1452 AND symb_decoder(16#f2#)) OR
 					(reg_q1452 AND symb_decoder(16#9a#)) OR
 					(reg_q1452 AND symb_decoder(16#38#)) OR
 					(reg_q1452 AND symb_decoder(16#8a#)) OR
 					(reg_q1452 AND symb_decoder(16#86#)) OR
 					(reg_q1452 AND symb_decoder(16#05#)) OR
 					(reg_q1452 AND symb_decoder(16#d3#)) OR
 					(reg_q1452 AND symb_decoder(16#81#)) OR
 					(reg_q1452 AND symb_decoder(16#b1#)) OR
 					(reg_q1452 AND symb_decoder(16#94#)) OR
 					(reg_q1452 AND symb_decoder(16#dc#)) OR
 					(reg_q1452 AND symb_decoder(16#e2#)) OR
 					(reg_q1452 AND symb_decoder(16#00#)) OR
 					(reg_q1452 AND symb_decoder(16#db#)) OR
 					(reg_q1452 AND symb_decoder(16#8d#)) OR
 					(reg_q1452 AND symb_decoder(16#66#)) OR
 					(reg_q1452 AND symb_decoder(16#1e#)) OR
 					(reg_q1452 AND symb_decoder(16#eb#)) OR
 					(reg_q1452 AND symb_decoder(16#01#)) OR
 					(reg_q1452 AND symb_decoder(16#55#)) OR
 					(reg_q1452 AND symb_decoder(16#18#)) OR
 					(reg_q1452 AND symb_decoder(16#99#)) OR
 					(reg_q1452 AND symb_decoder(16#48#)) OR
 					(reg_q1452 AND symb_decoder(16#46#)) OR
 					(reg_q1452 AND symb_decoder(16#d7#)) OR
 					(reg_q1452 AND symb_decoder(16#fe#)) OR
 					(reg_q1452 AND symb_decoder(16#0e#));
reg_fullgraph0_init <= "01";

reg_fullgraph0_sel <= "00" & reg_q1452_in & reg_q2695_in;

	--coder fullgraph0
with reg_fullgraph0_sel select
reg_fullgraph0_in <=
	"01" when "0001",
	"10" when "0010",
	"00" when others;
 --end coder

	p_reg_fullgraph0: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph0 <= reg_fullgraph0_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph0 <= reg_fullgraph0_init;
        else
          reg_fullgraph0 <= reg_fullgraph0_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph0

		reg_q2695 <= '1' when reg_fullgraph0 = "01" else '0'; 
		reg_q1452 <= '1' when reg_fullgraph0 = "10" else '0'; 
--end decoder 

reg_q1826_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1826 AND symb_decoder(16#23#)) OR
 					(reg_q1826 AND symb_decoder(16#e8#)) OR
 					(reg_q1826 AND symb_decoder(16#39#)) OR
 					(reg_q1826 AND symb_decoder(16#fa#)) OR
 					(reg_q1826 AND symb_decoder(16#57#)) OR
 					(reg_q1826 AND symb_decoder(16#21#)) OR
 					(reg_q1826 AND symb_decoder(16#e6#)) OR
 					(reg_q1826 AND symb_decoder(16#3b#)) OR
 					(reg_q1826 AND symb_decoder(16#9e#)) OR
 					(reg_q1826 AND symb_decoder(16#fc#)) OR
 					(reg_q1826 AND symb_decoder(16#56#)) OR
 					(reg_q1826 AND symb_decoder(16#95#)) OR
 					(reg_q1826 AND symb_decoder(16#f5#)) OR
 					(reg_q1826 AND symb_decoder(16#0a#)) OR
 					(reg_q1826 AND symb_decoder(16#26#)) OR
 					(reg_q1826 AND symb_decoder(16#c0#)) OR
 					(reg_q1826 AND symb_decoder(16#4e#)) OR
 					(reg_q1826 AND symb_decoder(16#8e#)) OR
 					(reg_q1826 AND symb_decoder(16#1a#)) OR
 					(reg_q1826 AND symb_decoder(16#53#)) OR
 					(reg_q1826 AND symb_decoder(16#25#)) OR
 					(reg_q1826 AND symb_decoder(16#17#)) OR
 					(reg_q1826 AND symb_decoder(16#bd#)) OR
 					(reg_q1826 AND symb_decoder(16#41#)) OR
 					(reg_q1826 AND symb_decoder(16#50#)) OR
 					(reg_q1826 AND symb_decoder(16#7e#)) OR
 					(reg_q1826 AND symb_decoder(16#14#)) OR
 					(reg_q1826 AND symb_decoder(16#04#)) OR
 					(reg_q1826 AND symb_decoder(16#31#)) OR
 					(reg_q1826 AND symb_decoder(16#70#)) OR
 					(reg_q1826 AND symb_decoder(16#2f#)) OR
 					(reg_q1826 AND symb_decoder(16#3a#)) OR
 					(reg_q1826 AND symb_decoder(16#e2#)) OR
 					(reg_q1826 AND symb_decoder(16#a4#)) OR
 					(reg_q1826 AND symb_decoder(16#c2#)) OR
 					(reg_q1826 AND symb_decoder(16#63#)) OR
 					(reg_q1826 AND symb_decoder(16#08#)) OR
 					(reg_q1826 AND symb_decoder(16#30#)) OR
 					(reg_q1826 AND symb_decoder(16#16#)) OR
 					(reg_q1826 AND symb_decoder(16#4a#)) OR
 					(reg_q1826 AND symb_decoder(16#d3#)) OR
 					(reg_q1826 AND symb_decoder(16#72#)) OR
 					(reg_q1826 AND symb_decoder(16#fe#)) OR
 					(reg_q1826 AND symb_decoder(16#d4#)) OR
 					(reg_q1826 AND symb_decoder(16#6c#)) OR
 					(reg_q1826 AND symb_decoder(16#3f#)) OR
 					(reg_q1826 AND symb_decoder(16#db#)) OR
 					(reg_q1826 AND symb_decoder(16#b7#)) OR
 					(reg_q1826 AND symb_decoder(16#e4#)) OR
 					(reg_q1826 AND symb_decoder(16#78#)) OR
 					(reg_q1826 AND symb_decoder(16#42#)) OR
 					(reg_q1826 AND symb_decoder(16#dd#)) OR
 					(reg_q1826 AND symb_decoder(16#5a#)) OR
 					(reg_q1826 AND symb_decoder(16#b9#)) OR
 					(reg_q1826 AND symb_decoder(16#00#)) OR
 					(reg_q1826 AND symb_decoder(16#d5#)) OR
 					(reg_q1826 AND symb_decoder(16#15#)) OR
 					(reg_q1826 AND symb_decoder(16#da#)) OR
 					(reg_q1826 AND symb_decoder(16#2b#)) OR
 					(reg_q1826 AND symb_decoder(16#49#)) OR
 					(reg_q1826 AND symb_decoder(16#84#)) OR
 					(reg_q1826 AND symb_decoder(16#40#)) OR
 					(reg_q1826 AND symb_decoder(16#47#)) OR
 					(reg_q1826 AND symb_decoder(16#be#)) OR
 					(reg_q1826 AND symb_decoder(16#fd#)) OR
 					(reg_q1826 AND symb_decoder(16#dc#)) OR
 					(reg_q1826 AND symb_decoder(16#f0#)) OR
 					(reg_q1826 AND symb_decoder(16#81#)) OR
 					(reg_q1826 AND symb_decoder(16#f6#)) OR
 					(reg_q1826 AND symb_decoder(16#8b#)) OR
 					(reg_q1826 AND symb_decoder(16#90#)) OR
 					(reg_q1826 AND symb_decoder(16#e5#)) OR
 					(reg_q1826 AND symb_decoder(16#b2#)) OR
 					(reg_q1826 AND symb_decoder(16#9c#)) OR
 					(reg_q1826 AND symb_decoder(16#f4#)) OR
 					(reg_q1826 AND symb_decoder(16#ca#)) OR
 					(reg_q1826 AND symb_decoder(16#9b#)) OR
 					(reg_q1826 AND symb_decoder(16#6a#)) OR
 					(reg_q1826 AND symb_decoder(16#2e#)) OR
 					(reg_q1826 AND symb_decoder(16#d2#)) OR
 					(reg_q1826 AND symb_decoder(16#f7#)) OR
 					(reg_q1826 AND symb_decoder(16#85#)) OR
 					(reg_q1826 AND symb_decoder(16#aa#)) OR
 					(reg_q1826 AND symb_decoder(16#73#)) OR
 					(reg_q1826 AND symb_decoder(16#3c#)) OR
 					(reg_q1826 AND symb_decoder(16#1f#)) OR
 					(reg_q1826 AND symb_decoder(16#0f#)) OR
 					(reg_q1826 AND symb_decoder(16#97#)) OR
 					(reg_q1826 AND symb_decoder(16#ab#)) OR
 					(reg_q1826 AND symb_decoder(16#37#)) OR
 					(reg_q1826 AND symb_decoder(16#d9#)) OR
 					(reg_q1826 AND symb_decoder(16#5f#)) OR
 					(reg_q1826 AND symb_decoder(16#ae#)) OR
 					(reg_q1826 AND symb_decoder(16#5c#)) OR
 					(reg_q1826 AND symb_decoder(16#58#)) OR
 					(reg_q1826 AND symb_decoder(16#eb#)) OR
 					(reg_q1826 AND symb_decoder(16#12#)) OR
 					(reg_q1826 AND symb_decoder(16#c6#)) OR
 					(reg_q1826 AND symb_decoder(16#2c#)) OR
 					(reg_q1826 AND symb_decoder(16#7d#)) OR
 					(reg_q1826 AND symb_decoder(16#54#)) OR
 					(reg_q1826 AND symb_decoder(16#cd#)) OR
 					(reg_q1826 AND symb_decoder(16#ea#)) OR
 					(reg_q1826 AND symb_decoder(16#94#)) OR
 					(reg_q1826 AND symb_decoder(16#5d#)) OR
 					(reg_q1826 AND symb_decoder(16#d7#)) OR
 					(reg_q1826 AND symb_decoder(16#20#)) OR
 					(reg_q1826 AND symb_decoder(16#10#)) OR
 					(reg_q1826 AND symb_decoder(16#5e#)) OR
 					(reg_q1826 AND symb_decoder(16#8a#)) OR
 					(reg_q1826 AND symb_decoder(16#a7#)) OR
 					(reg_q1826 AND symb_decoder(16#36#)) OR
 					(reg_q1826 AND symb_decoder(16#1e#)) OR
 					(reg_q1826 AND symb_decoder(16#65#)) OR
 					(reg_q1826 AND symb_decoder(16#bf#)) OR
 					(reg_q1826 AND symb_decoder(16#06#)) OR
 					(reg_q1826 AND symb_decoder(16#e0#)) OR
 					(reg_q1826 AND symb_decoder(16#ad#)) OR
 					(reg_q1826 AND symb_decoder(16#e1#)) OR
 					(reg_q1826 AND symb_decoder(16#fb#)) OR
 					(reg_q1826 AND symb_decoder(16#3d#)) OR
 					(reg_q1826 AND symb_decoder(16#f3#)) OR
 					(reg_q1826 AND symb_decoder(16#24#)) OR
 					(reg_q1826 AND symb_decoder(16#ed#)) OR
 					(reg_q1826 AND symb_decoder(16#c1#)) OR
 					(reg_q1826 AND symb_decoder(16#0c#)) OR
 					(reg_q1826 AND symb_decoder(16#ac#)) OR
 					(reg_q1826 AND symb_decoder(16#1c#)) OR
 					(reg_q1826 AND symb_decoder(16#b4#)) OR
 					(reg_q1826 AND symb_decoder(16#c4#)) OR
 					(reg_q1826 AND symb_decoder(16#e3#)) OR
 					(reg_q1826 AND symb_decoder(16#b6#)) OR
 					(reg_q1826 AND symb_decoder(16#52#)) OR
 					(reg_q1826 AND symb_decoder(16#a2#)) OR
 					(reg_q1826 AND symb_decoder(16#ff#)) OR
 					(reg_q1826 AND symb_decoder(16#2d#)) OR
 					(reg_q1826 AND symb_decoder(16#77#)) OR
 					(reg_q1826 AND symb_decoder(16#9d#)) OR
 					(reg_q1826 AND symb_decoder(16#6e#)) OR
 					(reg_q1826 AND symb_decoder(16#cc#)) OR
 					(reg_q1826 AND symb_decoder(16#a6#)) OR
 					(reg_q1826 AND symb_decoder(16#18#)) OR
 					(reg_q1826 AND symb_decoder(16#d0#)) OR
 					(reg_q1826 AND symb_decoder(16#7f#)) OR
 					(reg_q1826 AND symb_decoder(16#87#)) OR
 					(reg_q1826 AND symb_decoder(16#9a#)) OR
 					(reg_q1826 AND symb_decoder(16#de#)) OR
 					(reg_q1826 AND symb_decoder(16#59#)) OR
 					(reg_q1826 AND symb_decoder(16#5b#)) OR
 					(reg_q1826 AND symb_decoder(16#1d#)) OR
 					(reg_q1826 AND symb_decoder(16#bb#)) OR
 					(reg_q1826 AND symb_decoder(16#7c#)) OR
 					(reg_q1826 AND symb_decoder(16#34#)) OR
 					(reg_q1826 AND symb_decoder(16#7a#)) OR
 					(reg_q1826 AND symb_decoder(16#4d#)) OR
 					(reg_q1826 AND symb_decoder(16#98#)) OR
 					(reg_q1826 AND symb_decoder(16#91#)) OR
 					(reg_q1826 AND symb_decoder(16#b5#)) OR
 					(reg_q1826 AND symb_decoder(16#df#)) OR
 					(reg_q1826 AND symb_decoder(16#b1#)) OR
 					(reg_q1826 AND symb_decoder(16#f9#)) OR
 					(reg_q1826 AND symb_decoder(16#b3#)) OR
 					(reg_q1826 AND symb_decoder(16#69#)) OR
 					(reg_q1826 AND symb_decoder(16#19#)) OR
 					(reg_q1826 AND symb_decoder(16#b8#)) OR
 					(reg_q1826 AND symb_decoder(16#01#)) OR
 					(reg_q1826 AND symb_decoder(16#11#)) OR
 					(reg_q1826 AND symb_decoder(16#46#)) OR
 					(reg_q1826 AND symb_decoder(16#c9#)) OR
 					(reg_q1826 AND symb_decoder(16#8d#)) OR
 					(reg_q1826 AND symb_decoder(16#ec#)) OR
 					(reg_q1826 AND symb_decoder(16#74#)) OR
 					(reg_q1826 AND symb_decoder(16#e9#)) OR
 					(reg_q1826 AND symb_decoder(16#79#)) OR
 					(reg_q1826 AND symb_decoder(16#22#)) OR
 					(reg_q1826 AND symb_decoder(16#55#)) OR
 					(reg_q1826 AND symb_decoder(16#f2#)) OR
 					(reg_q1826 AND symb_decoder(16#44#)) OR
 					(reg_q1826 AND symb_decoder(16#13#)) OR
 					(reg_q1826 AND symb_decoder(16#51#)) OR
 					(reg_q1826 AND symb_decoder(16#d1#)) OR
 					(reg_q1826 AND symb_decoder(16#7b#)) OR
 					(reg_q1826 AND symb_decoder(16#93#)) OR
 					(reg_q1826 AND symb_decoder(16#43#)) OR
 					(reg_q1826 AND symb_decoder(16#45#)) OR
 					(reg_q1826 AND symb_decoder(16#76#)) OR
 					(reg_q1826 AND symb_decoder(16#cb#)) OR
 					(reg_q1826 AND symb_decoder(16#6b#)) OR
 					(reg_q1826 AND symb_decoder(16#33#)) OR
 					(reg_q1826 AND symb_decoder(16#4b#)) OR
 					(reg_q1826 AND symb_decoder(16#1b#)) OR
 					(reg_q1826 AND symb_decoder(16#d6#)) OR
 					(reg_q1826 AND symb_decoder(16#c5#)) OR
 					(reg_q1826 AND symb_decoder(16#0d#)) OR
 					(reg_q1826 AND symb_decoder(16#03#)) OR
 					(reg_q1826 AND symb_decoder(16#61#)) OR
 					(reg_q1826 AND symb_decoder(16#38#)) OR
 					(reg_q1826 AND symb_decoder(16#3e#)) OR
 					(reg_q1826 AND symb_decoder(16#89#)) OR
 					(reg_q1826 AND symb_decoder(16#71#)) OR
 					(reg_q1826 AND symb_decoder(16#99#)) OR
 					(reg_q1826 AND symb_decoder(16#32#)) OR
 					(reg_q1826 AND symb_decoder(16#29#)) OR
 					(reg_q1826 AND symb_decoder(16#6f#)) OR
 					(reg_q1826 AND symb_decoder(16#ce#)) OR
 					(reg_q1826 AND symb_decoder(16#35#)) OR
 					(reg_q1826 AND symb_decoder(16#67#)) OR
 					(reg_q1826 AND symb_decoder(16#a0#)) OR
 					(reg_q1826 AND symb_decoder(16#a5#)) OR
 					(reg_q1826 AND symb_decoder(16#f1#)) OR
 					(reg_q1826 AND symb_decoder(16#c7#)) OR
 					(reg_q1826 AND symb_decoder(16#f8#)) OR
 					(reg_q1826 AND symb_decoder(16#8f#)) OR
 					(reg_q1826 AND symb_decoder(16#82#)) OR
 					(reg_q1826 AND symb_decoder(16#92#)) OR
 					(reg_q1826 AND symb_decoder(16#83#)) OR
 					(reg_q1826 AND symb_decoder(16#6d#)) OR
 					(reg_q1826 AND symb_decoder(16#b0#)) OR
 					(reg_q1826 AND symb_decoder(16#80#)) OR
 					(reg_q1826 AND symb_decoder(16#07#)) OR
 					(reg_q1826 AND symb_decoder(16#ee#)) OR
 					(reg_q1826 AND symb_decoder(16#0b#)) OR
 					(reg_q1826 AND symb_decoder(16#a3#)) OR
 					(reg_q1826 AND symb_decoder(16#af#)) OR
 					(reg_q1826 AND symb_decoder(16#8c#)) OR
 					(reg_q1826 AND symb_decoder(16#e7#)) OR
 					(reg_q1826 AND symb_decoder(16#ef#)) OR
 					(reg_q1826 AND symb_decoder(16#ba#)) OR
 					(reg_q1826 AND symb_decoder(16#75#)) OR
 					(reg_q1826 AND symb_decoder(16#64#)) OR
 					(reg_q1826 AND symb_decoder(16#9f#)) OR
 					(reg_q1826 AND symb_decoder(16#86#)) OR
 					(reg_q1826 AND symb_decoder(16#a1#)) OR
 					(reg_q1826 AND symb_decoder(16#62#)) OR
 					(reg_q1826 AND symb_decoder(16#02#)) OR
 					(reg_q1826 AND symb_decoder(16#09#)) OR
 					(reg_q1826 AND symb_decoder(16#96#)) OR
 					(reg_q1826 AND symb_decoder(16#c3#)) OR
 					(reg_q1826 AND symb_decoder(16#4f#)) OR
 					(reg_q1826 AND symb_decoder(16#68#)) OR
 					(reg_q1826 AND symb_decoder(16#05#)) OR
 					(reg_q1826 AND symb_decoder(16#60#)) OR
 					(reg_q1826 AND symb_decoder(16#a8#)) OR
 					(reg_q1826 AND symb_decoder(16#88#)) OR
 					(reg_q1826 AND symb_decoder(16#4c#)) OR
 					(reg_q1826 AND symb_decoder(16#48#)) OR
 					(reg_q1826 AND symb_decoder(16#2a#)) OR
 					(reg_q1826 AND symb_decoder(16#28#)) OR
 					(reg_q1826 AND symb_decoder(16#27#)) OR
 					(reg_q1826 AND symb_decoder(16#66#)) OR
 					(reg_q1826 AND symb_decoder(16#cf#)) OR
 					(reg_q1826 AND symb_decoder(16#a9#)) OR
 					(reg_q1826 AND symb_decoder(16#d8#)) OR
 					(reg_q1826 AND symb_decoder(16#c8#)) OR
 					(reg_q1826 AND symb_decoder(16#bc#)) OR
 					(reg_q1826 AND symb_decoder(16#0e#));
reg_q1826_init <= '0' ;
	p_reg_q1826: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1826 <= reg_q1826_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1826 <= reg_q1826_init;
        else
          reg_q1826 <= reg_q1826_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph2

reg_q1139_in <= (reg_q1139 AND symb_decoder(16#36#)) OR
 					(reg_q1139 AND symb_decoder(16#32#)) OR
 					(reg_q1139 AND symb_decoder(16#38#)) OR
 					(reg_q1139 AND symb_decoder(16#39#)) OR
 					(reg_q1139 AND symb_decoder(16#31#)) OR
 					(reg_q1139 AND symb_decoder(16#34#)) OR
 					(reg_q1139 AND symb_decoder(16#37#)) OR
 					(reg_q1139 AND symb_decoder(16#35#)) OR
 					(reg_q1139 AND symb_decoder(16#30#)) OR
 					(reg_q1139 AND symb_decoder(16#33#)) OR
 					(reg_q1137 AND symb_decoder(16#37#)) OR
 					(reg_q1137 AND symb_decoder(16#35#)) OR
 					(reg_q1137 AND symb_decoder(16#39#)) OR
 					(reg_q1137 AND symb_decoder(16#30#)) OR
 					(reg_q1137 AND symb_decoder(16#33#)) OR
 					(reg_q1137 AND symb_decoder(16#31#)) OR
 					(reg_q1137 AND symb_decoder(16#34#)) OR
 					(reg_q1137 AND symb_decoder(16#32#)) OR
 					(reg_q1137 AND symb_decoder(16#38#)) OR
 					(reg_q1137 AND symb_decoder(16#36#));
reg_q828_in <= (reg_q826 AND symb_decoder(16#5e#));
reg_q848_in <= (reg_q828 AND symb_decoder(16#b6#)) OR
 					(reg_q828 AND symb_decoder(16#1d#)) OR
 					(reg_q828 AND symb_decoder(16#6f#)) OR
 					(reg_q828 AND symb_decoder(16#b1#)) OR
 					(reg_q828 AND symb_decoder(16#53#)) OR
 					(reg_q828 AND symb_decoder(16#8e#)) OR
 					(reg_q828 AND symb_decoder(16#56#)) OR
 					(reg_q828 AND symb_decoder(16#d4#)) OR
 					(reg_q828 AND symb_decoder(16#27#)) OR
 					(reg_q828 AND symb_decoder(16#d0#)) OR
 					(reg_q828 AND symb_decoder(16#61#)) OR
 					(reg_q828 AND symb_decoder(16#20#)) OR
 					(reg_q828 AND symb_decoder(16#59#)) OR
 					(reg_q828 AND symb_decoder(16#a4#)) OR
 					(reg_q828 AND symb_decoder(16#c7#)) OR
 					(reg_q828 AND symb_decoder(16#63#)) OR
 					(reg_q828 AND symb_decoder(16#2c#)) OR
 					(reg_q828 AND symb_decoder(16#87#)) OR
 					(reg_q828 AND symb_decoder(16#bd#)) OR
 					(reg_q828 AND symb_decoder(16#36#)) OR
 					(reg_q828 AND symb_decoder(16#05#)) OR
 					(reg_q828 AND symb_decoder(16#5f#)) OR
 					(reg_q828 AND symb_decoder(16#24#)) OR
 					(reg_q828 AND symb_decoder(16#84#)) OR
 					(reg_q828 AND symb_decoder(16#34#)) OR
 					(reg_q828 AND symb_decoder(16#b5#)) OR
 					(reg_q828 AND symb_decoder(16#9f#)) OR
 					(reg_q828 AND symb_decoder(16#37#)) OR
 					(reg_q828 AND symb_decoder(16#22#)) OR
 					(reg_q828 AND symb_decoder(16#e1#)) OR
 					(reg_q828 AND symb_decoder(16#70#)) OR
 					(reg_q828 AND symb_decoder(16#55#)) OR
 					(reg_q828 AND symb_decoder(16#c2#)) OR
 					(reg_q828 AND symb_decoder(16#c5#)) OR
 					(reg_q828 AND symb_decoder(16#7a#)) OR
 					(reg_q828 AND symb_decoder(16#ee#)) OR
 					(reg_q828 AND symb_decoder(16#67#)) OR
 					(reg_q828 AND symb_decoder(16#35#)) OR
 					(reg_q828 AND symb_decoder(16#bc#)) OR
 					(reg_q828 AND symb_decoder(16#85#)) OR
 					(reg_q828 AND symb_decoder(16#f5#)) OR
 					(reg_q828 AND symb_decoder(16#5e#)) OR
 					(reg_q828 AND symb_decoder(16#38#)) OR
 					(reg_q828 AND symb_decoder(16#fd#)) OR
 					(reg_q828 AND symb_decoder(16#df#)) OR
 					(reg_q828 AND symb_decoder(16#4c#)) OR
 					(reg_q828 AND symb_decoder(16#d2#)) OR
 					(reg_q828 AND symb_decoder(16#ed#)) OR
 					(reg_q828 AND symb_decoder(16#83#)) OR
 					(reg_q828 AND symb_decoder(16#57#)) OR
 					(reg_q828 AND symb_decoder(16#4d#)) OR
 					(reg_q828 AND symb_decoder(16#3f#)) OR
 					(reg_q828 AND symb_decoder(16#79#)) OR
 					(reg_q828 AND symb_decoder(16#64#)) OR
 					(reg_q828 AND symb_decoder(16#cb#)) OR
 					(reg_q828 AND symb_decoder(16#25#)) OR
 					(reg_q828 AND symb_decoder(16#95#)) OR
 					(reg_q828 AND symb_decoder(16#92#)) OR
 					(reg_q828 AND symb_decoder(16#6a#)) OR
 					(reg_q828 AND symb_decoder(16#76#)) OR
 					(reg_q828 AND symb_decoder(16#a9#)) OR
 					(reg_q828 AND symb_decoder(16#f9#)) OR
 					(reg_q828 AND symb_decoder(16#21#)) OR
 					(reg_q828 AND symb_decoder(16#5a#)) OR
 					(reg_q828 AND symb_decoder(16#e2#)) OR
 					(reg_q828 AND symb_decoder(16#29#)) OR
 					(reg_q828 AND symb_decoder(16#52#)) OR
 					(reg_q828 AND symb_decoder(16#c0#)) OR
 					(reg_q828 AND symb_decoder(16#10#)) OR
 					(reg_q828 AND symb_decoder(16#8f#)) OR
 					(reg_q828 AND symb_decoder(16#3b#)) OR
 					(reg_q828 AND symb_decoder(16#c6#)) OR
 					(reg_q828 AND symb_decoder(16#9a#)) OR
 					(reg_q828 AND symb_decoder(16#eb#)) OR
 					(reg_q828 AND symb_decoder(16#42#)) OR
 					(reg_q828 AND symb_decoder(16#1f#)) OR
 					(reg_q828 AND symb_decoder(16#2b#)) OR
 					(reg_q828 AND symb_decoder(16#3a#)) OR
 					(reg_q828 AND symb_decoder(16#06#)) OR
 					(reg_q828 AND symb_decoder(16#69#)) OR
 					(reg_q828 AND symb_decoder(16#8d#)) OR
 					(reg_q828 AND symb_decoder(16#90#)) OR
 					(reg_q828 AND symb_decoder(16#13#)) OR
 					(reg_q828 AND symb_decoder(16#d5#)) OR
 					(reg_q828 AND symb_decoder(16#7b#)) OR
 					(reg_q828 AND symb_decoder(16#66#)) OR
 					(reg_q828 AND symb_decoder(16#71#)) OR
 					(reg_q828 AND symb_decoder(16#d9#)) OR
 					(reg_q828 AND symb_decoder(16#39#)) OR
 					(reg_q828 AND symb_decoder(16#a5#)) OR
 					(reg_q828 AND symb_decoder(16#89#)) OR
 					(reg_q828 AND symb_decoder(16#b7#)) OR
 					(reg_q828 AND symb_decoder(16#b3#)) OR
 					(reg_q828 AND symb_decoder(16#82#)) OR
 					(reg_q828 AND symb_decoder(16#e3#)) OR
 					(reg_q828 AND symb_decoder(16#b4#)) OR
 					(reg_q828 AND symb_decoder(16#65#)) OR
 					(reg_q828 AND symb_decoder(16#7e#)) OR
 					(reg_q828 AND symb_decoder(16#c1#)) OR
 					(reg_q828 AND symb_decoder(16#f0#)) OR
 					(reg_q828 AND symb_decoder(16#0f#)) OR
 					(reg_q828 AND symb_decoder(16#86#)) OR
 					(reg_q828 AND symb_decoder(16#f4#)) OR
 					(reg_q828 AND symb_decoder(16#91#)) OR
 					(reg_q828 AND symb_decoder(16#12#)) OR
 					(reg_q828 AND symb_decoder(16#26#)) OR
 					(reg_q828 AND symb_decoder(16#a6#)) OR
 					(reg_q828 AND symb_decoder(16#ec#)) OR
 					(reg_q828 AND symb_decoder(16#5d#)) OR
 					(reg_q828 AND symb_decoder(16#8b#)) OR
 					(reg_q828 AND symb_decoder(16#18#)) OR
 					(reg_q828 AND symb_decoder(16#2a#)) OR
 					(reg_q828 AND symb_decoder(16#5b#)) OR
 					(reg_q828 AND symb_decoder(16#33#)) OR
 					(reg_q828 AND symb_decoder(16#a3#)) OR
 					(reg_q828 AND symb_decoder(16#4a#)) OR
 					(reg_q828 AND symb_decoder(16#9e#)) OR
 					(reg_q828 AND symb_decoder(16#14#)) OR
 					(reg_q828 AND symb_decoder(16#fe#)) OR
 					(reg_q828 AND symb_decoder(16#73#)) OR
 					(reg_q828 AND symb_decoder(16#ae#)) OR
 					(reg_q828 AND symb_decoder(16#88#)) OR
 					(reg_q828 AND symb_decoder(16#de#)) OR
 					(reg_q828 AND symb_decoder(16#03#)) OR
 					(reg_q828 AND symb_decoder(16#e5#)) OR
 					(reg_q828 AND symb_decoder(16#49#)) OR
 					(reg_q828 AND symb_decoder(16#a8#)) OR
 					(reg_q828 AND symb_decoder(16#44#)) OR
 					(reg_q828 AND symb_decoder(16#b0#)) OR
 					(reg_q828 AND symb_decoder(16#6c#)) OR
 					(reg_q828 AND symb_decoder(16#d3#)) OR
 					(reg_q828 AND symb_decoder(16#b2#)) OR
 					(reg_q828 AND symb_decoder(16#1b#)) OR
 					(reg_q828 AND symb_decoder(16#d7#)) OR
 					(reg_q828 AND symb_decoder(16#3d#)) OR
 					(reg_q828 AND symb_decoder(16#0b#)) OR
 					(reg_q828 AND symb_decoder(16#62#)) OR
 					(reg_q828 AND symb_decoder(16#a7#)) OR
 					(reg_q828 AND symb_decoder(16#f2#)) OR
 					(reg_q828 AND symb_decoder(16#54#)) OR
 					(reg_q828 AND symb_decoder(16#cd#)) OR
 					(reg_q828 AND symb_decoder(16#9b#)) OR
 					(reg_q828 AND symb_decoder(16#d6#)) OR
 					(reg_q828 AND symb_decoder(16#68#)) OR
 					(reg_q828 AND symb_decoder(16#e0#)) OR
 					(reg_q828 AND symb_decoder(16#c9#)) OR
 					(reg_q828 AND symb_decoder(16#d8#)) OR
 					(reg_q828 AND symb_decoder(16#e6#)) OR
 					(reg_q828 AND symb_decoder(16#b8#)) OR
 					(reg_q828 AND symb_decoder(16#fa#)) OR
 					(reg_q828 AND symb_decoder(16#6e#)) OR
 					(reg_q828 AND symb_decoder(16#cf#)) OR
 					(reg_q828 AND symb_decoder(16#ab#)) OR
 					(reg_q828 AND symb_decoder(16#19#)) OR
 					(reg_q828 AND symb_decoder(16#7d#)) OR
 					(reg_q828 AND symb_decoder(16#97#)) OR
 					(reg_q828 AND symb_decoder(16#17#)) OR
 					(reg_q828 AND symb_decoder(16#28#)) OR
 					(reg_q828 AND symb_decoder(16#32#)) OR
 					(reg_q828 AND symb_decoder(16#93#)) OR
 					(reg_q828 AND symb_decoder(16#1c#)) OR
 					(reg_q828 AND symb_decoder(16#07#)) OR
 					(reg_q828 AND symb_decoder(16#ad#)) OR
 					(reg_q828 AND symb_decoder(16#1a#)) OR
 					(reg_q828 AND symb_decoder(16#9c#)) OR
 					(reg_q828 AND symb_decoder(16#e9#)) OR
 					(reg_q828 AND symb_decoder(16#5c#)) OR
 					(reg_q828 AND symb_decoder(16#e8#)) OR
 					(reg_q828 AND symb_decoder(16#75#)) OR
 					(reg_q828 AND symb_decoder(16#7f#)) OR
 					(reg_q828 AND symb_decoder(16#4e#)) OR
 					(reg_q828 AND symb_decoder(16#96#)) OR
 					(reg_q828 AND symb_decoder(16#94#)) OR
 					(reg_q828 AND symb_decoder(16#81#)) OR
 					(reg_q828 AND symb_decoder(16#c4#)) OR
 					(reg_q828 AND symb_decoder(16#e7#)) OR
 					(reg_q828 AND symb_decoder(16#f6#)) OR
 					(reg_q828 AND symb_decoder(16#31#)) OR
 					(reg_q828 AND symb_decoder(16#0c#)) OR
 					(reg_q828 AND symb_decoder(16#99#)) OR
 					(reg_q828 AND symb_decoder(16#6b#)) OR
 					(reg_q828 AND symb_decoder(16#ac#)) OR
 					(reg_q828 AND symb_decoder(16#80#)) OR
 					(reg_q828 AND symb_decoder(16#a1#)) OR
 					(reg_q828 AND symb_decoder(16#da#)) OR
 					(reg_q828 AND symb_decoder(16#2d#)) OR
 					(reg_q828 AND symb_decoder(16#1e#)) OR
 					(reg_q828 AND symb_decoder(16#78#)) OR
 					(reg_q828 AND symb_decoder(16#cc#)) OR
 					(reg_q828 AND symb_decoder(16#f8#)) OR
 					(reg_q828 AND symb_decoder(16#74#)) OR
 					(reg_q828 AND symb_decoder(16#b9#)) OR
 					(reg_q828 AND symb_decoder(16#f3#)) OR
 					(reg_q828 AND symb_decoder(16#af#)) OR
 					(reg_q828 AND symb_decoder(16#fc#)) OR
 					(reg_q828 AND symb_decoder(16#98#)) OR
 					(reg_q828 AND symb_decoder(16#02#)) OR
 					(reg_q828 AND symb_decoder(16#dc#)) OR
 					(reg_q828 AND symb_decoder(16#46#)) OR
 					(reg_q828 AND symb_decoder(16#01#)) OR
 					(reg_q828 AND symb_decoder(16#60#)) OR
 					(reg_q828 AND symb_decoder(16#a0#)) OR
 					(reg_q828 AND symb_decoder(16#a2#)) OR
 					(reg_q828 AND symb_decoder(16#47#)) OR
 					(reg_q828 AND symb_decoder(16#f1#)) OR
 					(reg_q828 AND symb_decoder(16#2e#)) OR
 					(reg_q828 AND symb_decoder(16#bf#)) OR
 					(reg_q828 AND symb_decoder(16#0e#)) OR
 					(reg_q828 AND symb_decoder(16#08#)) OR
 					(reg_q828 AND symb_decoder(16#e4#)) OR
 					(reg_q828 AND symb_decoder(16#40#)) OR
 					(reg_q828 AND symb_decoder(16#04#)) OR
 					(reg_q828 AND symb_decoder(16#be#)) OR
 					(reg_q828 AND symb_decoder(16#fb#)) OR
 					(reg_q828 AND symb_decoder(16#43#)) OR
 					(reg_q828 AND symb_decoder(16#8a#)) OR
 					(reg_q828 AND symb_decoder(16#00#)) OR
 					(reg_q828 AND symb_decoder(16#41#)) OR
 					(reg_q828 AND symb_decoder(16#7c#)) OR
 					(reg_q828 AND symb_decoder(16#ca#)) OR
 					(reg_q828 AND symb_decoder(16#8c#)) OR
 					(reg_q828 AND symb_decoder(16#2f#)) OR
 					(reg_q828 AND symb_decoder(16#db#)) OR
 					(reg_q828 AND symb_decoder(16#9d#)) OR
 					(reg_q828 AND symb_decoder(16#51#)) OR
 					(reg_q828 AND symb_decoder(16#58#)) OR
 					(reg_q828 AND symb_decoder(16#77#)) OR
 					(reg_q828 AND symb_decoder(16#bb#)) OR
 					(reg_q828 AND symb_decoder(16#c3#)) OR
 					(reg_q828 AND symb_decoder(16#3c#)) OR
 					(reg_q828 AND symb_decoder(16#f7#)) OR
 					(reg_q828 AND symb_decoder(16#45#)) OR
 					(reg_q828 AND symb_decoder(16#50#)) OR
 					(reg_q828 AND symb_decoder(16#aa#)) OR
 					(reg_q828 AND symb_decoder(16#c8#)) OR
 					(reg_q828 AND symb_decoder(16#ba#)) OR
 					(reg_q828 AND symb_decoder(16#d1#)) OR
 					(reg_q828 AND symb_decoder(16#16#)) OR
 					(reg_q828 AND symb_decoder(16#30#)) OR
 					(reg_q828 AND symb_decoder(16#09#)) OR
 					(reg_q828 AND symb_decoder(16#6d#)) OR
 					(reg_q828 AND symb_decoder(16#ff#)) OR
 					(reg_q828 AND symb_decoder(16#48#)) OR
 					(reg_q828 AND symb_decoder(16#72#)) OR
 					(reg_q828 AND symb_decoder(16#23#)) OR
 					(reg_q828 AND symb_decoder(16#15#)) OR
 					(reg_q828 AND symb_decoder(16#11#)) OR
 					(reg_q828 AND symb_decoder(16#ea#)) OR
 					(reg_q828 AND symb_decoder(16#4f#)) OR
 					(reg_q828 AND symb_decoder(16#dd#)) OR
 					(reg_q828 AND symb_decoder(16#ce#)) OR
 					(reg_q828 AND symb_decoder(16#4b#)) OR
 					(reg_q828 AND symb_decoder(16#ef#)) OR
 					(reg_q828 AND symb_decoder(16#3e#)) OR
 					(reg_q848 AND symb_decoder(16#ce#)) OR
 					(reg_q848 AND symb_decoder(16#32#)) OR
 					(reg_q848 AND symb_decoder(16#0e#)) OR
 					(reg_q848 AND symb_decoder(16#8b#)) OR
 					(reg_q848 AND symb_decoder(16#e9#)) OR
 					(reg_q848 AND symb_decoder(16#02#)) OR
 					(reg_q848 AND symb_decoder(16#e8#)) OR
 					(reg_q848 AND symb_decoder(16#a8#)) OR
 					(reg_q848 AND symb_decoder(16#85#)) OR
 					(reg_q848 AND symb_decoder(16#a9#)) OR
 					(reg_q848 AND symb_decoder(16#f9#)) OR
 					(reg_q848 AND symb_decoder(16#22#)) OR
 					(reg_q848 AND symb_decoder(16#45#)) OR
 					(reg_q848 AND symb_decoder(16#33#)) OR
 					(reg_q848 AND symb_decoder(16#b8#)) OR
 					(reg_q848 AND symb_decoder(16#83#)) OR
 					(reg_q848 AND symb_decoder(16#08#)) OR
 					(reg_q848 AND symb_decoder(16#c2#)) OR
 					(reg_q848 AND symb_decoder(16#68#)) OR
 					(reg_q848 AND symb_decoder(16#86#)) OR
 					(reg_q848 AND symb_decoder(16#71#)) OR
 					(reg_q848 AND symb_decoder(16#9f#)) OR
 					(reg_q848 AND symb_decoder(16#96#)) OR
 					(reg_q848 AND symb_decoder(16#d0#)) OR
 					(reg_q848 AND symb_decoder(16#53#)) OR
 					(reg_q848 AND symb_decoder(16#2d#)) OR
 					(reg_q848 AND symb_decoder(16#64#)) OR
 					(reg_q848 AND symb_decoder(16#78#)) OR
 					(reg_q848 AND symb_decoder(16#51#)) OR
 					(reg_q848 AND symb_decoder(16#d5#)) OR
 					(reg_q848 AND symb_decoder(16#f2#)) OR
 					(reg_q848 AND symb_decoder(16#3c#)) OR
 					(reg_q848 AND symb_decoder(16#5a#)) OR
 					(reg_q848 AND symb_decoder(16#10#)) OR
 					(reg_q848 AND symb_decoder(16#2e#)) OR
 					(reg_q848 AND symb_decoder(16#4c#)) OR
 					(reg_q848 AND symb_decoder(16#df#)) OR
 					(reg_q848 AND symb_decoder(16#4d#)) OR
 					(reg_q848 AND symb_decoder(16#80#)) OR
 					(reg_q848 AND symb_decoder(16#a3#)) OR
 					(reg_q848 AND symb_decoder(16#18#)) OR
 					(reg_q848 AND symb_decoder(16#d6#)) OR
 					(reg_q848 AND symb_decoder(16#76#)) OR
 					(reg_q848 AND symb_decoder(16#0c#)) OR
 					(reg_q848 AND symb_decoder(16#47#)) OR
 					(reg_q848 AND symb_decoder(16#7d#)) OR
 					(reg_q848 AND symb_decoder(16#cd#)) OR
 					(reg_q848 AND symb_decoder(16#54#)) OR
 					(reg_q848 AND symb_decoder(16#8d#)) OR
 					(reg_q848 AND symb_decoder(16#57#)) OR
 					(reg_q848 AND symb_decoder(16#ed#)) OR
 					(reg_q848 AND symb_decoder(16#bb#)) OR
 					(reg_q848 AND symb_decoder(16#c4#)) OR
 					(reg_q848 AND symb_decoder(16#8f#)) OR
 					(reg_q848 AND symb_decoder(16#aa#)) OR
 					(reg_q848 AND symb_decoder(16#01#)) OR
 					(reg_q848 AND symb_decoder(16#e6#)) OR
 					(reg_q848 AND symb_decoder(16#fa#)) OR
 					(reg_q848 AND symb_decoder(16#15#)) OR
 					(reg_q848 AND symb_decoder(16#6f#)) OR
 					(reg_q848 AND symb_decoder(16#d7#)) OR
 					(reg_q848 AND symb_decoder(16#bd#)) OR
 					(reg_q848 AND symb_decoder(16#e2#)) OR
 					(reg_q848 AND symb_decoder(16#16#)) OR
 					(reg_q848 AND symb_decoder(16#00#)) OR
 					(reg_q848 AND symb_decoder(16#12#)) OR
 					(reg_q848 AND symb_decoder(16#bf#)) OR
 					(reg_q848 AND symb_decoder(16#9d#)) OR
 					(reg_q848 AND symb_decoder(16#bc#)) OR
 					(reg_q848 AND symb_decoder(16#4e#)) OR
 					(reg_q848 AND symb_decoder(16#db#)) OR
 					(reg_q848 AND symb_decoder(16#35#)) OR
 					(reg_q848 AND symb_decoder(16#97#)) OR
 					(reg_q848 AND symb_decoder(16#cb#)) OR
 					(reg_q848 AND symb_decoder(16#59#)) OR
 					(reg_q848 AND symb_decoder(16#f8#)) OR
 					(reg_q848 AND symb_decoder(16#62#)) OR
 					(reg_q848 AND symb_decoder(16#ae#)) OR
 					(reg_q848 AND symb_decoder(16#90#)) OR
 					(reg_q848 AND symb_decoder(16#1d#)) OR
 					(reg_q848 AND symb_decoder(16#ef#)) OR
 					(reg_q848 AND symb_decoder(16#21#)) OR
 					(reg_q848 AND symb_decoder(16#7f#)) OR
 					(reg_q848 AND symb_decoder(16#38#)) OR
 					(reg_q848 AND symb_decoder(16#f4#)) OR
 					(reg_q848 AND symb_decoder(16#30#)) OR
 					(reg_q848 AND symb_decoder(16#65#)) OR
 					(reg_q848 AND symb_decoder(16#73#)) OR
 					(reg_q848 AND symb_decoder(16#5c#)) OR
 					(reg_q848 AND symb_decoder(16#ca#)) OR
 					(reg_q848 AND symb_decoder(16#f3#)) OR
 					(reg_q848 AND symb_decoder(16#da#)) OR
 					(reg_q848 AND symb_decoder(16#ec#)) OR
 					(reg_q848 AND symb_decoder(16#55#)) OR
 					(reg_q848 AND symb_decoder(16#67#)) OR
 					(reg_q848 AND symb_decoder(16#75#)) OR
 					(reg_q848 AND symb_decoder(16#a0#)) OR
 					(reg_q848 AND symb_decoder(16#52#)) OR
 					(reg_q848 AND symb_decoder(16#e5#)) OR
 					(reg_q848 AND symb_decoder(16#fb#)) OR
 					(reg_q848 AND symb_decoder(16#37#)) OR
 					(reg_q848 AND symb_decoder(16#f0#)) OR
 					(reg_q848 AND symb_decoder(16#ee#)) OR
 					(reg_q848 AND symb_decoder(16#a4#)) OR
 					(reg_q848 AND symb_decoder(16#44#)) OR
 					(reg_q848 AND symb_decoder(16#d2#)) OR
 					(reg_q848 AND symb_decoder(16#70#)) OR
 					(reg_q848 AND symb_decoder(16#14#)) OR
 					(reg_q848 AND symb_decoder(16#4b#)) OR
 					(reg_q848 AND symb_decoder(16#6e#)) OR
 					(reg_q848 AND symb_decoder(16#b9#)) OR
 					(reg_q848 AND symb_decoder(16#72#)) OR
 					(reg_q848 AND symb_decoder(16#88#)) OR
 					(reg_q848 AND symb_decoder(16#f6#)) OR
 					(reg_q848 AND symb_decoder(16#99#)) OR
 					(reg_q848 AND symb_decoder(16#ff#)) OR
 					(reg_q848 AND symb_decoder(16#77#)) OR
 					(reg_q848 AND symb_decoder(16#dd#)) OR
 					(reg_q848 AND symb_decoder(16#cf#)) OR
 					(reg_q848 AND symb_decoder(16#63#)) OR
 					(reg_q848 AND symb_decoder(16#c1#)) OR
 					(reg_q848 AND symb_decoder(16#eb#)) OR
 					(reg_q848 AND symb_decoder(16#93#)) OR
 					(reg_q848 AND symb_decoder(16#34#)) OR
 					(reg_q848 AND symb_decoder(16#f5#)) OR
 					(reg_q848 AND symb_decoder(16#ad#)) OR
 					(reg_q848 AND symb_decoder(16#a1#)) OR
 					(reg_q848 AND symb_decoder(16#74#)) OR
 					(reg_q848 AND symb_decoder(16#81#)) OR
 					(reg_q848 AND symb_decoder(16#82#)) OR
 					(reg_q848 AND symb_decoder(16#e7#)) OR
 					(reg_q848 AND symb_decoder(16#e3#)) OR
 					(reg_q848 AND symb_decoder(16#91#)) OR
 					(reg_q848 AND symb_decoder(16#39#)) OR
 					(reg_q848 AND symb_decoder(16#11#)) OR
 					(reg_q848 AND symb_decoder(16#2b#)) OR
 					(reg_q848 AND symb_decoder(16#4f#)) OR
 					(reg_q848 AND symb_decoder(16#27#)) OR
 					(reg_q848 AND symb_decoder(16#94#)) OR
 					(reg_q848 AND symb_decoder(16#1a#)) OR
 					(reg_q848 AND symb_decoder(16#a2#)) OR
 					(reg_q848 AND symb_decoder(16#25#)) OR
 					(reg_q848 AND symb_decoder(16#4a#)) OR
 					(reg_q848 AND symb_decoder(16#6a#)) OR
 					(reg_q848 AND symb_decoder(16#f7#)) OR
 					(reg_q848 AND symb_decoder(16#58#)) OR
 					(reg_q848 AND symb_decoder(16#9c#)) OR
 					(reg_q848 AND symb_decoder(16#0b#)) OR
 					(reg_q848 AND symb_decoder(16#9a#)) OR
 					(reg_q848 AND symb_decoder(16#c3#)) OR
 					(reg_q848 AND symb_decoder(16#5e#)) OR
 					(reg_q848 AND symb_decoder(16#b3#)) OR
 					(reg_q848 AND symb_decoder(16#be#)) OR
 					(reg_q848 AND symb_decoder(16#06#)) OR
 					(reg_q848 AND symb_decoder(16#c7#)) OR
 					(reg_q848 AND symb_decoder(16#5b#)) OR
 					(reg_q848 AND symb_decoder(16#07#)) OR
 					(reg_q848 AND symb_decoder(16#b4#)) OR
 					(reg_q848 AND symb_decoder(16#17#)) OR
 					(reg_q848 AND symb_decoder(16#b2#)) OR
 					(reg_q848 AND symb_decoder(16#7e#)) OR
 					(reg_q848 AND symb_decoder(16#48#)) OR
 					(reg_q848 AND symb_decoder(16#7a#)) OR
 					(reg_q848 AND symb_decoder(16#36#)) OR
 					(reg_q848 AND symb_decoder(16#1c#)) OR
 					(reg_q848 AND symb_decoder(16#1e#)) OR
 					(reg_q848 AND symb_decoder(16#49#)) OR
 					(reg_q848 AND symb_decoder(16#fe#)) OR
 					(reg_q848 AND symb_decoder(16#43#)) OR
 					(reg_q848 AND symb_decoder(16#a7#)) OR
 					(reg_q848 AND symb_decoder(16#3b#)) OR
 					(reg_q848 AND symb_decoder(16#fc#)) OR
 					(reg_q848 AND symb_decoder(16#ea#)) OR
 					(reg_q848 AND symb_decoder(16#26#)) OR
 					(reg_q848 AND symb_decoder(16#24#)) OR
 					(reg_q848 AND symb_decoder(16#19#)) OR
 					(reg_q848 AND symb_decoder(16#d3#)) OR
 					(reg_q848 AND symb_decoder(16#9e#)) OR
 					(reg_q848 AND symb_decoder(16#2a#)) OR
 					(reg_q848 AND symb_decoder(16#c0#)) OR
 					(reg_q848 AND symb_decoder(16#66#)) OR
 					(reg_q848 AND symb_decoder(16#95#)) OR
 					(reg_q848 AND symb_decoder(16#e4#)) OR
 					(reg_q848 AND symb_decoder(16#6b#)) OR
 					(reg_q848 AND symb_decoder(16#60#)) OR
 					(reg_q848 AND symb_decoder(16#c6#)) OR
 					(reg_q848 AND symb_decoder(16#05#)) OR
 					(reg_q848 AND symb_decoder(16#b0#)) OR
 					(reg_q848 AND symb_decoder(16#69#)) OR
 					(reg_q848 AND symb_decoder(16#a5#)) OR
 					(reg_q848 AND symb_decoder(16#d1#)) OR
 					(reg_q848 AND symb_decoder(16#9b#)) OR
 					(reg_q848 AND symb_decoder(16#b7#)) OR
 					(reg_q848 AND symb_decoder(16#de#)) OR
 					(reg_q848 AND symb_decoder(16#5f#)) OR
 					(reg_q848 AND symb_decoder(16#3e#)) OR
 					(reg_q848 AND symb_decoder(16#8c#)) OR
 					(reg_q848 AND symb_decoder(16#1f#)) OR
 					(reg_q848 AND symb_decoder(16#ab#)) OR
 					(reg_q848 AND symb_decoder(16#cc#)) OR
 					(reg_q848 AND symb_decoder(16#0f#)) OR
 					(reg_q848 AND symb_decoder(16#09#)) OR
 					(reg_q848 AND symb_decoder(16#41#)) OR
 					(reg_q848 AND symb_decoder(16#13#)) OR
 					(reg_q848 AND symb_decoder(16#89#)) OR
 					(reg_q848 AND symb_decoder(16#2f#)) OR
 					(reg_q848 AND symb_decoder(16#28#)) OR
 					(reg_q848 AND symb_decoder(16#79#)) OR
 					(reg_q848 AND symb_decoder(16#fd#)) OR
 					(reg_q848 AND symb_decoder(16#e0#)) OR
 					(reg_q848 AND symb_decoder(16#8e#)) OR
 					(reg_q848 AND symb_decoder(16#98#)) OR
 					(reg_q848 AND symb_decoder(16#61#)) OR
 					(reg_q848 AND symb_decoder(16#5d#)) OR
 					(reg_q848 AND symb_decoder(16#b1#)) OR
 					(reg_q848 AND symb_decoder(16#3d#)) OR
 					(reg_q848 AND symb_decoder(16#6c#)) OR
 					(reg_q848 AND symb_decoder(16#b5#)) OR
 					(reg_q848 AND symb_decoder(16#23#)) OR
 					(reg_q848 AND symb_decoder(16#6d#)) OR
 					(reg_q848 AND symb_decoder(16#e1#)) OR
 					(reg_q848 AND symb_decoder(16#46#)) OR
 					(reg_q848 AND symb_decoder(16#40#)) OR
 					(reg_q848 AND symb_decoder(16#42#)) OR
 					(reg_q848 AND symb_decoder(16#dc#)) OR
 					(reg_q848 AND symb_decoder(16#1b#)) OR
 					(reg_q848 AND symb_decoder(16#8a#)) OR
 					(reg_q848 AND symb_decoder(16#31#)) OR
 					(reg_q848 AND symb_decoder(16#3a#)) OR
 					(reg_q848 AND symb_decoder(16#c5#)) OR
 					(reg_q848 AND symb_decoder(16#ba#)) OR
 					(reg_q848 AND symb_decoder(16#56#)) OR
 					(reg_q848 AND symb_decoder(16#b6#)) OR
 					(reg_q848 AND symb_decoder(16#92#)) OR
 					(reg_q848 AND symb_decoder(16#7c#)) OR
 					(reg_q848 AND symb_decoder(16#03#)) OR
 					(reg_q848 AND symb_decoder(16#f1#)) OR
 					(reg_q848 AND symb_decoder(16#7b#)) OR
 					(reg_q848 AND symb_decoder(16#50#)) OR
 					(reg_q848 AND symb_decoder(16#2c#)) OR
 					(reg_q848 AND symb_decoder(16#29#)) OR
 					(reg_q848 AND symb_decoder(16#af#)) OR
 					(reg_q848 AND symb_decoder(16#d9#)) OR
 					(reg_q848 AND symb_decoder(16#84#)) OR
 					(reg_q848 AND symb_decoder(16#04#)) OR
 					(reg_q848 AND symb_decoder(16#3f#)) OR
 					(reg_q848 AND symb_decoder(16#d8#)) OR
 					(reg_q848 AND symb_decoder(16#87#)) OR
 					(reg_q848 AND symb_decoder(16#c9#)) OR
 					(reg_q848 AND symb_decoder(16#c8#)) OR
 					(reg_q848 AND symb_decoder(16#d4#)) OR
 					(reg_q848 AND symb_decoder(16#ac#)) OR
 					(reg_q848 AND symb_decoder(16#a6#)) OR
 					(reg_q848 AND symb_decoder(16#20#));
reg_q2579_in <= (reg_q2579 AND symb_decoder(16#09#)) OR
 					(reg_q2579 AND symb_decoder(16#20#)) OR
 					(reg_q2579 AND symb_decoder(16#0c#)) OR
 					(reg_q2579 AND symb_decoder(16#0d#)) OR
 					(reg_q2579 AND symb_decoder(16#0a#)) OR
 					(reg_q2577 AND symb_decoder(16#0a#)) OR
 					(reg_q2577 AND symb_decoder(16#09#)) OR
 					(reg_q2577 AND symb_decoder(16#20#)) OR
 					(reg_q2577 AND symb_decoder(16#0d#)) OR
 					(reg_q2577 AND symb_decoder(16#0c#));
reg_q955_in <= (reg_q955 AND symb_decoder(16#1d#)) OR
 					(reg_q955 AND symb_decoder(16#48#)) OR
 					(reg_q955 AND symb_decoder(16#5f#)) OR
 					(reg_q955 AND symb_decoder(16#d5#)) OR
 					(reg_q955 AND symb_decoder(16#86#)) OR
 					(reg_q955 AND symb_decoder(16#6b#)) OR
 					(reg_q955 AND symb_decoder(16#9e#)) OR
 					(reg_q955 AND symb_decoder(16#c7#)) OR
 					(reg_q955 AND symb_decoder(16#97#)) OR
 					(reg_q955 AND symb_decoder(16#8c#)) OR
 					(reg_q955 AND symb_decoder(16#ef#)) OR
 					(reg_q955 AND symb_decoder(16#c5#)) OR
 					(reg_q955 AND symb_decoder(16#28#)) OR
 					(reg_q955 AND symb_decoder(16#ed#)) OR
 					(reg_q955 AND symb_decoder(16#0b#)) OR
 					(reg_q955 AND symb_decoder(16#aa#)) OR
 					(reg_q955 AND symb_decoder(16#70#)) OR
 					(reg_q955 AND symb_decoder(16#fc#)) OR
 					(reg_q955 AND symb_decoder(16#19#)) OR
 					(reg_q955 AND symb_decoder(16#88#)) OR
 					(reg_q955 AND symb_decoder(16#69#)) OR
 					(reg_q955 AND symb_decoder(16#12#)) OR
 					(reg_q955 AND symb_decoder(16#04#)) OR
 					(reg_q955 AND symb_decoder(16#e2#)) OR
 					(reg_q955 AND symb_decoder(16#4a#)) OR
 					(reg_q955 AND symb_decoder(16#74#)) OR
 					(reg_q955 AND symb_decoder(16#fb#)) OR
 					(reg_q955 AND symb_decoder(16#1e#)) OR
 					(reg_q955 AND symb_decoder(16#07#)) OR
 					(reg_q955 AND symb_decoder(16#2c#)) OR
 					(reg_q955 AND symb_decoder(16#0f#)) OR
 					(reg_q955 AND symb_decoder(16#da#)) OR
 					(reg_q955 AND symb_decoder(16#cf#)) OR
 					(reg_q955 AND symb_decoder(16#fe#)) OR
 					(reg_q955 AND symb_decoder(16#9c#)) OR
 					(reg_q955 AND symb_decoder(16#be#)) OR
 					(reg_q955 AND symb_decoder(16#4c#)) OR
 					(reg_q955 AND symb_decoder(16#d8#)) OR
 					(reg_q955 AND symb_decoder(16#87#)) OR
 					(reg_q955 AND symb_decoder(16#83#)) OR
 					(reg_q955 AND symb_decoder(16#f4#)) OR
 					(reg_q955 AND symb_decoder(16#52#)) OR
 					(reg_q955 AND symb_decoder(16#9d#)) OR
 					(reg_q955 AND symb_decoder(16#22#)) OR
 					(reg_q955 AND symb_decoder(16#29#)) OR
 					(reg_q955 AND symb_decoder(16#60#)) OR
 					(reg_q955 AND symb_decoder(16#31#)) OR
 					(reg_q955 AND symb_decoder(16#b8#)) OR
 					(reg_q955 AND symb_decoder(16#0c#)) OR
 					(reg_q955 AND symb_decoder(16#4f#)) OR
 					(reg_q955 AND symb_decoder(16#16#)) OR
 					(reg_q955 AND symb_decoder(16#9f#)) OR
 					(reg_q955 AND symb_decoder(16#c0#)) OR
 					(reg_q955 AND symb_decoder(16#ce#)) OR
 					(reg_q955 AND symb_decoder(16#d2#)) OR
 					(reg_q955 AND symb_decoder(16#e8#)) OR
 					(reg_q955 AND symb_decoder(16#3c#)) OR
 					(reg_q955 AND symb_decoder(16#27#)) OR
 					(reg_q955 AND symb_decoder(16#a7#)) OR
 					(reg_q955 AND symb_decoder(16#57#)) OR
 					(reg_q955 AND symb_decoder(16#d4#)) OR
 					(reg_q955 AND symb_decoder(16#c9#)) OR
 					(reg_q955 AND symb_decoder(16#6a#)) OR
 					(reg_q955 AND symb_decoder(16#f6#)) OR
 					(reg_q955 AND symb_decoder(16#41#)) OR
 					(reg_q955 AND symb_decoder(16#51#)) OR
 					(reg_q955 AND symb_decoder(16#06#)) OR
 					(reg_q955 AND symb_decoder(16#89#)) OR
 					(reg_q955 AND symb_decoder(16#b1#)) OR
 					(reg_q955 AND symb_decoder(16#17#)) OR
 					(reg_q955 AND symb_decoder(16#26#)) OR
 					(reg_q955 AND symb_decoder(16#e4#)) OR
 					(reg_q955 AND symb_decoder(16#3f#)) OR
 					(reg_q955 AND symb_decoder(16#44#)) OR
 					(reg_q955 AND symb_decoder(16#dd#)) OR
 					(reg_q955 AND symb_decoder(16#77#)) OR
 					(reg_q955 AND symb_decoder(16#62#)) OR
 					(reg_q955 AND symb_decoder(16#7c#)) OR
 					(reg_q955 AND symb_decoder(16#00#)) OR
 					(reg_q955 AND symb_decoder(16#b2#)) OR
 					(reg_q955 AND symb_decoder(16#73#)) OR
 					(reg_q955 AND symb_decoder(16#14#)) OR
 					(reg_q955 AND symb_decoder(16#72#)) OR
 					(reg_q955 AND symb_decoder(16#8d#)) OR
 					(reg_q955 AND symb_decoder(16#ca#)) OR
 					(reg_q955 AND symb_decoder(16#f2#)) OR
 					(reg_q955 AND symb_decoder(16#f9#)) OR
 					(reg_q955 AND symb_decoder(16#03#)) OR
 					(reg_q955 AND symb_decoder(16#3a#)) OR
 					(reg_q955 AND symb_decoder(16#2a#)) OR
 					(reg_q955 AND symb_decoder(16#01#)) OR
 					(reg_q955 AND symb_decoder(16#38#)) OR
 					(reg_q955 AND symb_decoder(16#c8#)) OR
 					(reg_q955 AND symb_decoder(16#96#)) OR
 					(reg_q955 AND symb_decoder(16#24#)) OR
 					(reg_q955 AND symb_decoder(16#c2#)) OR
 					(reg_q955 AND symb_decoder(16#d3#)) OR
 					(reg_q955 AND symb_decoder(16#e6#)) OR
 					(reg_q955 AND symb_decoder(16#09#)) OR
 					(reg_q955 AND symb_decoder(16#32#)) OR
 					(reg_q955 AND symb_decoder(16#58#)) OR
 					(reg_q955 AND symb_decoder(16#e9#)) OR
 					(reg_q955 AND symb_decoder(16#dc#)) OR
 					(reg_q955 AND symb_decoder(16#f8#)) OR
 					(reg_q955 AND symb_decoder(16#d9#)) OR
 					(reg_q955 AND symb_decoder(16#ab#)) OR
 					(reg_q955 AND symb_decoder(16#34#)) OR
 					(reg_q955 AND symb_decoder(16#47#)) OR
 					(reg_q955 AND symb_decoder(16#3d#)) OR
 					(reg_q955 AND symb_decoder(16#f7#)) OR
 					(reg_q955 AND symb_decoder(16#d6#)) OR
 					(reg_q955 AND symb_decoder(16#a5#)) OR
 					(reg_q955 AND symb_decoder(16#35#)) OR
 					(reg_q955 AND symb_decoder(16#d1#)) OR
 					(reg_q955 AND symb_decoder(16#98#)) OR
 					(reg_q955 AND symb_decoder(16#ad#)) OR
 					(reg_q955 AND symb_decoder(16#53#)) OR
 					(reg_q955 AND symb_decoder(16#92#)) OR
 					(reg_q955 AND symb_decoder(16#c1#)) OR
 					(reg_q955 AND symb_decoder(16#ff#)) OR
 					(reg_q955 AND symb_decoder(16#85#)) OR
 					(reg_q955 AND symb_decoder(16#bc#)) OR
 					(reg_q955 AND symb_decoder(16#b4#)) OR
 					(reg_q955 AND symb_decoder(16#c3#)) OR
 					(reg_q955 AND symb_decoder(16#a3#)) OR
 					(reg_q955 AND symb_decoder(16#56#)) OR
 					(reg_q955 AND symb_decoder(16#75#)) OR
 					(reg_q955 AND symb_decoder(16#c6#)) OR
 					(reg_q955 AND symb_decoder(16#02#)) OR
 					(reg_q955 AND symb_decoder(16#b9#)) OR
 					(reg_q955 AND symb_decoder(16#64#)) OR
 					(reg_q955 AND symb_decoder(16#6c#)) OR
 					(reg_q955 AND symb_decoder(16#1a#)) OR
 					(reg_q955 AND symb_decoder(16#e0#)) OR
 					(reg_q955 AND symb_decoder(16#f3#)) OR
 					(reg_q955 AND symb_decoder(16#45#)) OR
 					(reg_q955 AND symb_decoder(16#eb#)) OR
 					(reg_q955 AND symb_decoder(16#3e#)) OR
 					(reg_q955 AND symb_decoder(16#f1#)) OR
 					(reg_q955 AND symb_decoder(16#20#)) OR
 					(reg_q955 AND symb_decoder(16#91#)) OR
 					(reg_q955 AND symb_decoder(16#9a#)) OR
 					(reg_q955 AND symb_decoder(16#cc#)) OR
 					(reg_q955 AND symb_decoder(16#d7#)) OR
 					(reg_q955 AND symb_decoder(16#5a#)) OR
 					(reg_q955 AND symb_decoder(16#b6#)) OR
 					(reg_q955 AND symb_decoder(16#df#)) OR
 					(reg_q955 AND symb_decoder(16#43#)) OR
 					(reg_q955 AND symb_decoder(16#8b#)) OR
 					(reg_q955 AND symb_decoder(16#d0#)) OR
 					(reg_q955 AND symb_decoder(16#2d#)) OR
 					(reg_q955 AND symb_decoder(16#ee#)) OR
 					(reg_q955 AND symb_decoder(16#e1#)) OR
 					(reg_q955 AND symb_decoder(16#ec#)) OR
 					(reg_q955 AND symb_decoder(16#1f#)) OR
 					(reg_q955 AND symb_decoder(16#4b#)) OR
 					(reg_q955 AND symb_decoder(16#61#)) OR
 					(reg_q955 AND symb_decoder(16#55#)) OR
 					(reg_q955 AND symb_decoder(16#e7#)) OR
 					(reg_q955 AND symb_decoder(16#76#)) OR
 					(reg_q955 AND symb_decoder(16#82#)) OR
 					(reg_q955 AND symb_decoder(16#ae#)) OR
 					(reg_q955 AND symb_decoder(16#e3#)) OR
 					(reg_q955 AND symb_decoder(16#4d#)) OR
 					(reg_q955 AND symb_decoder(16#79#)) OR
 					(reg_q955 AND symb_decoder(16#49#)) OR
 					(reg_q955 AND symb_decoder(16#af#)) OR
 					(reg_q955 AND symb_decoder(16#63#)) OR
 					(reg_q955 AND symb_decoder(16#13#)) OR
 					(reg_q955 AND symb_decoder(16#b3#)) OR
 					(reg_q955 AND symb_decoder(16#33#)) OR
 					(reg_q955 AND symb_decoder(16#81#)) OR
 					(reg_q955 AND symb_decoder(16#a1#)) OR
 					(reg_q955 AND symb_decoder(16#59#)) OR
 					(reg_q955 AND symb_decoder(16#71#)) OR
 					(reg_q955 AND symb_decoder(16#6d#)) OR
 					(reg_q955 AND symb_decoder(16#7b#)) OR
 					(reg_q955 AND symb_decoder(16#65#)) OR
 					(reg_q955 AND symb_decoder(16#18#)) OR
 					(reg_q955 AND symb_decoder(16#37#)) OR
 					(reg_q955 AND symb_decoder(16#a8#)) OR
 					(reg_q955 AND symb_decoder(16#fa#)) OR
 					(reg_q955 AND symb_decoder(16#90#)) OR
 					(reg_q955 AND symb_decoder(16#9b#)) OR
 					(reg_q955 AND symb_decoder(16#bd#)) OR
 					(reg_q955 AND symb_decoder(16#a2#)) OR
 					(reg_q955 AND symb_decoder(16#f5#)) OR
 					(reg_q955 AND symb_decoder(16#78#)) OR
 					(reg_q955 AND symb_decoder(16#cb#)) OR
 					(reg_q955 AND symb_decoder(16#0e#)) OR
 					(reg_q955 AND symb_decoder(16#94#)) OR
 					(reg_q955 AND symb_decoder(16#15#)) OR
 					(reg_q955 AND symb_decoder(16#1b#)) OR
 					(reg_q955 AND symb_decoder(16#93#)) OR
 					(reg_q955 AND symb_decoder(16#f0#)) OR
 					(reg_q955 AND symb_decoder(16#84#)) OR
 					(reg_q955 AND symb_decoder(16#7d#)) OR
 					(reg_q955 AND symb_decoder(16#67#)) OR
 					(reg_q955 AND symb_decoder(16#2b#)) OR
 					(reg_q955 AND symb_decoder(16#bf#)) OR
 					(reg_q955 AND symb_decoder(16#8e#)) OR
 					(reg_q955 AND symb_decoder(16#68#)) OR
 					(reg_q955 AND symb_decoder(16#b7#)) OR
 					(reg_q955 AND symb_decoder(16#6f#)) OR
 					(reg_q955 AND symb_decoder(16#36#)) OR
 					(reg_q955 AND symb_decoder(16#23#)) OR
 					(reg_q955 AND symb_decoder(16#2f#)) OR
 					(reg_q955 AND symb_decoder(16#c4#)) OR
 					(reg_q955 AND symb_decoder(16#7f#)) OR
 					(reg_q955 AND symb_decoder(16#8a#)) OR
 					(reg_q955 AND symb_decoder(16#21#)) OR
 					(reg_q955 AND symb_decoder(16#95#)) OR
 					(reg_q955 AND symb_decoder(16#42#)) OR
 					(reg_q955 AND symb_decoder(16#25#)) OR
 					(reg_q955 AND symb_decoder(16#7e#)) OR
 					(reg_q955 AND symb_decoder(16#3b#)) OR
 					(reg_q955 AND symb_decoder(16#ac#)) OR
 					(reg_q955 AND symb_decoder(16#4e#)) OR
 					(reg_q955 AND symb_decoder(16#40#)) OR
 					(reg_q955 AND symb_decoder(16#cd#)) OR
 					(reg_q955 AND symb_decoder(16#54#)) OR
 					(reg_q955 AND symb_decoder(16#fd#)) OR
 					(reg_q955 AND symb_decoder(16#2e#)) OR
 					(reg_q955 AND symb_decoder(16#a4#)) OR
 					(reg_q955 AND symb_decoder(16#05#)) OR
 					(reg_q955 AND symb_decoder(16#ba#)) OR
 					(reg_q955 AND symb_decoder(16#80#)) OR
 					(reg_q955 AND symb_decoder(16#5e#)) OR
 					(reg_q955 AND symb_decoder(16#46#)) OR
 					(reg_q955 AND symb_decoder(16#e5#)) OR
 					(reg_q955 AND symb_decoder(16#a0#)) OR
 					(reg_q955 AND symb_decoder(16#5d#)) OR
 					(reg_q955 AND symb_decoder(16#a9#)) OR
 					(reg_q955 AND symb_decoder(16#de#)) OR
 					(reg_q955 AND symb_decoder(16#7a#)) OR
 					(reg_q955 AND symb_decoder(16#1c#)) OR
 					(reg_q955 AND symb_decoder(16#b5#)) OR
 					(reg_q955 AND symb_decoder(16#5c#)) OR
 					(reg_q955 AND symb_decoder(16#db#)) OR
 					(reg_q955 AND symb_decoder(16#8f#)) OR
 					(reg_q955 AND symb_decoder(16#11#)) OR
 					(reg_q955 AND symb_decoder(16#ea#)) OR
 					(reg_q955 AND symb_decoder(16#10#)) OR
 					(reg_q955 AND symb_decoder(16#6e#)) OR
 					(reg_q955 AND symb_decoder(16#5b#)) OR
 					(reg_q955 AND symb_decoder(16#66#)) OR
 					(reg_q955 AND symb_decoder(16#b0#)) OR
 					(reg_q955 AND symb_decoder(16#bb#)) OR
 					(reg_q955 AND symb_decoder(16#99#)) OR
 					(reg_q955 AND symb_decoder(16#30#)) OR
 					(reg_q955 AND symb_decoder(16#39#)) OR
 					(reg_q955 AND symb_decoder(16#08#)) OR
 					(reg_q955 AND symb_decoder(16#a6#)) OR
 					(reg_q955 AND symb_decoder(16#50#)) OR
 					(reg_q933 AND symb_decoder(16#45#)) OR
 					(reg_q933 AND symb_decoder(16#03#)) OR
 					(reg_q933 AND symb_decoder(16#eb#)) OR
 					(reg_q933 AND symb_decoder(16#3e#)) OR
 					(reg_q933 AND symb_decoder(16#2a#)) OR
 					(reg_q933 AND symb_decoder(16#01#)) OR
 					(reg_q933 AND symb_decoder(16#6d#)) OR
 					(reg_q933 AND symb_decoder(16#cc#)) OR
 					(reg_q933 AND symb_decoder(16#d7#)) OR
 					(reg_q933 AND symb_decoder(16#7b#)) OR
 					(reg_q933 AND symb_decoder(16#ad#)) OR
 					(reg_q933 AND symb_decoder(16#53#)) OR
 					(reg_q933 AND symb_decoder(16#92#)) OR
 					(reg_q933 AND symb_decoder(16#09#)) OR
 					(reg_q933 AND symb_decoder(16#fa#)) OR
 					(reg_q933 AND symb_decoder(16#9b#)) OR
 					(reg_q933 AND symb_decoder(16#58#)) OR
 					(reg_q933 AND symb_decoder(16#bc#)) OR
 					(reg_q933 AND symb_decoder(16#56#)) OR
 					(reg_q933 AND symb_decoder(16#2d#)) OR
 					(reg_q933 AND symb_decoder(16#dc#)) OR
 					(reg_q933 AND symb_decoder(16#4b#)) OR
 					(reg_q933 AND symb_decoder(16#61#)) OR
 					(reg_q933 AND symb_decoder(16#e7#)) OR
 					(reg_q933 AND symb_decoder(16#76#)) OR
 					(reg_q933 AND symb_decoder(16#f7#)) OR
 					(reg_q933 AND symb_decoder(16#64#)) OR
 					(reg_q933 AND symb_decoder(16#84#)) OR
 					(reg_q933 AND symb_decoder(16#1a#)) OR
 					(reg_q933 AND symb_decoder(16#7d#)) OR
 					(reg_q933 AND symb_decoder(16#79#)) OR
 					(reg_q933 AND symb_decoder(16#af#)) OR
 					(reg_q933 AND symb_decoder(16#8e#)) OR
 					(reg_q933 AND symb_decoder(16#35#)) OR
 					(reg_q933 AND symb_decoder(16#25#)) OR
 					(reg_q933 AND symb_decoder(16#18#)) OR
 					(reg_q933 AND symb_decoder(16#37#)) OR
 					(reg_q933 AND symb_decoder(16#ff#)) OR
 					(reg_q933 AND symb_decoder(16#bd#)) OR
 					(reg_q933 AND symb_decoder(16#f5#)) OR
 					(reg_q933 AND symb_decoder(16#43#)) OR
 					(reg_q933 AND symb_decoder(16#d0#)) OR
 					(reg_q933 AND symb_decoder(16#c3#)) OR
 					(reg_q933 AND symb_decoder(16#a3#)) OR
 					(reg_q933 AND symb_decoder(16#e1#)) OR
 					(reg_q933 AND symb_decoder(16#ec#)) OR
 					(reg_q933 AND symb_decoder(16#94#)) OR
 					(reg_q933 AND symb_decoder(16#75#)) OR
 					(reg_q933 AND symb_decoder(16#40#)) OR
 					(reg_q933 AND symb_decoder(16#02#)) OR
 					(reg_q933 AND symb_decoder(16#55#)) OR
 					(reg_q933 AND symb_decoder(16#e3#)) OR
 					(reg_q933 AND symb_decoder(16#05#)) OR
 					(reg_q933 AND symb_decoder(16#ba#)) OR
 					(reg_q933 AND symb_decoder(16#49#)) OR
 					(reg_q933 AND symb_decoder(16#46#)) OR
 					(reg_q933 AND symb_decoder(16#2b#)) OR
 					(reg_q933 AND symb_decoder(16#68#)) OR
 					(reg_q933 AND symb_decoder(16#63#)) OR
 					(reg_q933 AND symb_decoder(16#f3#)) OR
 					(reg_q933 AND symb_decoder(16#13#)) OR
 					(reg_q933 AND symb_decoder(16#6f#)) OR
 					(reg_q933 AND symb_decoder(16#a1#)) OR
 					(reg_q933 AND symb_decoder(16#23#)) OR
 					(reg_q933 AND symb_decoder(16#00#)) OR
 					(reg_q933 AND symb_decoder(16#5c#)) OR
 					(reg_q933 AND symb_decoder(16#c4#)) OR
 					(reg_q933 AND symb_decoder(16#71#)) OR
 					(reg_q933 AND symb_decoder(16#20#)) OR
 					(reg_q933 AND symb_decoder(16#11#)) OR
 					(reg_q933 AND symb_decoder(16#42#)) OR
 					(reg_q933 AND symb_decoder(16#df#)) OR
 					(reg_q933 AND symb_decoder(16#6e#)) OR
 					(reg_q933 AND symb_decoder(16#5b#)) OR
 					(reg_q933 AND symb_decoder(16#65#)) OR
 					(reg_q933 AND symb_decoder(16#90#)) OR
 					(reg_q933 AND symb_decoder(16#a2#)) OR
 					(reg_q933 AND symb_decoder(16#08#)) OR
 					(reg_q933 AND symb_decoder(16#8b#)) OR
 					(reg_q933 AND symb_decoder(16#ee#)) OR
 					(reg_q933 AND symb_decoder(16#0e#)) OR
 					(reg_q933 AND symb_decoder(16#1d#)) OR
 					(reg_q933 AND symb_decoder(16#15#)) OR
 					(reg_q933 AND symb_decoder(16#4e#)) OR
 					(reg_q933 AND symb_decoder(16#48#)) OR
 					(reg_q933 AND symb_decoder(16#d5#)) OR
 					(reg_q933 AND symb_decoder(16#93#)) OR
 					(reg_q933 AND symb_decoder(16#82#)) OR
 					(reg_q933 AND symb_decoder(16#2e#)) OR
 					(reg_q933 AND symb_decoder(16#f0#)) OR
 					(reg_q933 AND symb_decoder(16#8c#)) OR
 					(reg_q933 AND symb_decoder(16#ef#)) OR
 					(reg_q933 AND symb_decoder(16#ae#)) OR
 					(reg_q933 AND symb_decoder(16#67#)) OR
 					(reg_q933 AND symb_decoder(16#b7#)) OR
 					(reg_q933 AND symb_decoder(16#b3#)) OR
 					(reg_q933 AND symb_decoder(16#81#)) OR
 					(reg_q933 AND symb_decoder(16#36#)) OR
 					(reg_q933 AND symb_decoder(16#de#)) OR
 					(reg_q933 AND symb_decoder(16#2f#)) OR
 					(reg_q933 AND symb_decoder(16#59#)) OR
 					(reg_q933 AND symb_decoder(16#b5#)) OR
 					(reg_q933 AND symb_decoder(16#ea#)) OR
 					(reg_q933 AND symb_decoder(16#10#)) OR
 					(reg_q933 AND symb_decoder(16#a8#)) OR
 					(reg_q933 AND symb_decoder(16#bb#)) OR
 					(reg_q933 AND symb_decoder(16#fb#)) OR
 					(reg_q933 AND symb_decoder(16#1e#)) OR
 					(reg_q933 AND symb_decoder(16#a6#)) OR
 					(reg_q933 AND symb_decoder(16#78#)) OR
 					(reg_q933 AND symb_decoder(16#cb#)) OR
 					(reg_q933 AND symb_decoder(16#da#)) OR
 					(reg_q933 AND symb_decoder(16#cf#)) OR
 					(reg_q933 AND symb_decoder(16#3b#)) OR
 					(reg_q933 AND symb_decoder(16#1b#)) OR
 					(reg_q933 AND symb_decoder(16#5f#)) OR
 					(reg_q933 AND symb_decoder(16#4c#)) OR
 					(reg_q933 AND symb_decoder(16#87#)) OR
 					(reg_q933 AND symb_decoder(16#f4#)) OR
 					(reg_q933 AND symb_decoder(16#cd#)) OR
 					(reg_q933 AND symb_decoder(16#54#)) OR
 					(reg_q933 AND symb_decoder(16#9d#)) OR
 					(reg_q933 AND symb_decoder(16#29#)) OR
 					(reg_q933 AND symb_decoder(16#a4#)) OR
 					(reg_q933 AND symb_decoder(16#5e#)) OR
 					(reg_q933 AND symb_decoder(16#ed#)) OR
 					(reg_q933 AND symb_decoder(16#e5#)) OR
 					(reg_q933 AND symb_decoder(16#bf#)) OR
 					(reg_q933 AND symb_decoder(16#ce#)) OR
 					(reg_q933 AND symb_decoder(16#7a#)) OR
 					(reg_q933 AND symb_decoder(16#d2#)) OR
 					(reg_q933 AND symb_decoder(16#8f#)) OR
 					(reg_q933 AND symb_decoder(16#7f#)) OR
 					(reg_q933 AND symb_decoder(16#27#)) OR
 					(reg_q933 AND symb_decoder(16#a7#)) OR
 					(reg_q933 AND symb_decoder(16#88#)) OR
 					(reg_q933 AND symb_decoder(16#8a#)) OR
 					(reg_q933 AND symb_decoder(16#21#)) OR
 					(reg_q933 AND symb_decoder(16#95#)) OR
 					(reg_q933 AND symb_decoder(16#12#)) OR
 					(reg_q933 AND symb_decoder(16#04#)) OR
 					(reg_q933 AND symb_decoder(16#66#)) OR
 					(reg_q933 AND symb_decoder(16#6a#)) OR
 					(reg_q933 AND symb_decoder(16#b0#)) OR
 					(reg_q933 AND symb_decoder(16#30#)) OR
 					(reg_q933 AND symb_decoder(16#39#)) OR
 					(reg_q933 AND symb_decoder(16#89#)) OR
 					(reg_q933 AND symb_decoder(16#7e#)) OR
 					(reg_q933 AND symb_decoder(16#ac#)) OR
 					(reg_q933 AND symb_decoder(16#e4#)) OR
 					(reg_q933 AND symb_decoder(16#6b#)) OR
 					(reg_q933 AND symb_decoder(16#fd#)) OR
 					(reg_q933 AND symb_decoder(16#22#)) OR
 					(reg_q933 AND symb_decoder(16#97#)) OR
 					(reg_q933 AND symb_decoder(16#80#)) OR
 					(reg_q933 AND symb_decoder(16#44#)) OR
 					(reg_q933 AND symb_decoder(16#c5#)) OR
 					(reg_q933 AND symb_decoder(16#dd#)) OR
 					(reg_q933 AND symb_decoder(16#77#)) OR
 					(reg_q933 AND symb_decoder(16#28#)) OR
 					(reg_q933 AND symb_decoder(16#a0#)) OR
 					(reg_q933 AND symb_decoder(16#5d#)) OR
 					(reg_q933 AND symb_decoder(16#0b#)) OR
 					(reg_q933 AND symb_decoder(16#a9#)) OR
 					(reg_q933 AND symb_decoder(16#b2#)) OR
 					(reg_q933 AND symb_decoder(16#9f#)) OR
 					(reg_q933 AND symb_decoder(16#73#)) OR
 					(reg_q933 AND symb_decoder(16#ca#)) OR
 					(reg_q933 AND symb_decoder(16#1c#)) OR
 					(reg_q933 AND symb_decoder(16#db#)) OR
 					(reg_q933 AND symb_decoder(16#fc#)) OR
 					(reg_q933 AND symb_decoder(16#38#)) OR
 					(reg_q933 AND symb_decoder(16#69#)) OR
 					(reg_q933 AND symb_decoder(16#96#)) OR
 					(reg_q933 AND symb_decoder(16#e2#)) OR
 					(reg_q933 AND symb_decoder(16#c9#)) OR
 					(reg_q933 AND symb_decoder(16#f6#)) OR
 					(reg_q933 AND symb_decoder(16#99#)) OR
 					(reg_q933 AND symb_decoder(16#51#)) OR
 					(reg_q933 AND symb_decoder(16#0f#)) OR
 					(reg_q933 AND symb_decoder(16#50#)) OR
 					(reg_q933 AND symb_decoder(16#fe#)) OR
 					(reg_q933 AND symb_decoder(16#f8#)) OR
 					(reg_q933 AND symb_decoder(16#d9#)) OR
 					(reg_q933 AND symb_decoder(16#ab#)) OR
 					(reg_q933 AND symb_decoder(16#be#)) OR
 					(reg_q933 AND symb_decoder(16#34#)) OR
 					(reg_q933 AND symb_decoder(16#86#)) OR
 					(reg_q933 AND symb_decoder(16#d8#)) OR
 					(reg_q933 AND symb_decoder(16#52#)) OR
 					(reg_q933 AND symb_decoder(16#9e#)) OR
 					(reg_q933 AND symb_decoder(16#c7#)) OR
 					(reg_q933 AND symb_decoder(16#3f#)) OR
 					(reg_q933 AND symb_decoder(16#b8#)) OR
 					(reg_q933 AND symb_decoder(16#aa#)) OR
 					(reg_q933 AND symb_decoder(16#0c#)) OR
 					(reg_q933 AND symb_decoder(16#4f#)) OR
 					(reg_q933 AND symb_decoder(16#16#)) OR
 					(reg_q933 AND symb_decoder(16#d1#)) OR
 					(reg_q933 AND symb_decoder(16#c0#)) OR
 					(reg_q933 AND symb_decoder(16#98#)) OR
 					(reg_q933 AND symb_decoder(16#f2#)) OR
 					(reg_q933 AND symb_decoder(16#f9#)) OR
 					(reg_q933 AND symb_decoder(16#3a#)) OR
 					(reg_q933 AND symb_decoder(16#70#)) OR
 					(reg_q933 AND symb_decoder(16#3c#)) OR
 					(reg_q933 AND symb_decoder(16#19#)) OR
 					(reg_q933 AND symb_decoder(16#57#)) OR
 					(reg_q933 AND symb_decoder(16#d4#)) OR
 					(reg_q933 AND symb_decoder(16#e6#)) OR
 					(reg_q933 AND symb_decoder(16#4a#)) OR
 					(reg_q933 AND symb_decoder(16#c1#)) OR
 					(reg_q933 AND symb_decoder(16#74#)) OR
 					(reg_q933 AND symb_decoder(16#85#)) OR
 					(reg_q933 AND symb_decoder(16#06#)) OR
 					(reg_q933 AND symb_decoder(16#07#)) OR
 					(reg_q933 AND symb_decoder(16#2c#)) OR
 					(reg_q933 AND symb_decoder(16#b1#)) OR
 					(reg_q933 AND symb_decoder(16#26#)) OR
 					(reg_q933 AND symb_decoder(16#c6#)) OR
 					(reg_q933 AND symb_decoder(16#9c#)) OR
 					(reg_q933 AND symb_decoder(16#47#)) OR
 					(reg_q933 AND symb_decoder(16#83#)) OR
 					(reg_q933 AND symb_decoder(16#b9#)) OR
 					(reg_q933 AND symb_decoder(16#3d#)) OR
 					(reg_q933 AND symb_decoder(16#6c#)) OR
 					(reg_q933 AND symb_decoder(16#60#)) OR
 					(reg_q933 AND symb_decoder(16#d6#)) OR
 					(reg_q933 AND symb_decoder(16#31#)) OR
 					(reg_q933 AND symb_decoder(16#e0#)) OR
 					(reg_q933 AND symb_decoder(16#7c#)) OR
 					(reg_q933 AND symb_decoder(16#14#)) OR
 					(reg_q933 AND symb_decoder(16#72#)) OR
 					(reg_q933 AND symb_decoder(16#8d#)) OR
 					(reg_q933 AND symb_decoder(16#e8#)) OR
 					(reg_q933 AND symb_decoder(16#f1#)) OR
 					(reg_q933 AND symb_decoder(16#91#)) OR
 					(reg_q933 AND symb_decoder(16#9a#)) OR
 					(reg_q933 AND symb_decoder(16#5a#)) OR
 					(reg_q933 AND symb_decoder(16#c8#)) OR
 					(reg_q933 AND symb_decoder(16#b6#)) OR
 					(reg_q933 AND symb_decoder(16#24#)) OR
 					(reg_q933 AND symb_decoder(16#c2#)) OR
 					(reg_q933 AND symb_decoder(16#d3#)) OR
 					(reg_q933 AND symb_decoder(16#32#)) OR
 					(reg_q933 AND symb_decoder(16#41#)) OR
 					(reg_q933 AND symb_decoder(16#b4#)) OR
 					(reg_q933 AND symb_decoder(16#e9#)) OR
 					(reg_q933 AND symb_decoder(16#17#)) OR
 					(reg_q933 AND symb_decoder(16#1f#)) OR
 					(reg_q933 AND symb_decoder(16#4d#)) OR
 					(reg_q933 AND symb_decoder(16#a5#)) OR
 					(reg_q933 AND symb_decoder(16#62#)) OR
 					(reg_q933 AND symb_decoder(16#33#));
reg_q933_in <= (reg_q931 AND symb_decoder(16#00#));
reg_q251_in <= (reg_q249 AND symb_decoder(16#ff#));
reg_q253_in <= (reg_q251 AND symb_decoder(16#36#)) OR
 					(reg_q251 AND symb_decoder(16#39#)) OR
 					(reg_q251 AND symb_decoder(16#34#)) OR
 					(reg_q251 AND symb_decoder(16#33#)) OR
 					(reg_q251 AND symb_decoder(16#37#)) OR
 					(reg_q251 AND symb_decoder(16#30#)) OR
 					(reg_q251 AND symb_decoder(16#35#)) OR
 					(reg_q251 AND symb_decoder(16#38#)) OR
 					(reg_q251 AND symb_decoder(16#31#)) OR
 					(reg_q251 AND symb_decoder(16#32#)) OR
 					(reg_q253 AND symb_decoder(16#35#)) OR
 					(reg_q253 AND symb_decoder(16#31#)) OR
 					(reg_q253 AND symb_decoder(16#30#)) OR
 					(reg_q253 AND symb_decoder(16#33#)) OR
 					(reg_q253 AND symb_decoder(16#32#)) OR
 					(reg_q253 AND symb_decoder(16#38#)) OR
 					(reg_q253 AND symb_decoder(16#39#)) OR
 					(reg_q253 AND symb_decoder(16#37#)) OR
 					(reg_q253 AND symb_decoder(16#36#)) OR
 					(reg_q253 AND symb_decoder(16#34#));
reg_q1331_in <= (reg_q1329 AND symb_decoder(16#72#)) OR
 					(reg_q1329 AND symb_decoder(16#52#));
reg_q1333_in <= (reg_q1331 AND symb_decoder(16#09#)) OR
 					(reg_q1331 AND symb_decoder(16#0a#)) OR
 					(reg_q1331 AND symb_decoder(16#20#)) OR
 					(reg_q1331 AND symb_decoder(16#0c#)) OR
 					(reg_q1331 AND symb_decoder(16#0d#)) OR
 					(reg_q1333 AND symb_decoder(16#20#)) OR
 					(reg_q1333 AND symb_decoder(16#0c#)) OR
 					(reg_q1333 AND symb_decoder(16#09#)) OR
 					(reg_q1333 AND symb_decoder(16#0a#)) OR
 					(reg_q1333 AND symb_decoder(16#0d#));
reg_q1997_in <= (reg_q1997 AND symb_decoder(16#a1#)) OR
 					(reg_q1997 AND symb_decoder(16#3d#)) OR
 					(reg_q1997 AND symb_decoder(16#9b#)) OR
 					(reg_q1997 AND symb_decoder(16#af#)) OR
 					(reg_q1997 AND symb_decoder(16#96#)) OR
 					(reg_q1997 AND symb_decoder(16#ab#)) OR
 					(reg_q1997 AND symb_decoder(16#f2#)) OR
 					(reg_q1997 AND symb_decoder(16#18#)) OR
 					(reg_q1997 AND symb_decoder(16#58#)) OR
 					(reg_q1997 AND symb_decoder(16#d0#)) OR
 					(reg_q1997 AND symb_decoder(16#d5#)) OR
 					(reg_q1997 AND symb_decoder(16#bb#)) OR
 					(reg_q1997 AND symb_decoder(16#16#)) OR
 					(reg_q1997 AND symb_decoder(16#ce#)) OR
 					(reg_q1997 AND symb_decoder(16#11#)) OR
 					(reg_q1997 AND symb_decoder(16#be#)) OR
 					(reg_q1997 AND symb_decoder(16#bd#)) OR
 					(reg_q1997 AND symb_decoder(16#8d#)) OR
 					(reg_q1997 AND symb_decoder(16#f3#)) OR
 					(reg_q1997 AND symb_decoder(16#89#)) OR
 					(reg_q1997 AND symb_decoder(16#88#)) OR
 					(reg_q1997 AND symb_decoder(16#e9#)) OR
 					(reg_q1997 AND symb_decoder(16#57#)) OR
 					(reg_q1997 AND symb_decoder(16#35#)) OR
 					(reg_q1997 AND symb_decoder(16#e2#)) OR
 					(reg_q1997 AND symb_decoder(16#2e#)) OR
 					(reg_q1997 AND symb_decoder(16#fd#)) OR
 					(reg_q1997 AND symb_decoder(16#7d#)) OR
 					(reg_q1997 AND symb_decoder(16#71#)) OR
 					(reg_q1997 AND symb_decoder(16#b9#)) OR
 					(reg_q1997 AND symb_decoder(16#08#)) OR
 					(reg_q1997 AND symb_decoder(16#d7#)) OR
 					(reg_q1997 AND symb_decoder(16#55#)) OR
 					(reg_q1997 AND symb_decoder(16#b3#)) OR
 					(reg_q1997 AND symb_decoder(16#3e#)) OR
 					(reg_q1997 AND symb_decoder(16#ad#)) OR
 					(reg_q1997 AND symb_decoder(16#2f#)) OR
 					(reg_q1997 AND symb_decoder(16#63#)) OR
 					(reg_q1997 AND symb_decoder(16#1b#)) OR
 					(reg_q1997 AND symb_decoder(16#cd#)) OR
 					(reg_q1997 AND symb_decoder(16#54#)) OR
 					(reg_q1997 AND symb_decoder(16#29#)) OR
 					(reg_q1997 AND symb_decoder(16#4d#)) OR
 					(reg_q1997 AND symb_decoder(16#d3#)) OR
 					(reg_q1997 AND symb_decoder(16#e8#)) OR
 					(reg_q1997 AND symb_decoder(16#a4#)) OR
 					(reg_q1997 AND symb_decoder(16#c5#)) OR
 					(reg_q1997 AND symb_decoder(16#59#)) OR
 					(reg_q1997 AND symb_decoder(16#c4#)) OR
 					(reg_q1997 AND symb_decoder(16#91#)) OR
 					(reg_q1997 AND symb_decoder(16#fc#)) OR
 					(reg_q1997 AND symb_decoder(16#dc#)) OR
 					(reg_q1997 AND symb_decoder(16#81#)) OR
 					(reg_q1997 AND symb_decoder(16#bc#)) OR
 					(reg_q1997 AND symb_decoder(16#f9#)) OR
 					(reg_q1997 AND symb_decoder(16#27#)) OR
 					(reg_q1997 AND symb_decoder(16#98#)) OR
 					(reg_q1997 AND symb_decoder(16#26#)) OR
 					(reg_q1997 AND symb_decoder(16#e6#)) OR
 					(reg_q1997 AND symb_decoder(16#75#)) OR
 					(reg_q1997 AND symb_decoder(16#b6#)) OR
 					(reg_q1997 AND symb_decoder(16#b5#)) OR
 					(reg_q1997 AND symb_decoder(16#5d#)) OR
 					(reg_q1997 AND symb_decoder(16#49#)) OR
 					(reg_q1997 AND symb_decoder(16#76#)) OR
 					(reg_q1997 AND symb_decoder(16#12#)) OR
 					(reg_q1997 AND symb_decoder(16#19#)) OR
 					(reg_q1997 AND symb_decoder(16#ac#)) OR
 					(reg_q1997 AND symb_decoder(16#bf#)) OR
 					(reg_q1997 AND symb_decoder(16#f1#)) OR
 					(reg_q1997 AND symb_decoder(16#28#)) OR
 					(reg_q1997 AND symb_decoder(16#c6#)) OR
 					(reg_q1997 AND symb_decoder(16#e4#)) OR
 					(reg_q1997 AND symb_decoder(16#de#)) OR
 					(reg_q1997 AND symb_decoder(16#2c#)) OR
 					(reg_q1997 AND symb_decoder(16#73#)) OR
 					(reg_q1997 AND symb_decoder(16#d1#)) OR
 					(reg_q1997 AND symb_decoder(16#3c#)) OR
 					(reg_q1997 AND symb_decoder(16#5f#)) OR
 					(reg_q1997 AND symb_decoder(16#51#)) OR
 					(reg_q1997 AND symb_decoder(16#ca#)) OR
 					(reg_q1997 AND symb_decoder(16#52#)) OR
 					(reg_q1997 AND symb_decoder(16#07#)) OR
 					(reg_q1997 AND symb_decoder(16#45#)) OR
 					(reg_q1997 AND symb_decoder(16#6a#)) OR
 					(reg_q1997 AND symb_decoder(16#78#)) OR
 					(reg_q1997 AND symb_decoder(16#b7#)) OR
 					(reg_q1997 AND symb_decoder(16#50#)) OR
 					(reg_q1997 AND symb_decoder(16#79#)) OR
 					(reg_q1997 AND symb_decoder(16#6b#)) OR
 					(reg_q1997 AND symb_decoder(16#36#)) OR
 					(reg_q1997 AND symb_decoder(16#ed#)) OR
 					(reg_q1997 AND symb_decoder(16#7c#)) OR
 					(reg_q1997 AND symb_decoder(16#cb#)) OR
 					(reg_q1997 AND symb_decoder(16#3f#)) OR
 					(reg_q1997 AND symb_decoder(16#48#)) OR
 					(reg_q1997 AND symb_decoder(16#23#)) OR
 					(reg_q1997 AND symb_decoder(16#ff#)) OR
 					(reg_q1997 AND symb_decoder(16#85#)) OR
 					(reg_q1997 AND symb_decoder(16#6d#)) OR
 					(reg_q1997 AND symb_decoder(16#8c#)) OR
 					(reg_q1997 AND symb_decoder(16#32#)) OR
 					(reg_q1997 AND symb_decoder(16#f7#)) OR
 					(reg_q1997 AND symb_decoder(16#c1#)) OR
 					(reg_q1997 AND symb_decoder(16#84#)) OR
 					(reg_q1997 AND symb_decoder(16#f0#)) OR
 					(reg_q1997 AND symb_decoder(16#1e#)) OR
 					(reg_q1997 AND symb_decoder(16#31#)) OR
 					(reg_q1997 AND symb_decoder(16#38#)) OR
 					(reg_q1997 AND symb_decoder(16#04#)) OR
 					(reg_q1997 AND symb_decoder(16#1f#)) OR
 					(reg_q1997 AND symb_decoder(16#6f#)) OR
 					(reg_q1997 AND symb_decoder(16#21#)) OR
 					(reg_q1997 AND symb_decoder(16#b8#)) OR
 					(reg_q1997 AND symb_decoder(16#2b#)) OR
 					(reg_q1997 AND symb_decoder(16#4f#)) OR
 					(reg_q1997 AND symb_decoder(16#a8#)) OR
 					(reg_q1997 AND symb_decoder(16#83#)) OR
 					(reg_q1997 AND symb_decoder(16#72#)) OR
 					(reg_q1997 AND symb_decoder(16#62#)) OR
 					(reg_q1997 AND symb_decoder(16#14#)) OR
 					(reg_q1997 AND symb_decoder(16#d8#)) OR
 					(reg_q1997 AND symb_decoder(16#95#)) OR
 					(reg_q1997 AND symb_decoder(16#d2#)) OR
 					(reg_q1997 AND symb_decoder(16#3b#)) OR
 					(reg_q1997 AND symb_decoder(16#0b#)) OR
 					(reg_q1997 AND symb_decoder(16#9d#)) OR
 					(reg_q1997 AND symb_decoder(16#86#)) OR
 					(reg_q1997 AND symb_decoder(16#8b#)) OR
 					(reg_q1997 AND symb_decoder(16#13#)) OR
 					(reg_q1997 AND symb_decoder(16#0e#)) OR
 					(reg_q1997 AND symb_decoder(16#43#)) OR
 					(reg_q1997 AND symb_decoder(16#da#)) OR
 					(reg_q1997 AND symb_decoder(16#df#)) OR
 					(reg_q1997 AND symb_decoder(16#0c#)) OR
 					(reg_q1997 AND symb_decoder(16#2d#)) OR
 					(reg_q1997 AND symb_decoder(16#39#)) OR
 					(reg_q1997 AND symb_decoder(16#9e#)) OR
 					(reg_q1997 AND symb_decoder(16#ea#)) OR
 					(reg_q1997 AND symb_decoder(16#cc#)) OR
 					(reg_q1997 AND symb_decoder(16#22#)) OR
 					(reg_q1997 AND symb_decoder(16#47#)) OR
 					(reg_q1997 AND symb_decoder(16#c0#)) OR
 					(reg_q1997 AND symb_decoder(16#8a#)) OR
 					(reg_q1997 AND symb_decoder(16#4a#)) OR
 					(reg_q1997 AND symb_decoder(16#cf#)) OR
 					(reg_q1997 AND symb_decoder(16#8e#)) OR
 					(reg_q1997 AND symb_decoder(16#37#)) OR
 					(reg_q1997 AND symb_decoder(16#93#)) OR
 					(reg_q1997 AND symb_decoder(16#68#)) OR
 					(reg_q1997 AND symb_decoder(16#4b#)) OR
 					(reg_q1997 AND symb_decoder(16#c3#)) OR
 					(reg_q1997 AND symb_decoder(16#9f#)) OR
 					(reg_q1997 AND symb_decoder(16#65#)) OR
 					(reg_q1997 AND symb_decoder(16#f6#)) OR
 					(reg_q1997 AND symb_decoder(16#5e#)) OR
 					(reg_q1997 AND symb_decoder(16#8f#)) OR
 					(reg_q1997 AND symb_decoder(16#06#)) OR
 					(reg_q1997 AND symb_decoder(16#1c#)) OR
 					(reg_q1997 AND symb_decoder(16#e3#)) OR
 					(reg_q1997 AND symb_decoder(16#ba#)) OR
 					(reg_q1997 AND symb_decoder(16#41#)) OR
 					(reg_q1997 AND symb_decoder(16#67#)) OR
 					(reg_q1997 AND symb_decoder(16#4e#)) OR
 					(reg_q1997 AND symb_decoder(16#44#)) OR
 					(reg_q1997 AND symb_decoder(16#94#)) OR
 					(reg_q1997 AND symb_decoder(16#aa#)) OR
 					(reg_q1997 AND symb_decoder(16#90#)) OR
 					(reg_q1997 AND symb_decoder(16#c7#)) OR
 					(reg_q1997 AND symb_decoder(16#b4#)) OR
 					(reg_q1997 AND symb_decoder(16#99#)) OR
 					(reg_q1997 AND symb_decoder(16#66#)) OR
 					(reg_q1997 AND symb_decoder(16#20#)) OR
 					(reg_q1997 AND symb_decoder(16#5c#)) OR
 					(reg_q1997 AND symb_decoder(16#ec#)) OR
 					(reg_q1997 AND symb_decoder(16#9c#)) OR
 					(reg_q1997 AND symb_decoder(16#d6#)) OR
 					(reg_q1997 AND symb_decoder(16#2a#)) OR
 					(reg_q1997 AND symb_decoder(16#dd#)) OR
 					(reg_q1997 AND symb_decoder(16#f5#)) OR
 					(reg_q1997 AND symb_decoder(16#d9#)) OR
 					(reg_q1997 AND symb_decoder(16#7a#)) OR
 					(reg_q1997 AND symb_decoder(16#25#)) OR
 					(reg_q1997 AND symb_decoder(16#09#)) OR
 					(reg_q1997 AND symb_decoder(16#10#)) OR
 					(reg_q1997 AND symb_decoder(16#70#)) OR
 					(reg_q1997 AND symb_decoder(16#56#)) OR
 					(reg_q1997 AND symb_decoder(16#fe#)) OR
 					(reg_q1997 AND symb_decoder(16#97#)) OR
 					(reg_q1997 AND symb_decoder(16#46#)) OR
 					(reg_q1997 AND symb_decoder(16#a9#)) OR
 					(reg_q1997 AND symb_decoder(16#15#)) OR
 					(reg_q1997 AND symb_decoder(16#f4#)) OR
 					(reg_q1997 AND symb_decoder(16#5b#)) OR
 					(reg_q1997 AND symb_decoder(16#77#)) OR
 					(reg_q1997 AND symb_decoder(16#fa#)) OR
 					(reg_q1997 AND symb_decoder(16#b2#)) OR
 					(reg_q1997 AND symb_decoder(16#30#)) OR
 					(reg_q1997 AND symb_decoder(16#5a#)) OR
 					(reg_q1997 AND symb_decoder(16#33#)) OR
 					(reg_q1997 AND symb_decoder(16#d4#)) OR
 					(reg_q1997 AND symb_decoder(16#7e#)) OR
 					(reg_q1997 AND symb_decoder(16#01#)) OR
 					(reg_q1997 AND symb_decoder(16#82#)) OR
 					(reg_q1997 AND symb_decoder(16#42#)) OR
 					(reg_q1997 AND symb_decoder(16#02#)) OR
 					(reg_q1997 AND symb_decoder(16#a7#)) OR
 					(reg_q1997 AND symb_decoder(16#a0#)) OR
 					(reg_q1997 AND symb_decoder(16#34#)) OR
 					(reg_q1997 AND symb_decoder(16#ee#)) OR
 					(reg_q1997 AND symb_decoder(16#c2#)) OR
 					(reg_q1997 AND symb_decoder(16#17#)) OR
 					(reg_q1997 AND symb_decoder(16#6e#)) OR
 					(reg_q1997 AND symb_decoder(16#0f#)) OR
 					(reg_q1997 AND symb_decoder(16#db#)) OR
 					(reg_q1997 AND symb_decoder(16#a3#)) OR
 					(reg_q1997 AND symb_decoder(16#ae#)) OR
 					(reg_q1997 AND symb_decoder(16#64#)) OR
 					(reg_q1997 AND symb_decoder(16#e0#)) OR
 					(reg_q1997 AND symb_decoder(16#92#)) OR
 					(reg_q1997 AND symb_decoder(16#c8#)) OR
 					(reg_q1997 AND symb_decoder(16#a5#)) OR
 					(reg_q1997 AND symb_decoder(16#80#)) OR
 					(reg_q1997 AND symb_decoder(16#ef#)) OR
 					(reg_q1997 AND symb_decoder(16#eb#)) OR
 					(reg_q1997 AND symb_decoder(16#9a#)) OR
 					(reg_q1997 AND symb_decoder(16#3a#)) OR
 					(reg_q1997 AND symb_decoder(16#03#)) OR
 					(reg_q1997 AND symb_decoder(16#87#)) OR
 					(reg_q1997 AND symb_decoder(16#7b#)) OR
 					(reg_q1997 AND symb_decoder(16#4c#)) OR
 					(reg_q1997 AND symb_decoder(16#a6#)) OR
 					(reg_q1997 AND symb_decoder(16#69#)) OR
 					(reg_q1997 AND symb_decoder(16#c9#)) OR
 					(reg_q1997 AND symb_decoder(16#05#)) OR
 					(reg_q1997 AND symb_decoder(16#fb#)) OR
 					(reg_q1997 AND symb_decoder(16#6c#)) OR
 					(reg_q1997 AND symb_decoder(16#40#)) OR
 					(reg_q1997 AND symb_decoder(16#a2#)) OR
 					(reg_q1997 AND symb_decoder(16#b1#)) OR
 					(reg_q1997 AND symb_decoder(16#53#)) OR
 					(reg_q1997 AND symb_decoder(16#e5#)) OR
 					(reg_q1997 AND symb_decoder(16#e1#)) OR
 					(reg_q1997 AND symb_decoder(16#b0#)) OR
 					(reg_q1997 AND symb_decoder(16#74#)) OR
 					(reg_q1997 AND symb_decoder(16#e7#)) OR
 					(reg_q1997 AND symb_decoder(16#1a#)) OR
 					(reg_q1997 AND symb_decoder(16#f8#)) OR
 					(reg_q1997 AND symb_decoder(16#24#)) OR
 					(reg_q1997 AND symb_decoder(16#00#)) OR
 					(reg_q1997 AND symb_decoder(16#60#)) OR
 					(reg_q1997 AND symb_decoder(16#61#)) OR
 					(reg_q1997 AND symb_decoder(16#1d#)) OR
 					(reg_q1997 AND symb_decoder(16#7f#)) OR
 					(reg_q1975 AND symb_decoder(16#9e#)) OR
 					(reg_q1975 AND symb_decoder(16#4a#)) OR
 					(reg_q1975 AND symb_decoder(16#be#)) OR
 					(reg_q1975 AND symb_decoder(16#8a#)) OR
 					(reg_q1975 AND symb_decoder(16#5a#)) OR
 					(reg_q1975 AND symb_decoder(16#0e#)) OR
 					(reg_q1975 AND symb_decoder(16#43#)) OR
 					(reg_q1975 AND symb_decoder(16#d8#)) OR
 					(reg_q1975 AND symb_decoder(16#cf#)) OR
 					(reg_q1975 AND symb_decoder(16#6b#)) OR
 					(reg_q1975 AND symb_decoder(16#b3#)) OR
 					(reg_q1975 AND symb_decoder(16#3b#)) OR
 					(reg_q1975 AND symb_decoder(16#ff#)) OR
 					(reg_q1975 AND symb_decoder(16#35#)) OR
 					(reg_q1975 AND symb_decoder(16#ad#)) OR
 					(reg_q1975 AND symb_decoder(16#bf#)) OR
 					(reg_q1975 AND symb_decoder(16#f7#)) OR
 					(reg_q1975 AND symb_decoder(16#21#)) OR
 					(reg_q1975 AND symb_decoder(16#ce#)) OR
 					(reg_q1975 AND symb_decoder(16#48#)) OR
 					(reg_q1975 AND symb_decoder(16#52#)) OR
 					(reg_q1975 AND symb_decoder(16#71#)) OR
 					(reg_q1975 AND symb_decoder(16#a3#)) OR
 					(reg_q1975 AND symb_decoder(16#86#)) OR
 					(reg_q1975 AND symb_decoder(16#ae#)) OR
 					(reg_q1975 AND symb_decoder(16#f8#)) OR
 					(reg_q1975 AND symb_decoder(16#6d#)) OR
 					(reg_q1975 AND symb_decoder(16#13#)) OR
 					(reg_q1975 AND symb_decoder(16#f0#)) OR
 					(reg_q1975 AND symb_decoder(16#24#)) OR
 					(reg_q1975 AND symb_decoder(16#da#)) OR
 					(reg_q1975 AND symb_decoder(16#77#)) OR
 					(reg_q1975 AND symb_decoder(16#51#)) OR
 					(reg_q1975 AND symb_decoder(16#2b#)) OR
 					(reg_q1975 AND symb_decoder(16#c9#)) OR
 					(reg_q1975 AND symb_decoder(16#5c#)) OR
 					(reg_q1975 AND symb_decoder(16#7e#)) OR
 					(reg_q1975 AND symb_decoder(16#7d#)) OR
 					(reg_q1975 AND symb_decoder(16#a1#)) OR
 					(reg_q1975 AND symb_decoder(16#4e#)) OR
 					(reg_q1975 AND symb_decoder(16#a4#)) OR
 					(reg_q1975 AND symb_decoder(16#3a#)) OR
 					(reg_q1975 AND symb_decoder(16#73#)) OR
 					(reg_q1975 AND symb_decoder(16#f5#)) OR
 					(reg_q1975 AND symb_decoder(16#d9#)) OR
 					(reg_q1975 AND symb_decoder(16#e6#)) OR
 					(reg_q1975 AND symb_decoder(16#81#)) OR
 					(reg_q1975 AND symb_decoder(16#23#)) OR
 					(reg_q1975 AND symb_decoder(16#6a#)) OR
 					(reg_q1975 AND symb_decoder(16#6f#)) OR
 					(reg_q1975 AND symb_decoder(16#9d#)) OR
 					(reg_q1975 AND symb_decoder(16#9f#)) OR
 					(reg_q1975 AND symb_decoder(16#d2#)) OR
 					(reg_q1975 AND symb_decoder(16#80#)) OR
 					(reg_q1975 AND symb_decoder(16#36#)) OR
 					(reg_q1975 AND symb_decoder(16#fd#)) OR
 					(reg_q1975 AND symb_decoder(16#16#)) OR
 					(reg_q1975 AND symb_decoder(16#20#)) OR
 					(reg_q1975 AND symb_decoder(16#b4#)) OR
 					(reg_q1975 AND symb_decoder(16#1c#)) OR
 					(reg_q1975 AND symb_decoder(16#07#)) OR
 					(reg_q1975 AND symb_decoder(16#b6#)) OR
 					(reg_q1975 AND symb_decoder(16#c8#)) OR
 					(reg_q1975 AND symb_decoder(16#ea#)) OR
 					(reg_q1975 AND symb_decoder(16#ec#)) OR
 					(reg_q1975 AND symb_decoder(16#fb#)) OR
 					(reg_q1975 AND symb_decoder(16#06#)) OR
 					(reg_q1975 AND symb_decoder(16#5b#)) OR
 					(reg_q1975 AND symb_decoder(16#ef#)) OR
 					(reg_q1975 AND symb_decoder(16#28#)) OR
 					(reg_q1975 AND symb_decoder(16#d7#)) OR
 					(reg_q1975 AND symb_decoder(16#2d#)) OR
 					(reg_q1975 AND symb_decoder(16#f3#)) OR
 					(reg_q1975 AND symb_decoder(16#f6#)) OR
 					(reg_q1975 AND symb_decoder(16#68#)) OR
 					(reg_q1975 AND symb_decoder(16#70#)) OR
 					(reg_q1975 AND symb_decoder(16#e9#)) OR
 					(reg_q1975 AND symb_decoder(16#a9#)) OR
 					(reg_q1975 AND symb_decoder(16#fa#)) OR
 					(reg_q1975 AND symb_decoder(16#83#)) OR
 					(reg_q1975 AND symb_decoder(16#7c#)) OR
 					(reg_q1975 AND symb_decoder(16#17#)) OR
 					(reg_q1975 AND symb_decoder(16#3f#)) OR
 					(reg_q1975 AND symb_decoder(16#ca#)) OR
 					(reg_q1975 AND symb_decoder(16#7b#)) OR
 					(reg_q1975 AND symb_decoder(16#1b#)) OR
 					(reg_q1975 AND symb_decoder(16#14#)) OR
 					(reg_q1975 AND symb_decoder(16#63#)) OR
 					(reg_q1975 AND symb_decoder(16#42#)) OR
 					(reg_q1975 AND symb_decoder(16#31#)) OR
 					(reg_q1975 AND symb_decoder(16#8f#)) OR
 					(reg_q1975 AND symb_decoder(16#25#)) OR
 					(reg_q1975 AND symb_decoder(16#b7#)) OR
 					(reg_q1975 AND symb_decoder(16#85#)) OR
 					(reg_q1975 AND symb_decoder(16#fe#)) OR
 					(reg_q1975 AND symb_decoder(16#d4#)) OR
 					(reg_q1975 AND symb_decoder(16#dd#)) OR
 					(reg_q1975 AND symb_decoder(16#05#)) OR
 					(reg_q1975 AND symb_decoder(16#60#)) OR
 					(reg_q1975 AND symb_decoder(16#4d#)) OR
 					(reg_q1975 AND symb_decoder(16#1e#)) OR
 					(reg_q1975 AND symb_decoder(16#94#)) OR
 					(reg_q1975 AND symb_decoder(16#8e#)) OR
 					(reg_q1975 AND symb_decoder(16#e8#)) OR
 					(reg_q1975 AND symb_decoder(16#e1#)) OR
 					(reg_q1975 AND symb_decoder(16#96#)) OR
 					(reg_q1975 AND symb_decoder(16#8b#)) OR
 					(reg_q1975 AND symb_decoder(16#11#)) OR
 					(reg_q1975 AND symb_decoder(16#91#)) OR
 					(reg_q1975 AND symb_decoder(16#b8#)) OR
 					(reg_q1975 AND symb_decoder(16#65#)) OR
 					(reg_q1975 AND symb_decoder(16#46#)) OR
 					(reg_q1975 AND symb_decoder(16#5e#)) OR
 					(reg_q1975 AND symb_decoder(16#c2#)) OR
 					(reg_q1975 AND symb_decoder(16#22#)) OR
 					(reg_q1975 AND symb_decoder(16#59#)) OR
 					(reg_q1975 AND symb_decoder(16#87#)) OR
 					(reg_q1975 AND symb_decoder(16#00#)) OR
 					(reg_q1975 AND symb_decoder(16#5f#)) OR
 					(reg_q1975 AND symb_decoder(16#92#)) OR
 					(reg_q1975 AND symb_decoder(16#29#)) OR
 					(reg_q1975 AND symb_decoder(16#8d#)) OR
 					(reg_q1975 AND symb_decoder(16#cb#)) OR
 					(reg_q1975 AND symb_decoder(16#ee#)) OR
 					(reg_q1975 AND symb_decoder(16#78#)) OR
 					(reg_q1975 AND symb_decoder(16#95#)) OR
 					(reg_q1975 AND symb_decoder(16#9b#)) OR
 					(reg_q1975 AND symb_decoder(16#27#)) OR
 					(reg_q1975 AND symb_decoder(16#76#)) OR
 					(reg_q1975 AND symb_decoder(16#61#)) OR
 					(reg_q1975 AND symb_decoder(16#e7#)) OR
 					(reg_q1975 AND symb_decoder(16#93#)) OR
 					(reg_q1975 AND symb_decoder(16#e4#)) OR
 					(reg_q1975 AND symb_decoder(16#9c#)) OR
 					(reg_q1975 AND symb_decoder(16#90#)) OR
 					(reg_q1975 AND symb_decoder(16#a7#)) OR
 					(reg_q1975 AND symb_decoder(16#66#)) OR
 					(reg_q1975 AND symb_decoder(16#b1#)) OR
 					(reg_q1975 AND symb_decoder(16#b2#)) OR
 					(reg_q1975 AND symb_decoder(16#0f#)) OR
 					(reg_q1975 AND symb_decoder(16#dc#)) OR
 					(reg_q1975 AND symb_decoder(16#41#)) OR
 					(reg_q1975 AND symb_decoder(16#15#)) OR
 					(reg_q1975 AND symb_decoder(16#a2#)) OR
 					(reg_q1975 AND symb_decoder(16#5d#)) OR
 					(reg_q1975 AND symb_decoder(16#62#)) OR
 					(reg_q1975 AND symb_decoder(16#7f#)) OR
 					(reg_q1975 AND symb_decoder(16#b5#)) OR
 					(reg_q1975 AND symb_decoder(16#33#)) OR
 					(reg_q1975 AND symb_decoder(16#f4#)) OR
 					(reg_q1975 AND symb_decoder(16#88#)) OR
 					(reg_q1975 AND symb_decoder(16#03#)) OR
 					(reg_q1975 AND symb_decoder(16#b0#)) OR
 					(reg_q1975 AND symb_decoder(16#75#)) OR
 					(reg_q1975 AND symb_decoder(16#c1#)) OR
 					(reg_q1975 AND symb_decoder(16#64#)) OR
 					(reg_q1975 AND symb_decoder(16#97#)) OR
 					(reg_q1975 AND symb_decoder(16#37#)) OR
 					(reg_q1975 AND symb_decoder(16#ab#)) OR
 					(reg_q1975 AND symb_decoder(16#c6#)) OR
 					(reg_q1975 AND symb_decoder(16#45#)) OR
 					(reg_q1975 AND symb_decoder(16#57#)) OR
 					(reg_q1975 AND symb_decoder(16#2c#)) OR
 					(reg_q1975 AND symb_decoder(16#7a#)) OR
 					(reg_q1975 AND symb_decoder(16#1d#)) OR
 					(reg_q1975 AND symb_decoder(16#69#)) OR
 					(reg_q1975 AND symb_decoder(16#32#)) OR
 					(reg_q1975 AND symb_decoder(16#bd#)) OR
 					(reg_q1975 AND symb_decoder(16#49#)) OR
 					(reg_q1975 AND symb_decoder(16#2e#)) OR
 					(reg_q1975 AND symb_decoder(16#ed#)) OR
 					(reg_q1975 AND symb_decoder(16#a8#)) OR
 					(reg_q1975 AND symb_decoder(16#02#)) OR
 					(reg_q1975 AND symb_decoder(16#aa#)) OR
 					(reg_q1975 AND symb_decoder(16#53#)) OR
 					(reg_q1975 AND symb_decoder(16#01#)) OR
 					(reg_q1975 AND symb_decoder(16#e5#)) OR
 					(reg_q1975 AND symb_decoder(16#d1#)) OR
 					(reg_q1975 AND symb_decoder(16#79#)) OR
 					(reg_q1975 AND symb_decoder(16#c3#)) OR
 					(reg_q1975 AND symb_decoder(16#c0#)) OR
 					(reg_q1975 AND symb_decoder(16#10#)) OR
 					(reg_q1975 AND symb_decoder(16#34#)) OR
 					(reg_q1975 AND symb_decoder(16#9a#)) OR
 					(reg_q1975 AND symb_decoder(16#a0#)) OR
 					(reg_q1975 AND symb_decoder(16#1f#)) OR
 					(reg_q1975 AND symb_decoder(16#e3#)) OR
 					(reg_q1975 AND symb_decoder(16#a5#)) OR
 					(reg_q1975 AND symb_decoder(16#12#)) OR
 					(reg_q1975 AND symb_decoder(16#6e#)) OR
 					(reg_q1975 AND symb_decoder(16#26#)) OR
 					(reg_q1975 AND symb_decoder(16#18#)) OR
 					(reg_q1975 AND symb_decoder(16#1a#)) OR
 					(reg_q1975 AND symb_decoder(16#58#)) OR
 					(reg_q1975 AND symb_decoder(16#c7#)) OR
 					(reg_q1975 AND symb_decoder(16#67#)) OR
 					(reg_q1975 AND symb_decoder(16#2a#)) OR
 					(reg_q1975 AND symb_decoder(16#3d#)) OR
 					(reg_q1975 AND symb_decoder(16#6c#)) OR
 					(reg_q1975 AND symb_decoder(16#cc#)) OR
 					(reg_q1975 AND symb_decoder(16#e2#)) OR
 					(reg_q1975 AND symb_decoder(16#8c#)) OR
 					(reg_q1975 AND symb_decoder(16#0b#)) OR
 					(reg_q1975 AND symb_decoder(16#f9#)) OR
 					(reg_q1975 AND symb_decoder(16#de#)) OR
 					(reg_q1975 AND symb_decoder(16#c5#)) OR
 					(reg_q1975 AND symb_decoder(16#bb#)) OR
 					(reg_q1975 AND symb_decoder(16#55#)) OR
 					(reg_q1975 AND symb_decoder(16#04#)) OR
 					(reg_q1975 AND symb_decoder(16#bc#)) OR
 					(reg_q1975 AND symb_decoder(16#df#)) OR
 					(reg_q1975 AND symb_decoder(16#d5#)) OR
 					(reg_q1975 AND symb_decoder(16#3c#)) OR
 					(reg_q1975 AND symb_decoder(16#b9#)) OR
 					(reg_q1975 AND symb_decoder(16#72#)) OR
 					(reg_q1975 AND symb_decoder(16#40#)) OR
 					(reg_q1975 AND symb_decoder(16#30#)) OR
 					(reg_q1975 AND symb_decoder(16#39#)) OR
 					(reg_q1975 AND symb_decoder(16#98#)) OR
 					(reg_q1975 AND symb_decoder(16#0c#)) OR
 					(reg_q1975 AND symb_decoder(16#e0#)) OR
 					(reg_q1975 AND symb_decoder(16#2f#)) OR
 					(reg_q1975 AND symb_decoder(16#4b#)) OR
 					(reg_q1975 AND symb_decoder(16#09#)) OR
 					(reg_q1975 AND symb_decoder(16#f2#)) OR
 					(reg_q1975 AND symb_decoder(16#89#)) OR
 					(reg_q1975 AND symb_decoder(16#c4#)) OR
 					(reg_q1975 AND symb_decoder(16#99#)) OR
 					(reg_q1975 AND symb_decoder(16#4c#)) OR
 					(reg_q1975 AND symb_decoder(16#fc#)) OR
 					(reg_q1975 AND symb_decoder(16#ac#)) OR
 					(reg_q1975 AND symb_decoder(16#d3#)) OR
 					(reg_q1975 AND symb_decoder(16#4f#)) OR
 					(reg_q1975 AND symb_decoder(16#84#)) OR
 					(reg_q1975 AND symb_decoder(16#ba#)) OR
 					(reg_q1975 AND symb_decoder(16#d0#)) OR
 					(reg_q1975 AND symb_decoder(16#56#)) OR
 					(reg_q1975 AND symb_decoder(16#cd#)) OR
 					(reg_q1975 AND symb_decoder(16#54#)) OR
 					(reg_q1975 AND symb_decoder(16#db#)) OR
 					(reg_q1975 AND symb_decoder(16#47#)) OR
 					(reg_q1975 AND symb_decoder(16#38#)) OR
 					(reg_q1975 AND symb_decoder(16#f1#)) OR
 					(reg_q1975 AND symb_decoder(16#82#)) OR
 					(reg_q1975 AND symb_decoder(16#19#)) OR
 					(reg_q1975 AND symb_decoder(16#50#)) OR
 					(reg_q1975 AND symb_decoder(16#d6#)) OR
 					(reg_q1975 AND symb_decoder(16#08#)) OR
 					(reg_q1975 AND symb_decoder(16#3e#)) OR
 					(reg_q1975 AND symb_decoder(16#eb#)) OR
 					(reg_q1975 AND symb_decoder(16#af#)) OR
 					(reg_q1975 AND symb_decoder(16#44#)) OR
 					(reg_q1975 AND symb_decoder(16#a6#)) OR
 					(reg_q1975 AND symb_decoder(16#74#));
reg_q2302_in <= (reg_q2302 AND symb_decoder(16#0a#)) OR
 					(reg_q2302 AND symb_decoder(16#0d#)) OR
 					(reg_q2302 AND symb_decoder(16#09#)) OR
 					(reg_q2302 AND symb_decoder(16#0c#)) OR
 					(reg_q2302 AND symb_decoder(16#20#)) OR
 					(reg_q2300 AND symb_decoder(16#0a#)) OR
 					(reg_q2300 AND symb_decoder(16#09#)) OR
 					(reg_q2300 AND symb_decoder(16#20#)) OR
 					(reg_q2300 AND symb_decoder(16#0c#)) OR
 					(reg_q2300 AND symb_decoder(16#0d#));
reg_q361_in <= (reg_q359 AND symb_decoder(16#72#)) OR
 					(reg_q359 AND symb_decoder(16#52#));
reg_q363_in <= (reg_q361 AND symb_decoder(16#0a#)) OR
 					(reg_q361 AND symb_decoder(16#0d#)) OR
 					(reg_q361 AND symb_decoder(16#20#)) OR
 					(reg_q361 AND symb_decoder(16#0c#)) OR
 					(reg_q361 AND symb_decoder(16#09#)) OR
 					(reg_q363 AND symb_decoder(16#0d#)) OR
 					(reg_q363 AND symb_decoder(16#0a#)) OR
 					(reg_q363 AND symb_decoder(16#20#)) OR
 					(reg_q363 AND symb_decoder(16#0c#)) OR
 					(reg_q363 AND symb_decoder(16#09#));
reg_q1104_in <= (reg_q1102 AND symb_decoder(16#54#)) OR
 					(reg_q1102 AND symb_decoder(16#74#));
reg_q1106_in <= (reg_q1104 AND symb_decoder(16#0c#)) OR
 					(reg_q1104 AND symb_decoder(16#0d#)) OR
 					(reg_q1104 AND symb_decoder(16#09#)) OR
 					(reg_q1104 AND symb_decoder(16#0a#)) OR
 					(reg_q1104 AND symb_decoder(16#20#)) OR
 					(reg_q1106 AND symb_decoder(16#0d#)) OR
 					(reg_q1106 AND symb_decoder(16#0a#)) OR
 					(reg_q1106 AND symb_decoder(16#0c#)) OR
 					(reg_q1106 AND symb_decoder(16#09#)) OR
 					(reg_q1106 AND symb_decoder(16#20#));
reg_q1668_in <= (reg_q1666 AND symb_decoder(16#2e#));
reg_q1670_in <= (reg_q1668 AND symb_decoder(16#35#)) OR
 					(reg_q1668 AND symb_decoder(16#34#)) OR
 					(reg_q1668 AND symb_decoder(16#38#)) OR
 					(reg_q1668 AND symb_decoder(16#31#)) OR
 					(reg_q1668 AND symb_decoder(16#30#)) OR
 					(reg_q1668 AND symb_decoder(16#36#)) OR
 					(reg_q1668 AND symb_decoder(16#33#)) OR
 					(reg_q1668 AND symb_decoder(16#39#)) OR
 					(reg_q1668 AND symb_decoder(16#37#)) OR
 					(reg_q1668 AND symb_decoder(16#32#)) OR
 					(reg_q1670 AND symb_decoder(16#36#)) OR
 					(reg_q1670 AND symb_decoder(16#37#)) OR
 					(reg_q1670 AND symb_decoder(16#39#)) OR
 					(reg_q1670 AND symb_decoder(16#30#)) OR
 					(reg_q1670 AND symb_decoder(16#32#)) OR
 					(reg_q1670 AND symb_decoder(16#34#)) OR
 					(reg_q1670 AND symb_decoder(16#31#)) OR
 					(reg_q1670 AND symb_decoder(16#35#)) OR
 					(reg_q1670 AND symb_decoder(16#38#)) OR
 					(reg_q1670 AND symb_decoder(16#33#));
reg_q2351_in <= (reg_q2351 AND symb_decoder(16#0d#)) OR
 					(reg_q2351 AND symb_decoder(16#0a#)) OR
 					(reg_q2351 AND symb_decoder(16#09#)) OR
 					(reg_q2351 AND symb_decoder(16#0c#)) OR
 					(reg_q2351 AND symb_decoder(16#20#)) OR
 					(reg_q2349 AND symb_decoder(16#0d#)) OR
 					(reg_q2349 AND symb_decoder(16#09#)) OR
 					(reg_q2349 AND symb_decoder(16#0c#)) OR
 					(reg_q2349 AND symb_decoder(16#20#)) OR
 					(reg_q2349 AND symb_decoder(16#0a#));
reg_q420_in <= (reg_q418 AND symb_decoder(16#61#)) OR
 					(reg_q418 AND symb_decoder(16#41#));
reg_q422_in <= (reg_q420 AND symb_decoder(16#64#)) OR
 					(reg_q420 AND symb_decoder(16#44#));
reg_q1147_in <= (reg_q1147 AND symb_decoder(16#39#)) OR
 					(reg_q1147 AND symb_decoder(16#32#)) OR
 					(reg_q1147 AND symb_decoder(16#30#)) OR
 					(reg_q1147 AND symb_decoder(16#33#)) OR
 					(reg_q1147 AND symb_decoder(16#36#)) OR
 					(reg_q1147 AND symb_decoder(16#35#)) OR
 					(reg_q1147 AND symb_decoder(16#34#)) OR
 					(reg_q1147 AND symb_decoder(16#37#)) OR
 					(reg_q1147 AND symb_decoder(16#31#)) OR
 					(reg_q1147 AND symb_decoder(16#38#)) OR
 					(reg_q1145 AND symb_decoder(16#32#)) OR
 					(reg_q1145 AND symb_decoder(16#39#)) OR
 					(reg_q1145 AND symb_decoder(16#34#)) OR
 					(reg_q1145 AND symb_decoder(16#31#)) OR
 					(reg_q1145 AND symb_decoder(16#30#)) OR
 					(reg_q1145 AND symb_decoder(16#38#)) OR
 					(reg_q1145 AND symb_decoder(16#36#)) OR
 					(reg_q1145 AND symb_decoder(16#35#)) OR
 					(reg_q1145 AND symb_decoder(16#37#)) OR
 					(reg_q1145 AND symb_decoder(16#33#));
reg_q982_in <= (reg_q980 AND symb_decoder(16#54#)) OR
 					(reg_q980 AND symb_decoder(16#74#));
reg_q984_in <= (reg_q982 AND symb_decoder(16#6f#)) OR
 					(reg_q982 AND symb_decoder(16#4f#));
reg_q1299_in <= (reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1298 AND symb_decoder(16#67#)) OR
 					(reg_q1298 AND symb_decoder(16#47#));
reg_q2603_in <= (reg_q2601 AND symb_decoder(16#75#)) OR
 					(reg_q2601 AND symb_decoder(16#55#));
reg_q2605_in <= (reg_q2603 AND symb_decoder(16#53#)) OR
 					(reg_q2603 AND symb_decoder(16#73#));
reg_q2172_in <= (reg_q2170 AND symb_decoder(16#4e#)) OR
 					(reg_q2170 AND symb_decoder(16#6e#));
reg_q2274_in <= (reg_q2272 AND symb_decoder(16#52#)) OR
 					(reg_q2272 AND symb_decoder(16#72#));
reg_q2276_in <= (reg_q2274 AND symb_decoder(16#6f#)) OR
 					(reg_q2274 AND symb_decoder(16#4f#));
reg_q1035_in <= (reg_q1035 AND symb_decoder(16#0d#)) OR
 					(reg_q1035 AND symb_decoder(16#0a#)) OR
 					(reg_q1035 AND symb_decoder(16#09#)) OR
 					(reg_q1035 AND symb_decoder(16#20#)) OR
 					(reg_q1035 AND symb_decoder(16#0c#)) OR
 					(reg_q1033 AND symb_decoder(16#0a#)) OR
 					(reg_q1033 AND symb_decoder(16#09#)) OR
 					(reg_q1033 AND symb_decoder(16#0d#)) OR
 					(reg_q1033 AND symb_decoder(16#20#)) OR
 					(reg_q1033 AND symb_decoder(16#0c#));
reg_q1037_in <= (reg_q1035 AND symb_decoder(16#73#)) OR
 					(reg_q1035 AND symb_decoder(16#53#));
reg_q671_in <= (reg_q669 AND symb_decoder(16#66#)) OR
 					(reg_q669 AND symb_decoder(16#46#));
reg_q673_in <= (reg_q671 AND symb_decoder(16#6b#)) OR
 					(reg_q671 AND symb_decoder(16#64#)) OR
 					(reg_q671 AND symb_decoder(16#57#)) OR
 					(reg_q671 AND symb_decoder(16#50#)) OR
 					(reg_q671 AND symb_decoder(16#47#)) OR
 					(reg_q671 AND symb_decoder(16#44#)) OR
 					(reg_q671 AND symb_decoder(16#73#)) OR
 					(reg_q671 AND symb_decoder(16#79#)) OR
 					(reg_q671 AND symb_decoder(16#6f#)) OR
 					(reg_q671 AND symb_decoder(16#43#)) OR
 					(reg_q671 AND symb_decoder(16#78#)) OR
 					(reg_q671 AND symb_decoder(16#6c#)) OR
 					(reg_q671 AND symb_decoder(16#75#)) OR
 					(reg_q671 AND symb_decoder(16#4e#)) OR
 					(reg_q671 AND symb_decoder(16#71#)) OR
 					(reg_q671 AND symb_decoder(16#53#)) OR
 					(reg_q671 AND symb_decoder(16#4c#)) OR
 					(reg_q671 AND symb_decoder(16#63#)) OR
 					(reg_q671 AND symb_decoder(16#74#)) OR
 					(reg_q671 AND symb_decoder(16#4a#)) OR
 					(reg_q671 AND symb_decoder(16#6d#)) OR
 					(reg_q671 AND symb_decoder(16#77#)) OR
 					(reg_q671 AND symb_decoder(16#72#)) OR
 					(reg_q671 AND symb_decoder(16#67#)) OR
 					(reg_q671 AND symb_decoder(16#55#)) OR
 					(reg_q671 AND symb_decoder(16#69#)) OR
 					(reg_q671 AND symb_decoder(16#61#)) OR
 					(reg_q671 AND symb_decoder(16#65#)) OR
 					(reg_q671 AND symb_decoder(16#5a#)) OR
 					(reg_q671 AND symb_decoder(16#56#)) OR
 					(reg_q671 AND symb_decoder(16#46#)) OR
 					(reg_q671 AND symb_decoder(16#52#)) OR
 					(reg_q671 AND symb_decoder(16#49#)) OR
 					(reg_q671 AND symb_decoder(16#42#)) OR
 					(reg_q671 AND symb_decoder(16#41#)) OR
 					(reg_q671 AND symb_decoder(16#58#)) OR
 					(reg_q671 AND symb_decoder(16#45#)) OR
 					(reg_q671 AND symb_decoder(16#48#)) OR
 					(reg_q671 AND symb_decoder(16#76#)) OR
 					(reg_q671 AND symb_decoder(16#6e#)) OR
 					(reg_q671 AND symb_decoder(16#59#)) OR
 					(reg_q671 AND symb_decoder(16#4b#)) OR
 					(reg_q671 AND symb_decoder(16#54#)) OR
 					(reg_q671 AND symb_decoder(16#6a#)) OR
 					(reg_q671 AND symb_decoder(16#70#)) OR
 					(reg_q671 AND symb_decoder(16#4d#)) OR
 					(reg_q671 AND symb_decoder(16#68#)) OR
 					(reg_q671 AND symb_decoder(16#66#)) OR
 					(reg_q671 AND symb_decoder(16#4f#)) OR
 					(reg_q671 AND symb_decoder(16#7a#)) OR
 					(reg_q671 AND symb_decoder(16#51#)) OR
 					(reg_q671 AND symb_decoder(16#62#));
reg_q1478_in <= (reg_q1476 AND symb_decoder(16#64#)) OR
 					(reg_q1476 AND symb_decoder(16#44#));
reg_q1480_in <= (reg_q1478 AND symb_decoder(16#79#)) OR
 					(reg_q1478 AND symb_decoder(16#59#));
reg_q2018_in <= (reg_q2016 AND symb_decoder(16#45#)) OR
 					(reg_q2016 AND symb_decoder(16#65#));
reg_q2020_in <= (reg_q2018 AND symb_decoder(16#72#)) OR
 					(reg_q2018 AND symb_decoder(16#52#));
reg_q1527_in <= (reg_q1525 AND symb_decoder(16#74#)) OR
 					(reg_q1525 AND symb_decoder(16#54#));
reg_q1529_in <= (reg_q1527 AND symb_decoder(16#62#)) OR
 					(reg_q1527 AND symb_decoder(16#42#));
reg_q1301_in <= (reg_q1299 AND symb_decoder(16#49#)) OR
 					(reg_q1299 AND symb_decoder(16#69#));
reg_q1660_in <= (reg_q1660 AND symb_decoder(16#0a#)) OR
 					(reg_q1660 AND symb_decoder(16#20#)) OR
 					(reg_q1660 AND symb_decoder(16#0c#)) OR
 					(reg_q1660 AND symb_decoder(16#0d#)) OR
 					(reg_q1660 AND symb_decoder(16#09#)) OR
 					(reg_q1658 AND symb_decoder(16#0c#)) OR
 					(reg_q1658 AND symb_decoder(16#0a#)) OR
 					(reg_q1658 AND symb_decoder(16#0d#)) OR
 					(reg_q1658 AND symb_decoder(16#20#)) OR
 					(reg_q1658 AND symb_decoder(16#09#));
reg_q1662_in <= (reg_q1660 AND symb_decoder(16#76#)) OR
 					(reg_q1660 AND symb_decoder(16#56#));
reg_q1441_in <= (reg_q1439 AND symb_decoder(16#59#)) OR
 					(reg_q1439 AND symb_decoder(16#79#));
reg_q1443_in <= (reg_q1441 AND symb_decoder(16#73#)) OR
 					(reg_q1441 AND symb_decoder(16#53#));
reg_q2353_in <= (reg_q2351 AND symb_decoder(16#4d#)) OR
 					(reg_q2351 AND symb_decoder(16#6d#));
reg_q2278_in <= (reg_q2276 AND symb_decoder(16#0c#)) OR
 					(reg_q2276 AND symb_decoder(16#20#)) OR
 					(reg_q2276 AND symb_decoder(16#0d#)) OR
 					(reg_q2276 AND symb_decoder(16#09#)) OR
 					(reg_q2276 AND symb_decoder(16#0a#)) OR
 					(reg_q2278 AND symb_decoder(16#09#)) OR
 					(reg_q2278 AND symb_decoder(16#0a#)) OR
 					(reg_q2278 AND symb_decoder(16#0c#)) OR
 					(reg_q2278 AND symb_decoder(16#0d#)) OR
 					(reg_q2278 AND symb_decoder(16#20#));
reg_q1027_in <= (reg_q1027 AND symb_decoder(16#09#)) OR
 					(reg_q1027 AND symb_decoder(16#0d#)) OR
 					(reg_q1027 AND symb_decoder(16#0c#)) OR
 					(reg_q1027 AND symb_decoder(16#20#)) OR
 					(reg_q1027 AND symb_decoder(16#0a#)) OR
 					(reg_q1025 AND symb_decoder(16#0d#)) OR
 					(reg_q1025 AND symb_decoder(16#0c#)) OR
 					(reg_q1025 AND symb_decoder(16#09#)) OR
 					(reg_q1025 AND symb_decoder(16#20#)) OR
 					(reg_q1025 AND symb_decoder(16#0a#));
reg_q1029_in <= (reg_q1027 AND symb_decoder(16#73#)) OR
 					(reg_q1027 AND symb_decoder(16#53#));
reg_q1084_in <= (reg_q1084 AND symb_decoder(16#0a#)) OR
 					(reg_q1084 AND symb_decoder(16#20#)) OR
 					(reg_q1084 AND symb_decoder(16#0c#)) OR
 					(reg_q1084 AND symb_decoder(16#0d#)) OR
 					(reg_q1084 AND symb_decoder(16#09#)) OR
 					(reg_q1082 AND symb_decoder(16#20#)) OR
 					(reg_q1082 AND symb_decoder(16#0d#)) OR
 					(reg_q1082 AND symb_decoder(16#09#)) OR
 					(reg_q1082 AND symb_decoder(16#0c#)) OR
 					(reg_q1082 AND symb_decoder(16#0a#));
reg_q1086_in <= (reg_q1084 AND symb_decoder(16#38#)) OR
 					(reg_q1084 AND symb_decoder(16#35#)) OR
 					(reg_q1084 AND symb_decoder(16#39#)) OR
 					(reg_q1084 AND symb_decoder(16#30#)) OR
 					(reg_q1084 AND symb_decoder(16#36#)) OR
 					(reg_q1084 AND symb_decoder(16#34#)) OR
 					(reg_q1084 AND symb_decoder(16#31#)) OR
 					(reg_q1084 AND symb_decoder(16#37#)) OR
 					(reg_q1084 AND symb_decoder(16#33#)) OR
 					(reg_q1084 AND symb_decoder(16#32#)) OR
 					(reg_q1086 AND symb_decoder(16#35#)) OR
 					(reg_q1086 AND symb_decoder(16#30#)) OR
 					(reg_q1086 AND symb_decoder(16#38#)) OR
 					(reg_q1086 AND symb_decoder(16#37#)) OR
 					(reg_q1086 AND symb_decoder(16#33#)) OR
 					(reg_q1086 AND symb_decoder(16#31#)) OR
 					(reg_q1086 AND symb_decoder(16#39#)) OR
 					(reg_q1086 AND symb_decoder(16#34#)) OR
 					(reg_q1086 AND symb_decoder(16#32#)) OR
 					(reg_q1086 AND symb_decoder(16#36#));
reg_q2514_in <= (reg_q2512 AND symb_decoder(16#2a#));
reg_q2516_in <= (reg_q2514 AND symb_decoder(16#36#)) OR
 					(reg_q2514 AND symb_decoder(16#38#)) OR
 					(reg_q2514 AND symb_decoder(16#39#)) OR
 					(reg_q2514 AND symb_decoder(16#37#)) OR
 					(reg_q2514 AND symb_decoder(16#32#)) OR
 					(reg_q2514 AND symb_decoder(16#33#)) OR
 					(reg_q2514 AND symb_decoder(16#30#)) OR
 					(reg_q2514 AND symb_decoder(16#34#)) OR
 					(reg_q2514 AND symb_decoder(16#31#)) OR
 					(reg_q2514 AND symb_decoder(16#35#)) OR
 					(reg_q2516 AND symb_decoder(16#34#)) OR
 					(reg_q2516 AND symb_decoder(16#39#)) OR
 					(reg_q2516 AND symb_decoder(16#37#)) OR
 					(reg_q2516 AND symb_decoder(16#30#)) OR
 					(reg_q2516 AND symb_decoder(16#35#)) OR
 					(reg_q2516 AND symb_decoder(16#36#)) OR
 					(reg_q2516 AND symb_decoder(16#31#)) OR
 					(reg_q2516 AND symb_decoder(16#33#)) OR
 					(reg_q2516 AND symb_decoder(16#32#)) OR
 					(reg_q2516 AND symb_decoder(16#38#));
reg_q1724_in <= (reg_q1722 AND symb_decoder(16#4f#)) OR
 					(reg_q1722 AND symb_decoder(16#6f#));
reg_q1726_in <= (reg_q1724 AND symb_decoder(16#75#)) OR
 					(reg_q1724 AND symb_decoder(16#55#));
reg_q1335_in <= (reg_q1333 AND symb_decoder(16#35#)) OR
 					(reg_q1333 AND symb_decoder(16#38#)) OR
 					(reg_q1333 AND symb_decoder(16#32#)) OR
 					(reg_q1333 AND symb_decoder(16#33#)) OR
 					(reg_q1333 AND symb_decoder(16#34#)) OR
 					(reg_q1333 AND symb_decoder(16#37#)) OR
 					(reg_q1333 AND symb_decoder(16#31#)) OR
 					(reg_q1333 AND symb_decoder(16#30#)) OR
 					(reg_q1333 AND symb_decoder(16#39#)) OR
 					(reg_q1333 AND symb_decoder(16#36#)) OR
 					(reg_q1335 AND symb_decoder(16#39#)) OR
 					(reg_q1335 AND symb_decoder(16#33#)) OR
 					(reg_q1335 AND symb_decoder(16#36#)) OR
 					(reg_q1335 AND symb_decoder(16#30#)) OR
 					(reg_q1335 AND symb_decoder(16#34#)) OR
 					(reg_q1335 AND symb_decoder(16#32#)) OR
 					(reg_q1335 AND symb_decoder(16#38#)) OR
 					(reg_q1335 AND symb_decoder(16#35#)) OR
 					(reg_q1335 AND symb_decoder(16#37#)) OR
 					(reg_q1335 AND symb_decoder(16#31#));
reg_q2109_in <= (reg_q2107 AND symb_decoder(16#58#)) OR
 					(reg_q2107 AND symb_decoder(16#78#));
reg_q2111_in <= (reg_q2109 AND symb_decoder(16#0d#)) OR
 					(reg_q2109 AND symb_decoder(16#09#)) OR
 					(reg_q2109 AND symb_decoder(16#20#)) OR
 					(reg_q2109 AND symb_decoder(16#0c#)) OR
 					(reg_q2109 AND symb_decoder(16#0a#)) OR
 					(reg_q2111 AND symb_decoder(16#09#)) OR
 					(reg_q2111 AND symb_decoder(16#20#)) OR
 					(reg_q2111 AND symb_decoder(16#0d#)) OR
 					(reg_q2111 AND symb_decoder(16#0c#)) OR
 					(reg_q2111 AND symb_decoder(16#0a#));
reg_q1355_in <= (reg_q1355 AND symb_decoder(16#0c#)) OR
 					(reg_q1355 AND symb_decoder(16#0d#)) OR
 					(reg_q1355 AND symb_decoder(16#09#)) OR
 					(reg_q1355 AND symb_decoder(16#0a#)) OR
 					(reg_q1355 AND symb_decoder(16#20#)) OR
 					(reg_q1353 AND symb_decoder(16#0a#)) OR
 					(reg_q1353 AND symb_decoder(16#09#)) OR
 					(reg_q1353 AND symb_decoder(16#0d#)) OR
 					(reg_q1353 AND symb_decoder(16#0c#)) OR
 					(reg_q1353 AND symb_decoder(16#20#));
reg_q1357_in <= (reg_q1355 AND symb_decoder(16#32#)) OR
 					(reg_q1355 AND symb_decoder(16#37#)) OR
 					(reg_q1355 AND symb_decoder(16#35#)) OR
 					(reg_q1355 AND symb_decoder(16#31#)) OR
 					(reg_q1355 AND symb_decoder(16#33#)) OR
 					(reg_q1355 AND symb_decoder(16#34#)) OR
 					(reg_q1355 AND symb_decoder(16#36#)) OR
 					(reg_q1355 AND symb_decoder(16#38#)) OR
 					(reg_q1355 AND symb_decoder(16#39#)) OR
 					(reg_q1355 AND symb_decoder(16#30#));
reg_q2004_in <= (reg_q2002 AND symb_decoder(16#66#)) OR
 					(reg_q2002 AND symb_decoder(16#46#));
reg_q1191_in <= (reg_q1189 AND symb_decoder(16#6c#)) OR
 					(reg_q1189 AND symb_decoder(16#4c#));
reg_q1193_in <= (reg_q1191 AND symb_decoder(16#45#)) OR
 					(reg_q1191 AND symb_decoder(16#65#));
reg_q1580_in <= (reg_q1580 AND symb_decoder(16#36#)) OR
 					(reg_q1580 AND symb_decoder(16#38#)) OR
 					(reg_q1580 AND symb_decoder(16#37#)) OR
 					(reg_q1580 AND symb_decoder(16#34#)) OR
 					(reg_q1580 AND symb_decoder(16#31#)) OR
 					(reg_q1580 AND symb_decoder(16#35#)) OR
 					(reg_q1580 AND symb_decoder(16#30#)) OR
 					(reg_q1580 AND symb_decoder(16#33#)) OR
 					(reg_q1580 AND symb_decoder(16#32#)) OR
 					(reg_q1580 AND symb_decoder(16#39#)) OR
 					(reg_q1578 AND symb_decoder(16#39#)) OR
 					(reg_q1578 AND symb_decoder(16#36#)) OR
 					(reg_q1578 AND symb_decoder(16#31#)) OR
 					(reg_q1578 AND symb_decoder(16#35#)) OR
 					(reg_q1578 AND symb_decoder(16#37#)) OR
 					(reg_q1578 AND symb_decoder(16#30#)) OR
 					(reg_q1578 AND symb_decoder(16#38#)) OR
 					(reg_q1578 AND symb_decoder(16#32#)) OR
 					(reg_q1578 AND symb_decoder(16#34#)) OR
 					(reg_q1578 AND symb_decoder(16#33#));
reg_q824_in <= (reg_q822 AND symb_decoder(16#4e#)) OR
 					(reg_q822 AND symb_decoder(16#6e#));
reg_q826_in <= (reg_q824 AND symb_decoder(16#66#)) OR
 					(reg_q824 AND symb_decoder(16#46#));
reg_q690_in <= (reg_q688 AND symb_decoder(16#2e#));
reg_q692_in <= (reg_q690 AND symb_decoder(16#35#)) OR
 					(reg_q690 AND symb_decoder(16#30#)) OR
 					(reg_q690 AND symb_decoder(16#37#)) OR
 					(reg_q690 AND symb_decoder(16#32#)) OR
 					(reg_q690 AND symb_decoder(16#38#)) OR
 					(reg_q690 AND symb_decoder(16#36#)) OR
 					(reg_q690 AND symb_decoder(16#34#)) OR
 					(reg_q690 AND symb_decoder(16#39#)) OR
 					(reg_q690 AND symb_decoder(16#31#)) OR
 					(reg_q690 AND symb_decoder(16#33#)) OR
 					(reg_q692 AND symb_decoder(16#39#)) OR
 					(reg_q692 AND symb_decoder(16#32#)) OR
 					(reg_q692 AND symb_decoder(16#31#)) OR
 					(reg_q692 AND symb_decoder(16#37#)) OR
 					(reg_q692 AND symb_decoder(16#33#)) OR
 					(reg_q692 AND symb_decoder(16#35#)) OR
 					(reg_q692 AND symb_decoder(16#38#)) OR
 					(reg_q692 AND symb_decoder(16#34#)) OR
 					(reg_q692 AND symb_decoder(16#30#)) OR
 					(reg_q692 AND symb_decoder(16#36#));
reg_q709_in <= (reg_q707 AND symb_decoder(16#0d#)) OR
 					(reg_q707 AND symb_decoder(16#0c#)) OR
 					(reg_q707 AND symb_decoder(16#0a#)) OR
 					(reg_q707 AND symb_decoder(16#20#)) OR
 					(reg_q707 AND symb_decoder(16#09#));
reg_q711_in <= (reg_q709 AND symb_decoder(16#35#)) OR
 					(reg_q709 AND symb_decoder(16#30#)) OR
 					(reg_q709 AND symb_decoder(16#39#)) OR
 					(reg_q709 AND symb_decoder(16#36#)) OR
 					(reg_q709 AND symb_decoder(16#31#)) OR
 					(reg_q709 AND symb_decoder(16#38#)) OR
 					(reg_q709 AND symb_decoder(16#32#)) OR
 					(reg_q709 AND symb_decoder(16#34#)) OR
 					(reg_q709 AND symb_decoder(16#33#)) OR
 					(reg_q709 AND symb_decoder(16#37#)) OR
 					(reg_q711 AND symb_decoder(16#32#)) OR
 					(reg_q711 AND symb_decoder(16#36#)) OR
 					(reg_q711 AND symb_decoder(16#38#)) OR
 					(reg_q711 AND symb_decoder(16#31#)) OR
 					(reg_q711 AND symb_decoder(16#33#)) OR
 					(reg_q711 AND symb_decoder(16#30#)) OR
 					(reg_q711 AND symb_decoder(16#35#)) OR
 					(reg_q711 AND symb_decoder(16#39#)) OR
 					(reg_q711 AND symb_decoder(16#34#)) OR
 					(reg_q711 AND symb_decoder(16#37#));
reg_q373_in <= (reg_q371 AND symb_decoder(16#22#));
reg_q375_in <= (reg_q373 AND symb_decoder(16#54#)) OR
 					(reg_q373 AND symb_decoder(16#74#));
reg_q247_in <= (reg_q245 AND symb_decoder(16#ff#));
reg_q249_in <= (reg_q247 AND symb_decoder(16#38#)) OR
 					(reg_q247 AND symb_decoder(16#36#)) OR
 					(reg_q247 AND symb_decoder(16#37#)) OR
 					(reg_q247 AND symb_decoder(16#33#)) OR
 					(reg_q247 AND symb_decoder(16#32#)) OR
 					(reg_q247 AND symb_decoder(16#39#)) OR
 					(reg_q247 AND symb_decoder(16#34#)) OR
 					(reg_q247 AND symb_decoder(16#30#)) OR
 					(reg_q247 AND symb_decoder(16#31#)) OR
 					(reg_q247 AND symb_decoder(16#35#)) OR
 					(reg_q249 AND symb_decoder(16#39#)) OR
 					(reg_q249 AND symb_decoder(16#37#)) OR
 					(reg_q249 AND symb_decoder(16#34#)) OR
 					(reg_q249 AND symb_decoder(16#35#)) OR
 					(reg_q249 AND symb_decoder(16#38#)) OR
 					(reg_q249 AND symb_decoder(16#32#)) OR
 					(reg_q249 AND symb_decoder(16#30#)) OR
 					(reg_q249 AND symb_decoder(16#31#)) OR
 					(reg_q249 AND symb_decoder(16#36#)) OR
 					(reg_q249 AND symb_decoder(16#33#));
reg_q2038_in <= (reg_q2036 AND symb_decoder(16#45#)) OR
 					(reg_q2036 AND symb_decoder(16#65#));
reg_q2040_in <= (reg_q2038 AND symb_decoder(16#0d#)) OR
 					(reg_q2038 AND symb_decoder(16#09#)) OR
 					(reg_q2038 AND symb_decoder(16#0c#)) OR
 					(reg_q2038 AND symb_decoder(16#0a#)) OR
 					(reg_q2038 AND symb_decoder(16#20#)) OR
 					(reg_q2040 AND symb_decoder(16#0c#)) OR
 					(reg_q2040 AND symb_decoder(16#09#)) OR
 					(reg_q2040 AND symb_decoder(16#0d#)) OR
 					(reg_q2040 AND symb_decoder(16#0a#)) OR
 					(reg_q2040 AND symb_decoder(16#20#));
reg_q1975_in <= (reg_q1973 AND symb_decoder(16#23#));
reg_q1248_in <= (reg_q1248 AND symb_decoder(16#0d#)) OR
 					(reg_q1248 AND symb_decoder(16#0c#)) OR
 					(reg_q1248 AND symb_decoder(16#0a#)) OR
 					(reg_q1248 AND symb_decoder(16#09#)) OR
 					(reg_q1248 AND symb_decoder(16#20#)) OR
 					(reg_q1246 AND symb_decoder(16#0a#)) OR
 					(reg_q1246 AND symb_decoder(16#0d#)) OR
 					(reg_q1246 AND symb_decoder(16#09#)) OR
 					(reg_q1246 AND symb_decoder(16#20#)) OR
 					(reg_q1246 AND symb_decoder(16#0c#));
reg_q2369_in <= (reg_q2369 AND symb_decoder(16#0a#)) OR
 					(reg_q2369 AND symb_decoder(16#09#)) OR
 					(reg_q2369 AND symb_decoder(16#20#)) OR
 					(reg_q2369 AND symb_decoder(16#0d#)) OR
 					(reg_q2369 AND symb_decoder(16#0c#)) OR
 					(reg_q2367 AND symb_decoder(16#0d#)) OR
 					(reg_q2367 AND symb_decoder(16#09#)) OR
 					(reg_q2367 AND symb_decoder(16#0c#)) OR
 					(reg_q2367 AND symb_decoder(16#0a#)) OR
 					(reg_q2367 AND symb_decoder(16#20#));
reg_q1094_in <= (reg_q1092 AND symb_decoder(16#2e#));
reg_q1096_in <= (reg_q1094 AND symb_decoder(16#0d#)) OR
 					(reg_q1094 AND symb_decoder(16#20#)) OR
 					(reg_q1094 AND symb_decoder(16#0a#)) OR
 					(reg_q1094 AND symb_decoder(16#0c#)) OR
 					(reg_q1094 AND symb_decoder(16#09#)) OR
 					(reg_q1096 AND symb_decoder(16#0c#)) OR
 					(reg_q1096 AND symb_decoder(16#0d#)) OR
 					(reg_q1096 AND symb_decoder(16#20#)) OR
 					(reg_q1096 AND symb_decoder(16#09#)) OR
 					(reg_q1096 AND symb_decoder(16#0a#));
reg_q1108_in <= (reg_q1106 AND symb_decoder(16#35#)) OR
 					(reg_q1106 AND symb_decoder(16#38#)) OR
 					(reg_q1106 AND symb_decoder(16#32#)) OR
 					(reg_q1106 AND symb_decoder(16#39#)) OR
 					(reg_q1106 AND symb_decoder(16#36#)) OR
 					(reg_q1106 AND symb_decoder(16#37#)) OR
 					(reg_q1106 AND symb_decoder(16#34#)) OR
 					(reg_q1106 AND symb_decoder(16#33#)) OR
 					(reg_q1106 AND symb_decoder(16#30#)) OR
 					(reg_q1106 AND symb_decoder(16#31#)) OR
 					(reg_q1108 AND symb_decoder(16#39#)) OR
 					(reg_q1108 AND symb_decoder(16#38#)) OR
 					(reg_q1108 AND symb_decoder(16#32#)) OR
 					(reg_q1108 AND symb_decoder(16#33#)) OR
 					(reg_q1108 AND symb_decoder(16#30#)) OR
 					(reg_q1108 AND symb_decoder(16#31#)) OR
 					(reg_q1108 AND symb_decoder(16#37#)) OR
 					(reg_q1108 AND symb_decoder(16#34#)) OR
 					(reg_q1108 AND symb_decoder(16#36#)) OR
 					(reg_q1108 AND symb_decoder(16#35#));
reg_q56_in <= (reg_q54 AND symb_decoder(16#6b#)) OR
 					(reg_q54 AND symb_decoder(16#4b#));
reg_q58_in <= (reg_q56 AND symb_decoder(16#20#)) OR
 					(reg_q56 AND symb_decoder(16#0c#)) OR
 					(reg_q56 AND symb_decoder(16#0d#)) OR
 					(reg_q56 AND symb_decoder(16#09#)) OR
 					(reg_q56 AND symb_decoder(16#0a#)) OR
 					(reg_q58 AND symb_decoder(16#09#)) OR
 					(reg_q58 AND symb_decoder(16#0a#)) OR
 					(reg_q58 AND symb_decoder(16#20#)) OR
 					(reg_q58 AND symb_decoder(16#0d#)) OR
 					(reg_q58 AND symb_decoder(16#0c#));
reg_q101_in <= (reg_q99 AND symb_decoder(16#4f#)) OR
 					(reg_q99 AND symb_decoder(16#6f#));
reg_q103_in <= (reg_q101 AND symb_decoder(16#50#)) OR
 					(reg_q101 AND symb_decoder(16#70#));
reg_q2480_in <= (reg_q2478 AND symb_decoder(16#2a#));
reg_q2482_in <= (reg_q2480 AND symb_decoder(16#36#)) OR
 					(reg_q2480 AND symb_decoder(16#32#)) OR
 					(reg_q2480 AND symb_decoder(16#34#)) OR
 					(reg_q2480 AND symb_decoder(16#33#)) OR
 					(reg_q2480 AND symb_decoder(16#35#)) OR
 					(reg_q2480 AND symb_decoder(16#30#)) OR
 					(reg_q2480 AND symb_decoder(16#38#)) OR
 					(reg_q2480 AND symb_decoder(16#39#)) OR
 					(reg_q2480 AND symb_decoder(16#31#)) OR
 					(reg_q2480 AND symb_decoder(16#37#)) OR
 					(reg_q2482 AND symb_decoder(16#30#)) OR
 					(reg_q2482 AND symb_decoder(16#34#)) OR
 					(reg_q2482 AND symb_decoder(16#33#)) OR
 					(reg_q2482 AND symb_decoder(16#38#)) OR
 					(reg_q2482 AND symb_decoder(16#35#)) OR
 					(reg_q2482 AND symb_decoder(16#39#)) OR
 					(reg_q2482 AND symb_decoder(16#36#)) OR
 					(reg_q2482 AND symb_decoder(16#32#)) OR
 					(reg_q2482 AND symb_decoder(16#31#)) OR
 					(reg_q2482 AND symb_decoder(16#37#));
reg_q1482_in <= (reg_q1480 AND symb_decoder(16#09#)) OR
 					(reg_q1480 AND symb_decoder(16#0a#)) OR
 					(reg_q1480 AND symb_decoder(16#0d#)) OR
 					(reg_q1480 AND symb_decoder(16#0c#)) OR
 					(reg_q1480 AND symb_decoder(16#20#)) OR
 					(reg_q1482 AND symb_decoder(16#0a#)) OR
 					(reg_q1482 AND symb_decoder(16#20#)) OR
 					(reg_q1482 AND symb_decoder(16#09#)) OR
 					(reg_q1482 AND symb_decoder(16#0d#)) OR
 					(reg_q1482 AND symb_decoder(16#0c#));
reg_q367_in <= (reg_q365 AND symb_decoder(16#2e#));
reg_q369_in <= (reg_q367 AND symb_decoder(16#30#)) OR
 					(reg_q367 AND symb_decoder(16#39#)) OR
 					(reg_q367 AND symb_decoder(16#38#)) OR
 					(reg_q367 AND symb_decoder(16#37#)) OR
 					(reg_q367 AND symb_decoder(16#33#)) OR
 					(reg_q367 AND symb_decoder(16#35#)) OR
 					(reg_q367 AND symb_decoder(16#34#)) OR
 					(reg_q367 AND symb_decoder(16#31#)) OR
 					(reg_q367 AND symb_decoder(16#36#)) OR
 					(reg_q367 AND symb_decoder(16#32#)) OR
 					(reg_q369 AND symb_decoder(16#38#)) OR
 					(reg_q369 AND symb_decoder(16#32#)) OR
 					(reg_q369 AND symb_decoder(16#39#)) OR
 					(reg_q369 AND symb_decoder(16#31#)) OR
 					(reg_q369 AND symb_decoder(16#34#)) OR
 					(reg_q369 AND symb_decoder(16#33#)) OR
 					(reg_q369 AND symb_decoder(16#30#)) OR
 					(reg_q369 AND symb_decoder(16#35#)) OR
 					(reg_q369 AND symb_decoder(16#37#)) OR
 					(reg_q369 AND symb_decoder(16#36#));
reg_q700_in <= (reg_q700 AND symb_decoder(16#34#)) OR
 					(reg_q700 AND symb_decoder(16#33#)) OR
 					(reg_q700 AND symb_decoder(16#36#)) OR
 					(reg_q700 AND symb_decoder(16#38#)) OR
 					(reg_q700 AND symb_decoder(16#39#)) OR
 					(reg_q700 AND symb_decoder(16#31#)) OR
 					(reg_q700 AND symb_decoder(16#37#)) OR
 					(reg_q700 AND symb_decoder(16#32#)) OR
 					(reg_q700 AND symb_decoder(16#35#)) OR
 					(reg_q700 AND symb_decoder(16#30#)) OR
 					(reg_q698 AND symb_decoder(16#39#)) OR
 					(reg_q698 AND symb_decoder(16#31#)) OR
 					(reg_q698 AND symb_decoder(16#30#)) OR
 					(reg_q698 AND symb_decoder(16#35#)) OR
 					(reg_q698 AND symb_decoder(16#36#)) OR
 					(reg_q698 AND symb_decoder(16#32#)) OR
 					(reg_q698 AND symb_decoder(16#34#)) OR
 					(reg_q698 AND symb_decoder(16#37#)) OR
 					(reg_q698 AND symb_decoder(16#33#)) OR
 					(reg_q698 AND symb_decoder(16#38#));
reg_q196_in <= (reg_q194 AND symb_decoder(16#45#)) OR
 					(reg_q194 AND symb_decoder(16#65#));
reg_q198_in <= (reg_q196 AND symb_decoder(16#4e#)) OR
 					(reg_q196 AND symb_decoder(16#6e#));
reg_q418_in <= (reg_q416 AND symb_decoder(16#4c#)) OR
 					(reg_q416 AND symb_decoder(16#6c#));
reg_q1688_in <= (reg_q1686 AND symb_decoder(16#6c#)) OR
 					(reg_q1686 AND symb_decoder(16#4c#));
reg_q1690_in <= (reg_q1688 AND symb_decoder(16#6c#)) OR
 					(reg_q1688 AND symb_decoder(16#4c#));
reg_q357_in <= (reg_q355 AND symb_decoder(16#56#)) OR
 					(reg_q355 AND symb_decoder(16#76#));
reg_q359_in <= (reg_q357 AND symb_decoder(16#45#)) OR
 					(reg_q357 AND symb_decoder(16#65#));
reg_q2101_in <= (reg_q2099 AND symb_decoder(16#61#)) OR
 					(reg_q2099 AND symb_decoder(16#41#));
reg_q2103_in <= (reg_q2101 AND symb_decoder(16#0c#)) OR
 					(reg_q2101 AND symb_decoder(16#0d#)) OR
 					(reg_q2101 AND symb_decoder(16#09#)) OR
 					(reg_q2101 AND symb_decoder(16#0a#)) OR
 					(reg_q2101 AND symb_decoder(16#20#)) OR
 					(reg_q2103 AND symb_decoder(16#09#)) OR
 					(reg_q2103 AND symb_decoder(16#0d#)) OR
 					(reg_q2103 AND symb_decoder(16#0c#)) OR
 					(reg_q2103 AND symb_decoder(16#20#)) OR
 					(reg_q2103 AND symb_decoder(16#0a#));
reg_q2375_in <= (reg_q2373 AND symb_decoder(16#2e#));
reg_q2377_in <= (reg_q2375 AND symb_decoder(16#35#)) OR
 					(reg_q2375 AND symb_decoder(16#31#)) OR
 					(reg_q2375 AND symb_decoder(16#36#)) OR
 					(reg_q2375 AND symb_decoder(16#30#)) OR
 					(reg_q2375 AND symb_decoder(16#39#)) OR
 					(reg_q2375 AND symb_decoder(16#37#)) OR
 					(reg_q2375 AND symb_decoder(16#38#)) OR
 					(reg_q2375 AND symb_decoder(16#32#)) OR
 					(reg_q2375 AND symb_decoder(16#33#)) OR
 					(reg_q2375 AND symb_decoder(16#34#)) OR
 					(reg_q2377 AND symb_decoder(16#33#)) OR
 					(reg_q2377 AND symb_decoder(16#37#)) OR
 					(reg_q2377 AND symb_decoder(16#30#)) OR
 					(reg_q2377 AND symb_decoder(16#36#)) OR
 					(reg_q2377 AND symb_decoder(16#39#)) OR
 					(reg_q2377 AND symb_decoder(16#31#)) OR
 					(reg_q2377 AND symb_decoder(16#32#)) OR
 					(reg_q2377 AND symb_decoder(16#34#)) OR
 					(reg_q2377 AND symb_decoder(16#35#)) OR
 					(reg_q2377 AND symb_decoder(16#38#));
reg_q2361_in <= (reg_q2359 AND symb_decoder(16#47#)) OR
 					(reg_q2359 AND symb_decoder(16#67#));
reg_q2363_in <= (reg_q2361 AND symb_decoder(16#65#)) OR
 					(reg_q2361 AND symb_decoder(16#45#));
reg_q121_in <= (reg_q119 AND symb_decoder(16#56#)) OR
 					(reg_q119 AND symb_decoder(16#76#));
reg_q123_in <= (reg_q121 AND symb_decoder(16#34#)) OR
 					(reg_q121 AND symb_decoder(16#36#)) OR
 					(reg_q121 AND symb_decoder(16#32#)) OR
 					(reg_q121 AND symb_decoder(16#31#)) OR
 					(reg_q121 AND symb_decoder(16#33#)) OR
 					(reg_q121 AND symb_decoder(16#30#)) OR
 					(reg_q121 AND symb_decoder(16#37#)) OR
 					(reg_q121 AND symb_decoder(16#38#)) OR
 					(reg_q121 AND symb_decoder(16#39#)) OR
 					(reg_q121 AND symb_decoder(16#35#)) OR
 					(reg_q123 AND symb_decoder(16#37#)) OR
 					(reg_q123 AND symb_decoder(16#31#)) OR
 					(reg_q123 AND symb_decoder(16#35#)) OR
 					(reg_q123 AND symb_decoder(16#39#)) OR
 					(reg_q123 AND symb_decoder(16#33#)) OR
 					(reg_q123 AND symb_decoder(16#34#)) OR
 					(reg_q123 AND symb_decoder(16#36#)) OR
 					(reg_q123 AND symb_decoder(16#30#)) OR
 					(reg_q123 AND symb_decoder(16#32#)) OR
 					(reg_q123 AND symb_decoder(16#38#));
reg_q2613_in <= (reg_q2613 AND symb_decoder(16#20#)) OR
 					(reg_q2613 AND symb_decoder(16#09#)) OR
 					(reg_q2613 AND symb_decoder(16#0d#)) OR
 					(reg_q2613 AND symb_decoder(16#0a#)) OR
 					(reg_q2613 AND symb_decoder(16#0c#)) OR
 					(reg_q2611 AND symb_decoder(16#0c#)) OR
 					(reg_q2611 AND symb_decoder(16#09#)) OR
 					(reg_q2611 AND symb_decoder(16#0d#)) OR
 					(reg_q2611 AND symb_decoder(16#20#)) OR
 					(reg_q2611 AND symb_decoder(16#0a#));
reg_q818_in <= (reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q817 AND symb_decoder(16#44#)) OR
 					(reg_q817 AND symb_decoder(16#64#));
reg_q2593_in <= (reg_q2591 AND symb_decoder(16#72#)) OR
 					(reg_q2591 AND symb_decoder(16#52#));
reg_q2595_in <= (reg_q2593 AND symb_decoder(16#65#)) OR
 					(reg_q2593 AND symb_decoder(16#45#));
reg_q426_in <= (reg_q426 AND symb_decoder(16#0a#)) OR
 					(reg_q426 AND symb_decoder(16#20#)) OR
 					(reg_q426 AND symb_decoder(16#0c#)) OR
 					(reg_q426 AND symb_decoder(16#09#)) OR
 					(reg_q426 AND symb_decoder(16#0d#)) OR
 					(reg_q424 AND symb_decoder(16#0a#)) OR
 					(reg_q424 AND symb_decoder(16#0d#)) OR
 					(reg_q424 AND symb_decoder(16#20#)) OR
 					(reg_q424 AND symb_decoder(16#09#)) OR
 					(reg_q424 AND symb_decoder(16#0c#));
reg_q428_in <= (reg_q426 AND symb_decoder(16#72#)) OR
 					(reg_q426 AND symb_decoder(16#52#));
reg_q2337_in <= (reg_q2337 AND symb_decoder(16#09#)) OR
 					(reg_q2337 AND symb_decoder(16#20#)) OR
 					(reg_q2337 AND symb_decoder(16#0c#)) OR
 					(reg_q2337 AND symb_decoder(16#0a#)) OR
 					(reg_q2337 AND symb_decoder(16#0d#)) OR
 					(reg_q2335 AND symb_decoder(16#09#)) OR
 					(reg_q2335 AND symb_decoder(16#0c#)) OR
 					(reg_q2335 AND symb_decoder(16#0d#)) OR
 					(reg_q2335 AND symb_decoder(16#20#)) OR
 					(reg_q2335 AND symb_decoder(16#0a#));
reg_q127_in <= (reg_q127 AND symb_decoder(16#33#)) OR
 					(reg_q127 AND symb_decoder(16#38#)) OR
 					(reg_q127 AND symb_decoder(16#39#)) OR
 					(reg_q127 AND symb_decoder(16#37#)) OR
 					(reg_q127 AND symb_decoder(16#31#)) OR
 					(reg_q127 AND symb_decoder(16#36#)) OR
 					(reg_q127 AND symb_decoder(16#30#)) OR
 					(reg_q127 AND symb_decoder(16#34#)) OR
 					(reg_q127 AND symb_decoder(16#35#)) OR
 					(reg_q127 AND symb_decoder(16#32#)) OR
 					(reg_q125 AND symb_decoder(16#31#)) OR
 					(reg_q125 AND symb_decoder(16#32#)) OR
 					(reg_q125 AND symb_decoder(16#30#)) OR
 					(reg_q125 AND symb_decoder(16#34#)) OR
 					(reg_q125 AND symb_decoder(16#38#)) OR
 					(reg_q125 AND symb_decoder(16#33#)) OR
 					(reg_q125 AND symb_decoder(16#39#)) OR
 					(reg_q125 AND symb_decoder(16#36#)) OR
 					(reg_q125 AND symb_decoder(16#37#)) OR
 					(reg_q125 AND symb_decoder(16#35#));
reg_q1337_in <= (reg_q1335 AND symb_decoder(16#2e#));
reg_q2341_in <= (reg_q2339 AND symb_decoder(16#45#)) OR
 					(reg_q2339 AND symb_decoder(16#65#));
reg_q2343_in <= (reg_q2341 AND symb_decoder(16#4d#)) OR
 					(reg_q2341 AND symb_decoder(16#6d#));
reg_q966_in <= (reg_q964 AND symb_decoder(16#57#)) OR
 					(reg_q964 AND symb_decoder(16#77#));
reg_q968_in <= (reg_q966 AND symb_decoder(16#45#)) OR
 					(reg_q966 AND symb_decoder(16#65#));
reg_q1676_in <= (reg_q1674 AND symb_decoder(16#66#)) OR
 					(reg_q1674 AND symb_decoder(16#46#));
reg_q1678_in <= (reg_q1676 AND symb_decoder(16#69#)) OR
 					(reg_q1676 AND symb_decoder(16#49#));
reg_q379_in <= (reg_q377 AND symb_decoder(16#45#)) OR
 					(reg_q377 AND symb_decoder(16#65#));
reg_q381_in <= (reg_q379 AND symb_decoder(16#0d#)) OR
 					(reg_q379 AND symb_decoder(16#0c#)) OR
 					(reg_q379 AND symb_decoder(16#0a#)) OR
 					(reg_q379 AND symb_decoder(16#20#)) OR
 					(reg_q379 AND symb_decoder(16#09#)) OR
 					(reg_q381 AND symb_decoder(16#20#)) OR
 					(reg_q381 AND symb_decoder(16#0d#)) OR
 					(reg_q381 AND symb_decoder(16#0c#)) OR
 					(reg_q381 AND symb_decoder(16#09#)) OR
 					(reg_q381 AND symb_decoder(16#0a#));
reg_q2577_in <= (reg_q2575 AND symb_decoder(16#3a#));
reg_q2688_in <= (reg_q2686 AND symb_decoder(16#64#)) OR
 					(reg_q2686 AND symb_decoder(16#44#));
reg_q2690_in <= (reg_q2688 AND symb_decoder(16#5c#));
reg_q1531_in <= (reg_q1529 AND symb_decoder(16#75#)) OR
 					(reg_q1529 AND symb_decoder(16#55#));
reg_q1674_in <= (reg_q1674 AND symb_decoder(16#0a#)) OR
 					(reg_q1674 AND symb_decoder(16#0d#)) OR
 					(reg_q1674 AND symb_decoder(16#09#)) OR
 					(reg_q1674 AND symb_decoder(16#20#)) OR
 					(reg_q1674 AND symb_decoder(16#0c#)) OR
 					(reg_q1672 AND symb_decoder(16#09#)) OR
 					(reg_q1672 AND symb_decoder(16#20#)) OR
 					(reg_q1672 AND symb_decoder(16#0a#)) OR
 					(reg_q1672 AND symb_decoder(16#0d#)) OR
 					(reg_q1672 AND symb_decoder(16#0c#));
reg_q756_in <= (reg_q756 AND symb_decoder(16#09#)) OR
 					(reg_q756 AND symb_decoder(16#20#)) OR
 					(reg_q756 AND symb_decoder(16#0d#)) OR
 					(reg_q756 AND symb_decoder(16#0a#)) OR
 					(reg_q756 AND symb_decoder(16#0c#)) OR
 					(reg_q754 AND symb_decoder(16#0c#)) OR
 					(reg_q754 AND symb_decoder(16#0a#)) OR
 					(reg_q754 AND symb_decoder(16#0d#)) OR
 					(reg_q754 AND symb_decoder(16#09#)) OR
 					(reg_q754 AND symb_decoder(16#20#));
reg_q1305_in <= (reg_q1303 AND symb_decoder(16#4c#)) OR
 					(reg_q1303 AND symb_decoder(16#6c#));
reg_q1307_in <= (reg_q1305 AND symb_decoder(16#66#)) OR
 					(reg_q1305 AND symb_decoder(16#46#));
reg_q1425_in <= (reg_q1423 AND symb_decoder(16#52#)) OR
 					(reg_q1423 AND symb_decoder(16#72#));
reg_q1427_in <= (reg_q1425 AND symb_decoder(16#41#)) OR
 					(reg_q1425 AND symb_decoder(16#61#));
reg_q194_in <= (reg_q192 AND symb_decoder(16#47#)) OR
 					(reg_q192 AND symb_decoder(16#67#));
reg_q115_in <= (reg_q113 AND symb_decoder(16#72#)) OR
 					(reg_q113 AND symb_decoder(16#52#));
reg_q117_in <= (reg_q115 AND symb_decoder(16#4f#)) OR
 					(reg_q115 AND symb_decoder(16#6f#));
reg_q1250_in <= (reg_q1248 AND symb_decoder(16#76#)) OR
 					(reg_q1248 AND symb_decoder(16#56#));
reg_q1252_in <= (reg_q1250 AND symb_decoder(16#36#)) OR
 					(reg_q1250 AND symb_decoder(16#37#)) OR
 					(reg_q1250 AND symb_decoder(16#31#)) OR
 					(reg_q1250 AND symb_decoder(16#34#)) OR
 					(reg_q1250 AND symb_decoder(16#32#)) OR
 					(reg_q1250 AND symb_decoder(16#35#)) OR
 					(reg_q1250 AND symb_decoder(16#39#)) OR
 					(reg_q1250 AND symb_decoder(16#38#)) OR
 					(reg_q1250 AND symb_decoder(16#33#)) OR
 					(reg_q1250 AND symb_decoder(16#30#)) OR
 					(reg_q1252 AND symb_decoder(16#37#)) OR
 					(reg_q1252 AND symb_decoder(16#39#)) OR
 					(reg_q1252 AND symb_decoder(16#33#)) OR
 					(reg_q1252 AND symb_decoder(16#36#)) OR
 					(reg_q1252 AND symb_decoder(16#38#)) OR
 					(reg_q1252 AND symb_decoder(16#32#)) OR
 					(reg_q1252 AND symb_decoder(16#35#)) OR
 					(reg_q1252 AND symb_decoder(16#31#)) OR
 					(reg_q1252 AND symb_decoder(16#30#)) OR
 					(reg_q1252 AND symb_decoder(16#34#));
reg_q2620_in <= (reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2619 AND symb_decoder(16#c0#));
reg_q2622_in <= (reg_q2620 AND symb_decoder(16#53#)) OR
 					(reg_q2620 AND symb_decoder(16#73#));
reg_q2042_in <= (reg_q2040 AND symb_decoder(16#46#)) OR
 					(reg_q2040 AND symb_decoder(16#66#));
reg_q1421_in <= (reg_q1419 AND symb_decoder(16#70#)) OR
 					(reg_q1419 AND symb_decoder(16#50#));
reg_q1423_in <= (reg_q1421 AND symb_decoder(16#65#)) OR
 					(reg_q1421 AND symb_decoder(16#45#));
reg_q1680_in <= (reg_q1678 AND symb_decoder(16#52#)) OR
 					(reg_q1678 AND symb_decoder(16#72#));
reg_q1682_in <= (reg_q1680 AND symb_decoder(16#65#)) OR
 					(reg_q1680 AND symb_decoder(16#45#));
reg_q74_in <= (reg_q72 AND symb_decoder(16#53#)) OR
 					(reg_q72 AND symb_decoder(16#73#));
reg_q76_in <= (reg_q74 AND symb_decoder(16#45#)) OR
 					(reg_q74 AND symb_decoder(16#65#));
reg_q113_in <= (reg_q111 AND symb_decoder(16#50#)) OR
 					(reg_q111 AND symb_decoder(16#70#));
reg_q1187_in <= (reg_q1185 AND symb_decoder(16#41#)) OR
 					(reg_q1185 AND symb_decoder(16#61#));
reg_q1189_in <= (reg_q1187 AND symb_decoder(16#62#)) OR
 					(reg_q1187 AND symb_decoder(16#42#));
reg_q1714_in <= (reg_q1712 AND symb_decoder(16#72#)) OR
 					(reg_q1712 AND symb_decoder(16#52#));
reg_q1716_in <= (reg_q1714 AND symb_decoder(16#54#)) OR
 					(reg_q1714 AND symb_decoder(16#74#));
reg_q341_in <= (reg_q339 AND symb_decoder(16#74#)) OR
 					(reg_q339 AND symb_decoder(16#54#));
reg_q343_in <= (reg_q341 AND symb_decoder(16#72#)) OR
 					(reg_q341 AND symb_decoder(16#52#));
reg_q2117_in <= (reg_q2115 AND symb_decoder(16#4e#)) OR
 					(reg_q2115 AND symb_decoder(16#6e#));
reg_q2119_in <= (reg_q2117 AND symb_decoder(16#45#)) OR
 					(reg_q2117 AND symb_decoder(16#65#));
reg_q1574_in <= (reg_q1574 AND symb_decoder(16#20#)) OR
 					(reg_q1574 AND symb_decoder(16#0d#)) OR
 					(reg_q1574 AND symb_decoder(16#0c#)) OR
 					(reg_q1574 AND symb_decoder(16#0a#)) OR
 					(reg_q1574 AND symb_decoder(16#09#)) OR
 					(reg_q1572 AND symb_decoder(16#0c#)) OR
 					(reg_q1572 AND symb_decoder(16#09#)) OR
 					(reg_q1572 AND symb_decoder(16#0a#)) OR
 					(reg_q1572 AND symb_decoder(16#20#)) OR
 					(reg_q1572 AND symb_decoder(16#0d#));
reg_q1576_in <= (reg_q1574 AND symb_decoder(16#30#)) OR
 					(reg_q1574 AND symb_decoder(16#32#)) OR
 					(reg_q1574 AND symb_decoder(16#39#)) OR
 					(reg_q1574 AND symb_decoder(16#33#)) OR
 					(reg_q1574 AND symb_decoder(16#31#)) OR
 					(reg_q1574 AND symb_decoder(16#37#)) OR
 					(reg_q1574 AND symb_decoder(16#34#)) OR
 					(reg_q1574 AND symb_decoder(16#36#)) OR
 					(reg_q1574 AND symb_decoder(16#35#)) OR
 					(reg_q1574 AND symb_decoder(16#38#)) OR
 					(reg_q1576 AND symb_decoder(16#35#)) OR
 					(reg_q1576 AND symb_decoder(16#38#)) OR
 					(reg_q1576 AND symb_decoder(16#31#)) OR
 					(reg_q1576 AND symb_decoder(16#37#)) OR
 					(reg_q1576 AND symb_decoder(16#39#)) OR
 					(reg_q1576 AND symb_decoder(16#30#)) OR
 					(reg_q1576 AND symb_decoder(16#36#)) OR
 					(reg_q1576 AND symb_decoder(16#33#)) OR
 					(reg_q1576 AND symb_decoder(16#34#)) OR
 					(reg_q1576 AND symb_decoder(16#32#));
reg_q2215_in <= (reg_q2213 AND symb_decoder(16#49#)) OR
 					(reg_q2213 AND symb_decoder(16#69#));
reg_q2217_in <= (reg_q2215 AND symb_decoder(16#6e#)) OR
 					(reg_q2215 AND symb_decoder(16#4e#));
reg_q2609_in <= (reg_q2607 AND symb_decoder(16#52#)) OR
 					(reg_q2607 AND symb_decoder(16#72#));
reg_q2611_in <= (reg_q2609 AND symb_decoder(16#3a#));
reg_q2168_in <= (reg_q2166 AND symb_decoder(16#4d#)) OR
 					(reg_q2166 AND symb_decoder(16#6d#));
reg_q2170_in <= (reg_q2168 AND symb_decoder(16#6f#)) OR
 					(reg_q2168 AND symb_decoder(16#4f#));
reg_q994_in <= (reg_q992 AND symb_decoder(16#4c#)) OR
 					(reg_q992 AND symb_decoder(16#6c#));
reg_q996_in <= (reg_q994 AND symb_decoder(16#46#)) OR
 					(reg_q994 AND symb_decoder(16#66#));
reg_q237_in <= (reg_q237 AND symb_decoder(16#39#)) OR
 					(reg_q237 AND symb_decoder(16#34#)) OR
 					(reg_q237 AND symb_decoder(16#36#)) OR
 					(reg_q237 AND symb_decoder(16#30#)) OR
 					(reg_q237 AND symb_decoder(16#33#)) OR
 					(reg_q237 AND symb_decoder(16#31#)) OR
 					(reg_q237 AND symb_decoder(16#37#)) OR
 					(reg_q237 AND symb_decoder(16#38#)) OR
 					(reg_q237 AND symb_decoder(16#32#)) OR
 					(reg_q237 AND symb_decoder(16#35#)) OR
 					(reg_q235 AND symb_decoder(16#34#)) OR
 					(reg_q235 AND symb_decoder(16#36#)) OR
 					(reg_q235 AND symb_decoder(16#38#)) OR
 					(reg_q235 AND symb_decoder(16#30#)) OR
 					(reg_q235 AND symb_decoder(16#32#)) OR
 					(reg_q235 AND symb_decoder(16#33#)) OR
 					(reg_q235 AND symb_decoder(16#37#)) OR
 					(reg_q235 AND symb_decoder(16#39#)) OR
 					(reg_q235 AND symb_decoder(16#35#)) OR
 					(reg_q235 AND symb_decoder(16#31#));
reg_q257_in <= (reg_q257 AND symb_decoder(16#35#)) OR
 					(reg_q257 AND symb_decoder(16#33#)) OR
 					(reg_q257 AND symb_decoder(16#39#)) OR
 					(reg_q257 AND symb_decoder(16#36#)) OR
 					(reg_q257 AND symb_decoder(16#32#)) OR
 					(reg_q257 AND symb_decoder(16#37#)) OR
 					(reg_q257 AND symb_decoder(16#38#)) OR
 					(reg_q257 AND symb_decoder(16#34#)) OR
 					(reg_q257 AND symb_decoder(16#30#)) OR
 					(reg_q257 AND symb_decoder(16#31#)) OR
 					(reg_q255 AND symb_decoder(16#37#)) OR
 					(reg_q255 AND symb_decoder(16#39#)) OR
 					(reg_q255 AND symb_decoder(16#36#)) OR
 					(reg_q255 AND symb_decoder(16#34#)) OR
 					(reg_q255 AND symb_decoder(16#31#)) OR
 					(reg_q255 AND symb_decoder(16#35#)) OR
 					(reg_q255 AND symb_decoder(16#33#)) OR
 					(reg_q255 AND symb_decoder(16#32#)) OR
 					(reg_q255 AND symb_decoder(16#30#)) OR
 					(reg_q255 AND symb_decoder(16#38#));
reg_q2535_in <= (reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2534 AND symb_decoder(16#2f#));
reg_q2537_in <= (reg_q2535 AND symb_decoder(16#6e#)) OR
 					(reg_q2535 AND symb_decoder(16#4e#));
reg_q2284_in <= (reg_q2282 AND symb_decoder(16#2e#));
reg_q2286_in <= (reg_q2284 AND symb_decoder(16#39#)) OR
 					(reg_q2284 AND symb_decoder(16#34#)) OR
 					(reg_q2284 AND symb_decoder(16#37#)) OR
 					(reg_q2284 AND symb_decoder(16#31#)) OR
 					(reg_q2284 AND symb_decoder(16#32#)) OR
 					(reg_q2284 AND symb_decoder(16#36#)) OR
 					(reg_q2284 AND symb_decoder(16#35#)) OR
 					(reg_q2284 AND symb_decoder(16#38#)) OR
 					(reg_q2284 AND symb_decoder(16#30#)) OR
 					(reg_q2284 AND symb_decoder(16#33#)) OR
 					(reg_q2286 AND symb_decoder(16#36#)) OR
 					(reg_q2286 AND symb_decoder(16#30#)) OR
 					(reg_q2286 AND symb_decoder(16#39#)) OR
 					(reg_q2286 AND symb_decoder(16#35#)) OR
 					(reg_q2286 AND symb_decoder(16#32#)) OR
 					(reg_q2286 AND symb_decoder(16#37#)) OR
 					(reg_q2286 AND symb_decoder(16#34#)) OR
 					(reg_q2286 AND symb_decoder(16#33#)) OR
 					(reg_q2286 AND symb_decoder(16#38#)) OR
 					(reg_q2286 AND symb_decoder(16#31#));
reg_q682_in <= (reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q681 AND symb_decoder(16#63#)) OR
 					(reg_q681 AND symb_decoder(16#43#));
reg_q998_in <= (reg_q996 AND symb_decoder(16#74#)) OR
 					(reg_q996 AND symb_decoder(16#54#));
reg_q1000_in <= (reg_q998 AND symb_decoder(16#70#)) OR
 					(reg_q998 AND symb_decoder(16#50#));
reg_q1698_in <= (reg_q1696 AND symb_decoder(16#41#)) OR
 					(reg_q1696 AND symb_decoder(16#61#));
reg_q1700_in <= (reg_q1698 AND symb_decoder(16#52#)) OR
 					(reg_q1698 AND symb_decoder(16#72#));
reg_q2243_in <= (reg_q2243 AND symb_decoder(16#0c#)) OR
 					(reg_q2243 AND symb_decoder(16#20#)) OR
 					(reg_q2243 AND symb_decoder(16#0a#)) OR
 					(reg_q2243 AND symb_decoder(16#0d#)) OR
 					(reg_q2243 AND symb_decoder(16#09#)) OR
 					(reg_q2241 AND symb_decoder(16#0c#)) OR
 					(reg_q2241 AND symb_decoder(16#0d#)) OR
 					(reg_q2241 AND symb_decoder(16#20#)) OR
 					(reg_q2241 AND symb_decoder(16#09#)) OR
 					(reg_q2241 AND symb_decoder(16#0a#));
reg_q2245_in <= (reg_q2243 AND symb_decoder(16#32#)) OR
 					(reg_q2243 AND symb_decoder(16#31#)) OR
 					(reg_q2243 AND symb_decoder(16#34#)) OR
 					(reg_q2243 AND symb_decoder(16#36#)) OR
 					(reg_q2243 AND symb_decoder(16#38#)) OR
 					(reg_q2243 AND symb_decoder(16#33#)) OR
 					(reg_q2243 AND symb_decoder(16#39#)) OR
 					(reg_q2243 AND symb_decoder(16#37#)) OR
 					(reg_q2243 AND symb_decoder(16#35#)) OR
 					(reg_q2243 AND symb_decoder(16#30#)) OR
 					(reg_q2245 AND symb_decoder(16#34#)) OR
 					(reg_q2245 AND symb_decoder(16#37#)) OR
 					(reg_q2245 AND symb_decoder(16#38#)) OR
 					(reg_q2245 AND symb_decoder(16#35#)) OR
 					(reg_q2245 AND symb_decoder(16#31#)) OR
 					(reg_q2245 AND symb_decoder(16#32#)) OR
 					(reg_q2245 AND symb_decoder(16#39#)) OR
 					(reg_q2245 AND symb_decoder(16#36#)) OR
 					(reg_q2245 AND symb_decoder(16#30#)) OR
 					(reg_q2245 AND symb_decoder(16#33#));
reg_q1578_in <= (reg_q1576 AND symb_decoder(16#2e#));
reg_q1145_in <= (reg_q1143 AND symb_decoder(16#2e#));
reg_q1736_in <= (reg_q1736 AND symb_decoder(16#0c#)) OR
 					(reg_q1736 AND symb_decoder(16#0d#)) OR
 					(reg_q1736 AND symb_decoder(16#09#)) OR
 					(reg_q1736 AND symb_decoder(16#20#)) OR
 					(reg_q1736 AND symb_decoder(16#0a#)) OR
 					(reg_q1734 AND symb_decoder(16#0c#)) OR
 					(reg_q1734 AND symb_decoder(16#0a#)) OR
 					(reg_q1734 AND symb_decoder(16#0d#)) OR
 					(reg_q1734 AND symb_decoder(16#20#)) OR
 					(reg_q1734 AND symb_decoder(16#09#));
reg_q1738_in <= (reg_q1736 AND symb_decoder(16#69#)) OR
 					(reg_q1736 AND symb_decoder(16#49#));
reg_q2670_in <= (reg_q2668 AND symb_decoder(16#4e#)) OR
 					(reg_q2668 AND symb_decoder(16#6e#));
reg_q2672_in <= (reg_q2670 AND symb_decoder(16#47#)) OR
 					(reg_q2670 AND symb_decoder(16#67#));
reg_q288_in <= (reg_q286 AND symb_decoder(16#57#)) OR
 					(reg_q286 AND symb_decoder(16#77#));
reg_q290_in <= (reg_q288 AND symb_decoder(16#45#)) OR
 					(reg_q288 AND symb_decoder(16#65#));
reg_q125_in <= (reg_q123 AND symb_decoder(16#2e#));
reg_q1002_in <= (reg_q1000 AND symb_decoder(16#0a#)) OR
 					(reg_q1000 AND symb_decoder(16#09#)) OR
 					(reg_q1000 AND symb_decoder(16#0c#)) OR
 					(reg_q1000 AND symb_decoder(16#0d#)) OR
 					(reg_q1000 AND symb_decoder(16#20#)) OR
 					(reg_q1002 AND symb_decoder(16#09#)) OR
 					(reg_q1002 AND symb_decoder(16#0a#)) OR
 					(reg_q1002 AND symb_decoder(16#0d#)) OR
 					(reg_q1002 AND symb_decoder(16#20#)) OR
 					(reg_q1002 AND symb_decoder(16#0c#));
reg_q980_in <= (reg_q980 AND symb_decoder(16#20#)) OR
 					(reg_q980 AND symb_decoder(16#09#)) OR
 					(reg_q980 AND symb_decoder(16#0a#)) OR
 					(reg_q980 AND symb_decoder(16#0c#)) OR
 					(reg_q980 AND symb_decoder(16#0d#)) OR
 					(reg_q978 AND symb_decoder(16#0a#)) OR
 					(reg_q978 AND symb_decoder(16#0d#)) OR
 					(reg_q978 AND symb_decoder(16#0c#)) OR
 					(reg_q978 AND symb_decoder(16#20#)) OR
 					(reg_q978 AND symb_decoder(16#09#));
reg_q1702_in <= (reg_q1700 AND symb_decoder(16#44#)) OR
 					(reg_q1700 AND symb_decoder(16#64#));
reg_q371_in <= (reg_q369 AND symb_decoder(16#09#)) OR
 					(reg_q369 AND symb_decoder(16#0c#)) OR
 					(reg_q369 AND symb_decoder(16#20#)) OR
 					(reg_q369 AND symb_decoder(16#0d#)) OR
 					(reg_q369 AND symb_decoder(16#0a#)) OR
 					(reg_q371 AND symb_decoder(16#0d#)) OR
 					(reg_q371 AND symb_decoder(16#20#)) OR
 					(reg_q371 AND symb_decoder(16#0c#)) OR
 					(reg_q371 AND symb_decoder(16#09#)) OR
 					(reg_q371 AND symb_decoder(16#0a#));
reg_q919_in <= (reg_q919 AND symb_decoder(16#0d#)) OR
 					(reg_q919 AND symb_decoder(16#09#)) OR
 					(reg_q919 AND symb_decoder(16#0c#)) OR
 					(reg_q919 AND symb_decoder(16#20#)) OR
 					(reg_q919 AND symb_decoder(16#0a#)) OR
 					(reg_q917 AND symb_decoder(16#09#)) OR
 					(reg_q917 AND symb_decoder(16#0c#)) OR
 					(reg_q917 AND symb_decoder(16#20#)) OR
 					(reg_q917 AND symb_decoder(16#0d#)) OR
 					(reg_q917 AND symb_decoder(16#0a#));
reg_q921_in <= (reg_q919 AND symb_decoder(16#53#)) OR
 					(reg_q919 AND symb_decoder(16#73#));
reg_q1582_in <= (reg_q1580 AND symb_decoder(16#0d#));
reg_q931_in <= (reg_q929 AND symb_decoder(16#72#)) OR
 					(reg_q929 AND symb_decoder(16#52#));
reg_q1315_in <= (reg_q1313 AND symb_decoder(16#4e#)) OR
 					(reg_q1313 AND symb_decoder(16#6e#));
reg_q1317_in <= (reg_q1315 AND symb_decoder(16#64#)) OR
 					(reg_q1315 AND symb_decoder(16#44#));
reg_q1102_in <= (reg_q1100 AND symb_decoder(16#72#)) OR
 					(reg_q1100 AND symb_decoder(16#52#));
reg_q2692_in <= (reg_q2690 AND symb_decoder(16#21#));
reg_q2371_in <= (reg_q2369 AND symb_decoder(16#76#)) OR
 					(reg_q2369 AND symb_decoder(16#56#));
reg_q2373_in <= (reg_q2371 AND symb_decoder(16#33#)) OR
 					(reg_q2371 AND symb_decoder(16#37#)) OR
 					(reg_q2371 AND symb_decoder(16#32#)) OR
 					(reg_q2371 AND symb_decoder(16#31#)) OR
 					(reg_q2371 AND symb_decoder(16#38#)) OR
 					(reg_q2371 AND symb_decoder(16#35#)) OR
 					(reg_q2371 AND symb_decoder(16#30#)) OR
 					(reg_q2371 AND symb_decoder(16#39#)) OR
 					(reg_q2371 AND symb_decoder(16#36#)) OR
 					(reg_q2371 AND symb_decoder(16#34#)) OR
 					(reg_q2373 AND symb_decoder(16#36#)) OR
 					(reg_q2373 AND symb_decoder(16#34#)) OR
 					(reg_q2373 AND symb_decoder(16#30#)) OR
 					(reg_q2373 AND symb_decoder(16#31#)) OR
 					(reg_q2373 AND symb_decoder(16#38#)) OR
 					(reg_q2373 AND symb_decoder(16#32#)) OR
 					(reg_q2373 AND symb_decoder(16#39#)) OR
 					(reg_q2373 AND symb_decoder(16#37#)) OR
 					(reg_q2373 AND symb_decoder(16#35#)) OR
 					(reg_q2373 AND symb_decoder(16#33#));
reg_q2589_in <= (reg_q2587 AND symb_decoder(16#55#)) OR
 					(reg_q2587 AND symb_decoder(16#75#));
reg_q2591_in <= (reg_q2589 AND symb_decoder(16#72#)) OR
 					(reg_q2589 AND symb_decoder(16#52#));
reg_q2030_in <= (reg_q2030 AND symb_decoder(16#0d#)) OR
 					(reg_q2030 AND symb_decoder(16#0a#)) OR
 					(reg_q2030 AND symb_decoder(16#20#)) OR
 					(reg_q2030 AND symb_decoder(16#09#)) OR
 					(reg_q2030 AND symb_decoder(16#0c#)) OR
 					(reg_q2028 AND symb_decoder(16#0c#)) OR
 					(reg_q2028 AND symb_decoder(16#0d#)) OR
 					(reg_q2028 AND symb_decoder(16#20#)) OR
 					(reg_q2028 AND symb_decoder(16#0a#)) OR
 					(reg_q2028 AND symb_decoder(16#09#));
reg_q1339_in <= (reg_q1337 AND symb_decoder(16#32#)) OR
 					(reg_q1337 AND symb_decoder(16#35#)) OR
 					(reg_q1337 AND symb_decoder(16#36#)) OR
 					(reg_q1337 AND symb_decoder(16#31#)) OR
 					(reg_q1337 AND symb_decoder(16#39#)) OR
 					(reg_q1337 AND symb_decoder(16#30#)) OR
 					(reg_q1337 AND symb_decoder(16#33#)) OR
 					(reg_q1337 AND symb_decoder(16#37#)) OR
 					(reg_q1337 AND symb_decoder(16#34#)) OR
 					(reg_q1337 AND symb_decoder(16#38#)) OR
 					(reg_q1339 AND symb_decoder(16#33#)) OR
 					(reg_q1339 AND symb_decoder(16#34#)) OR
 					(reg_q1339 AND symb_decoder(16#37#)) OR
 					(reg_q1339 AND symb_decoder(16#30#)) OR
 					(reg_q1339 AND symb_decoder(16#31#)) OR
 					(reg_q1339 AND symb_decoder(16#35#)) OR
 					(reg_q1339 AND symb_decoder(16#32#)) OR
 					(reg_q1339 AND symb_decoder(16#39#)) OR
 					(reg_q1339 AND symb_decoder(16#38#)) OR
 					(reg_q1339 AND symb_decoder(16#36#));
reg_q1341_in <= (reg_q1339 AND symb_decoder(16#0a#)) OR
 					(reg_q1339 AND symb_decoder(16#0d#)) OR
 					(reg_q1339 AND symb_decoder(16#20#)) OR
 					(reg_q1339 AND symb_decoder(16#09#)) OR
 					(reg_q1339 AND symb_decoder(16#0c#)) OR
 					(reg_q1341 AND symb_decoder(16#0c#)) OR
 					(reg_q1341 AND symb_decoder(16#09#)) OR
 					(reg_q1341 AND symb_decoder(16#20#)) OR
 					(reg_q1341 AND symb_decoder(16#0d#)) OR
 					(reg_q1341 AND symb_decoder(16#0a#));
reg_q167_in <= (reg_q165 AND symb_decoder(16#75#)) OR
 					(reg_q165 AND symb_decoder(16#55#));
reg_q169_in <= (reg_q167 AND symb_decoder(16#4c#)) OR
 					(reg_q167 AND symb_decoder(16#6c#));
reg_q450_in <= (reg_q450 AND symb_decoder(16#32#)) OR
 					(reg_q450 AND symb_decoder(16#33#)) OR
 					(reg_q450 AND symb_decoder(16#30#)) OR
 					(reg_q450 AND symb_decoder(16#36#)) OR
 					(reg_q450 AND symb_decoder(16#39#)) OR
 					(reg_q450 AND symb_decoder(16#35#)) OR
 					(reg_q450 AND symb_decoder(16#31#)) OR
 					(reg_q450 AND symb_decoder(16#38#)) OR
 					(reg_q450 AND symb_decoder(16#37#)) OR
 					(reg_q450 AND symb_decoder(16#34#)) OR
 					(reg_q448 AND symb_decoder(16#30#)) OR
 					(reg_q448 AND symb_decoder(16#31#)) OR
 					(reg_q448 AND symb_decoder(16#33#)) OR
 					(reg_q448 AND symb_decoder(16#38#)) OR
 					(reg_q448 AND symb_decoder(16#35#)) OR
 					(reg_q448 AND symb_decoder(16#34#)) OR
 					(reg_q448 AND symb_decoder(16#36#)) OR
 					(reg_q448 AND symb_decoder(16#37#)) OR
 					(reg_q448 AND symb_decoder(16#39#)) OR
 					(reg_q448 AND symb_decoder(16#32#));
reg_q2221_in <= (reg_q2219 AND symb_decoder(16#52#)) OR
 					(reg_q2219 AND symb_decoder(16#72#));
reg_q2223_in <= (reg_q2221 AND symb_decoder(16#41#)) OR
 					(reg_q2221 AND symb_decoder(16#61#));
reg_q2634_in <= (reg_q2632 AND symb_decoder(16#c0#));
reg_q2636_in <= (reg_q2634 AND symb_decoder(16#73#)) OR
 					(reg_q2634 AND symb_decoder(16#53#));
reg_q2272_in <= (reg_q2270 AND symb_decoder(16#70#)) OR
 					(reg_q2270 AND symb_decoder(16#50#));
reg_q2115_in <= (reg_q2113 AND symb_decoder(16#41#)) OR
 					(reg_q2113 AND symb_decoder(16#61#));
reg_q333_in <= (reg_q331 AND symb_decoder(16#54#)) OR
 					(reg_q331 AND symb_decoder(16#74#));
reg_q335_in <= (reg_q333 AND symb_decoder(16#63#)) OR
 					(reg_q333 AND symb_decoder(16#43#));
reg_q1460_in <= (reg_q1458 AND symb_decoder(16#54#)) OR
 					(reg_q1458 AND symb_decoder(16#74#));
reg_q1462_in <= (reg_q1460 AND symb_decoder(16#0a#)) OR
 					(reg_q1460 AND symb_decoder(16#09#)) OR
 					(reg_q1460 AND symb_decoder(16#0d#)) OR
 					(reg_q1460 AND symb_decoder(16#20#)) OR
 					(reg_q1460 AND symb_decoder(16#0c#)) OR
 					(reg_q1462 AND symb_decoder(16#0c#)) OR
 					(reg_q1462 AND symb_decoder(16#09#)) OR
 					(reg_q1462 AND symb_decoder(16#0d#)) OR
 					(reg_q1462 AND symb_decoder(16#20#)) OR
 					(reg_q1462 AND symb_decoder(16#0a#));
reg_q2333_in <= (reg_q2331 AND symb_decoder(16#4c#)) OR
 					(reg_q2331 AND symb_decoder(16#6c#));
reg_q2335_in <= (reg_q2333 AND symb_decoder(16#46#)) OR
 					(reg_q2333 AND symb_decoder(16#66#));
reg_q2227_in <= (reg_q2225 AND symb_decoder(16#68#)) OR
 					(reg_q2225 AND symb_decoder(16#48#));
reg_q2229_in <= (reg_q2227 AND symb_decoder(16#09#)) OR
 					(reg_q2227 AND symb_decoder(16#0a#)) OR
 					(reg_q2227 AND symb_decoder(16#0c#)) OR
 					(reg_q2227 AND symb_decoder(16#0d#)) OR
 					(reg_q2227 AND symb_decoder(16#20#)) OR
 					(reg_q2229 AND symb_decoder(16#0c#)) OR
 					(reg_q2229 AND symb_decoder(16#0a#)) OR
 					(reg_q2229 AND symb_decoder(16#09#)) OR
 					(reg_q2229 AND symb_decoder(16#20#)) OR
 					(reg_q2229 AND symb_decoder(16#0d#));
reg_q1466_in <= (reg_q1464 AND symb_decoder(16#72#)) OR
 					(reg_q1464 AND symb_decoder(16#52#));
reg_q1468_in <= (reg_q1466 AND symb_decoder(16#45#)) OR
 					(reg_q1466 AND symb_decoder(16#65#));
reg_q1072_in <= (reg_q1070 AND symb_decoder(16#53#)) OR
 					(reg_q1070 AND symb_decoder(16#73#));
reg_q1074_in <= (reg_q1072 AND symb_decoder(16#65#)) OR
 					(reg_q1072 AND symb_decoder(16#45#));
reg_q2474_in <= (reg_q2472 AND symb_decoder(16#52#));
reg_q2476_in <= (reg_q2474 AND symb_decoder(16#54#));
reg_q1560_in <= (reg_q1558 AND symb_decoder(16#76#)) OR
 					(reg_q1558 AND symb_decoder(16#56#));
reg_q1562_in <= (reg_q1560 AND symb_decoder(16#65#)) OR
 					(reg_q1560 AND symb_decoder(16#45#));
reg_q686_in <= (reg_q684 AND symb_decoder(16#20#)) OR
 					(reg_q684 AND symb_decoder(16#0c#)) OR
 					(reg_q684 AND symb_decoder(16#0a#)) OR
 					(reg_q684 AND symb_decoder(16#0d#)) OR
 					(reg_q684 AND symb_decoder(16#09#));
reg_q688_in <= (reg_q686 AND symb_decoder(16#35#)) OR
 					(reg_q686 AND symb_decoder(16#39#)) OR
 					(reg_q686 AND symb_decoder(16#36#)) OR
 					(reg_q686 AND symb_decoder(16#34#)) OR
 					(reg_q686 AND symb_decoder(16#30#)) OR
 					(reg_q686 AND symb_decoder(16#31#)) OR
 					(reg_q686 AND symb_decoder(16#33#)) OR
 					(reg_q686 AND symb_decoder(16#37#)) OR
 					(reg_q686 AND symb_decoder(16#38#)) OR
 					(reg_q686 AND symb_decoder(16#32#)) OR
 					(reg_q688 AND symb_decoder(16#37#)) OR
 					(reg_q688 AND symb_decoder(16#38#)) OR
 					(reg_q688 AND symb_decoder(16#33#)) OR
 					(reg_q688 AND symb_decoder(16#36#)) OR
 					(reg_q688 AND symb_decoder(16#35#)) OR
 					(reg_q688 AND symb_decoder(16#34#)) OR
 					(reg_q688 AND symb_decoder(16#31#)) OR
 					(reg_q688 AND symb_decoder(16#30#)) OR
 					(reg_q688 AND symb_decoder(16#32#)) OR
 					(reg_q688 AND symb_decoder(16#39#));
reg_q1734_in <= (reg_q1732 AND symb_decoder(16#70#)) OR
 					(reg_q1732 AND symb_decoder(16#50#));
reg_q1704_in <= (reg_q1702 AND symb_decoder(16#65#)) OR
 					(reg_q1702 AND symb_decoder(16#45#));
reg_q305_in <= (reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q304 AND symb_decoder(16#41#)) OR
 					(reg_q304 AND symb_decoder(16#61#));
reg_q2028_in <= (reg_q2026 AND symb_decoder(16#47#)) OR
 					(reg_q2026 AND symb_decoder(16#67#));
reg_q235_in <= (reg_q233 AND symb_decoder(16#ff#));
reg_q1143_in <= (reg_q1143 AND symb_decoder(16#34#)) OR
 					(reg_q1143 AND symb_decoder(16#35#)) OR
 					(reg_q1143 AND symb_decoder(16#33#)) OR
 					(reg_q1143 AND symb_decoder(16#38#)) OR
 					(reg_q1143 AND symb_decoder(16#32#)) OR
 					(reg_q1143 AND symb_decoder(16#36#)) OR
 					(reg_q1143 AND symb_decoder(16#37#)) OR
 					(reg_q1143 AND symb_decoder(16#39#)) OR
 					(reg_q1143 AND symb_decoder(16#30#)) OR
 					(reg_q1143 AND symb_decoder(16#31#)) OR
 					(reg_q1141 AND symb_decoder(16#39#)) OR
 					(reg_q1141 AND symb_decoder(16#37#)) OR
 					(reg_q1141 AND symb_decoder(16#35#)) OR
 					(reg_q1141 AND symb_decoder(16#31#)) OR
 					(reg_q1141 AND symb_decoder(16#38#)) OR
 					(reg_q1141 AND symb_decoder(16#30#)) OR
 					(reg_q1141 AND symb_decoder(16#33#)) OR
 					(reg_q1141 AND symb_decoder(16#32#)) OR
 					(reg_q1141 AND symb_decoder(16#34#)) OR
 					(reg_q1141 AND symb_decoder(16#36#));
reg_q1541_in <= (reg_q1541 AND symb_decoder(16#39#)) OR
 					(reg_q1541 AND symb_decoder(16#38#)) OR
 					(reg_q1541 AND symb_decoder(16#32#)) OR
 					(reg_q1541 AND symb_decoder(16#30#)) OR
 					(reg_q1541 AND symb_decoder(16#36#)) OR
 					(reg_q1541 AND symb_decoder(16#33#)) OR
 					(reg_q1541 AND symb_decoder(16#34#)) OR
 					(reg_q1541 AND symb_decoder(16#37#)) OR
 					(reg_q1541 AND symb_decoder(16#31#)) OR
 					(reg_q1541 AND symb_decoder(16#35#)) OR
 					(reg_q1539 AND symb_decoder(16#35#)) OR
 					(reg_q1539 AND symb_decoder(16#34#)) OR
 					(reg_q1539 AND symb_decoder(16#32#)) OR
 					(reg_q1539 AND symb_decoder(16#39#)) OR
 					(reg_q1539 AND symb_decoder(16#37#)) OR
 					(reg_q1539 AND symb_decoder(16#30#)) OR
 					(reg_q1539 AND symb_decoder(16#33#)) OR
 					(reg_q1539 AND symb_decoder(16#36#)) OR
 					(reg_q1539 AND symb_decoder(16#38#)) OR
 					(reg_q1539 AND symb_decoder(16#31#));
reg_q1546_in <= (reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q1545 AND symb_decoder(16#6e#)) OR
 					(reg_q1545 AND symb_decoder(16#4e#));
reg_q1548_in <= (reg_q1546 AND symb_decoder(16#45#)) OR
 					(reg_q1546 AND symb_decoder(16#65#));
reg_q2022_in <= (reg_q2020 AND symb_decoder(16#52#)) OR
 					(reg_q2020 AND symb_decoder(16#72#));
reg_q2024_in <= (reg_q2022 AND symb_decoder(16#69#)) OR
 					(reg_q2022 AND symb_decoder(16#49#));
reg_q1730_in <= (reg_q1730 AND symb_decoder(16#20#)) OR
 					(reg_q1730 AND symb_decoder(16#0a#)) OR
 					(reg_q1730 AND symb_decoder(16#09#)) OR
 					(reg_q1730 AND symb_decoder(16#0c#)) OR
 					(reg_q1730 AND symb_decoder(16#0d#)) OR
 					(reg_q1728 AND symb_decoder(16#0d#)) OR
 					(reg_q1728 AND symb_decoder(16#0c#)) OR
 					(reg_q1728 AND symb_decoder(16#09#)) OR
 					(reg_q1728 AND symb_decoder(16#0a#)) OR
 					(reg_q1728 AND symb_decoder(16#20#));
reg_q1732_in <= (reg_q1730 AND symb_decoder(16#69#)) OR
 					(reg_q1730 AND symb_decoder(16#49#));
reg_q2225_in <= (reg_q2223 AND symb_decoder(16#53#)) OR
 					(reg_q2223 AND symb_decoder(16#73#));
reg_q1470_in <= (reg_q1468 AND symb_decoder(16#0a#)) OR
 					(reg_q1468 AND symb_decoder(16#20#)) OR
 					(reg_q1468 AND symb_decoder(16#0d#)) OR
 					(reg_q1468 AND symb_decoder(16#09#)) OR
 					(reg_q1468 AND symb_decoder(16#0c#)) OR
 					(reg_q1470 AND symb_decoder(16#0a#)) OR
 					(reg_q1470 AND symb_decoder(16#20#)) OR
 					(reg_q1470 AND symb_decoder(16#09#)) OR
 					(reg_q1470 AND symb_decoder(16#0d#)) OR
 					(reg_q1470 AND symb_decoder(16#0c#));
reg_q1472_in <= (reg_q1470 AND symb_decoder(16#72#)) OR
 					(reg_q1470 AND symb_decoder(16#52#));
reg_q111_in <= (reg_q111 AND symb_decoder(16#0a#)) OR
 					(reg_q111 AND symb_decoder(16#0c#)) OR
 					(reg_q111 AND symb_decoder(16#09#)) OR
 					(reg_q111 AND symb_decoder(16#20#)) OR
 					(reg_q111 AND symb_decoder(16#0d#)) OR
 					(reg_q109 AND symb_decoder(16#20#)) OR
 					(reg_q109 AND symb_decoder(16#09#)) OR
 					(reg_q109 AND symb_decoder(16#0c#)) OR
 					(reg_q109 AND symb_decoder(16#0a#)) OR
 					(reg_q109 AND symb_decoder(16#0d#));
reg_q133_in <= (reg_q131 AND symb_decoder(16#6f#)) OR
 					(reg_q131 AND symb_decoder(16#4f#));
reg_q135_in <= (reg_q133 AND symb_decoder(16#6e#)) OR
 					(reg_q133 AND symb_decoder(16#4e#));
reg_q2292_in <= (reg_q2290 AND symb_decoder(16#45#)) OR
 					(reg_q2290 AND symb_decoder(16#65#));
reg_q2294_in <= (reg_q2292 AND symb_decoder(16#72#)) OR
 					(reg_q2292 AND symb_decoder(16#52#));
reg_q1080_in <= (reg_q1078 AND symb_decoder(16#45#)) OR
 					(reg_q1078 AND symb_decoder(16#65#));
reg_q1082_in <= (reg_q1080 AND symb_decoder(16#52#)) OR
 					(reg_q1080 AND symb_decoder(16#72#));
reg_q2247_in <= (reg_q2245 AND symb_decoder(16#2e#));
reg_q2249_in <= (reg_q2247 AND symb_decoder(16#35#)) OR
 					(reg_q2247 AND symb_decoder(16#32#)) OR
 					(reg_q2247 AND symb_decoder(16#37#)) OR
 					(reg_q2247 AND symb_decoder(16#31#)) OR
 					(reg_q2247 AND symb_decoder(16#36#)) OR
 					(reg_q2247 AND symb_decoder(16#39#)) OR
 					(reg_q2247 AND symb_decoder(16#30#)) OR
 					(reg_q2247 AND symb_decoder(16#38#)) OR
 					(reg_q2247 AND symb_decoder(16#33#)) OR
 					(reg_q2247 AND symb_decoder(16#34#)) OR
 					(reg_q2249 AND symb_decoder(16#30#)) OR
 					(reg_q2249 AND symb_decoder(16#39#)) OR
 					(reg_q2249 AND symb_decoder(16#38#)) OR
 					(reg_q2249 AND symb_decoder(16#34#)) OR
 					(reg_q2249 AND symb_decoder(16#31#)) OR
 					(reg_q2249 AND symb_decoder(16#35#)) OR
 					(reg_q2249 AND symb_decoder(16#37#)) OR
 					(reg_q2249 AND symb_decoder(16#33#)) OR
 					(reg_q2249 AND symb_decoder(16#36#)) OR
 					(reg_q2249 AND symb_decoder(16#32#));
reg_q245_in <= (reg_q245 AND symb_decoder(16#37#)) OR
 					(reg_q245 AND symb_decoder(16#30#)) OR
 					(reg_q245 AND symb_decoder(16#32#)) OR
 					(reg_q245 AND symb_decoder(16#39#)) OR
 					(reg_q245 AND symb_decoder(16#36#)) OR
 					(reg_q245 AND symb_decoder(16#31#)) OR
 					(reg_q245 AND symb_decoder(16#33#)) OR
 					(reg_q245 AND symb_decoder(16#34#)) OR
 					(reg_q245 AND symb_decoder(16#38#)) OR
 					(reg_q245 AND symb_decoder(16#35#)) OR
 					(reg_q243 AND symb_decoder(16#32#)) OR
 					(reg_q243 AND symb_decoder(16#38#)) OR
 					(reg_q243 AND symb_decoder(16#30#)) OR
 					(reg_q243 AND symb_decoder(16#37#)) OR
 					(reg_q243 AND symb_decoder(16#39#)) OR
 					(reg_q243 AND symb_decoder(16#31#)) OR
 					(reg_q243 AND symb_decoder(16#34#)) OR
 					(reg_q243 AND symb_decoder(16#33#)) OR
 					(reg_q243 AND symb_decoder(16#35#)) OR
 					(reg_q243 AND symb_decoder(16#36#));
reg_q742_in <= (reg_q740 AND symb_decoder(16#74#)) OR
 					(reg_q740 AND symb_decoder(16#54#));
reg_q744_in <= (reg_q742 AND symb_decoder(16#65#)) OR
 					(reg_q742 AND symb_decoder(16#45#));
reg_q1090_in <= (reg_q1090 AND symb_decoder(16#31#)) OR
 					(reg_q1090 AND symb_decoder(16#36#)) OR
 					(reg_q1090 AND symb_decoder(16#35#)) OR
 					(reg_q1090 AND symb_decoder(16#39#)) OR
 					(reg_q1090 AND symb_decoder(16#37#)) OR
 					(reg_q1090 AND symb_decoder(16#34#)) OR
 					(reg_q1090 AND symb_decoder(16#38#)) OR
 					(reg_q1090 AND symb_decoder(16#32#)) OR
 					(reg_q1090 AND symb_decoder(16#33#)) OR
 					(reg_q1090 AND symb_decoder(16#30#)) OR
 					(reg_q1088 AND symb_decoder(16#39#)) OR
 					(reg_q1088 AND symb_decoder(16#30#)) OR
 					(reg_q1088 AND symb_decoder(16#31#)) OR
 					(reg_q1088 AND symb_decoder(16#34#)) OR
 					(reg_q1088 AND symb_decoder(16#38#)) OR
 					(reg_q1088 AND symb_decoder(16#32#)) OR
 					(reg_q1088 AND symb_decoder(16#36#)) OR
 					(reg_q1088 AND symb_decoder(16#35#)) OR
 					(reg_q1088 AND symb_decoder(16#37#)) OR
 					(reg_q1088 AND symb_decoder(16#33#));
reg_q129_in <= (reg_q127 AND symb_decoder(16#0c#)) OR
 					(reg_q127 AND symb_decoder(16#0d#)) OR
 					(reg_q127 AND symb_decoder(16#09#)) OR
 					(reg_q127 AND symb_decoder(16#0a#)) OR
 					(reg_q127 AND symb_decoder(16#20#)) OR
 					(reg_q129 AND symb_decoder(16#0a#)) OR
 					(reg_q129 AND symb_decoder(16#20#)) OR
 					(reg_q129 AND symb_decoder(16#0d#)) OR
 					(reg_q129 AND symb_decoder(16#0c#)) OR
 					(reg_q129 AND symb_decoder(16#09#));
reg_q1135_in <= (reg_q1133 AND symb_decoder(16#79#)) OR
 					(reg_q1133 AND symb_decoder(16#59#));
reg_q1137_in <= (reg_q1135 AND symb_decoder(16#0d#)) OR
 					(reg_q1135 AND symb_decoder(16#0a#)) OR
 					(reg_q1135 AND symb_decoder(16#09#)) OR
 					(reg_q1135 AND symb_decoder(16#20#)) OR
 					(reg_q1135 AND symb_decoder(16#0c#)) OR
 					(reg_q1137 AND symb_decoder(16#09#)) OR
 					(reg_q1137 AND symb_decoder(16#0c#)) OR
 					(reg_q1137 AND symb_decoder(16#0d#)) OR
 					(reg_q1137 AND symb_decoder(16#0a#)) OR
 					(reg_q1137 AND symb_decoder(16#20#));
reg_q1431_in <= (reg_q1429 AND symb_decoder(16#49#)) OR
 					(reg_q1429 AND symb_decoder(16#69#));
reg_q1433_in <= (reg_q1431 AND symb_decoder(16#4e#)) OR
 					(reg_q1431 AND symb_decoder(16#6e#));
reg_q2308_in <= (reg_q2306 AND symb_decoder(16#6c#)) OR
 					(reg_q2306 AND symb_decoder(16#4c#));
reg_q2310_in <= (reg_q2308 AND symb_decoder(16#69#)) OR
 					(reg_q2308 AND symb_decoder(16#49#));
reg_q2597_in <= (reg_q2595 AND symb_decoder(16#6e#)) OR
 					(reg_q2595 AND symb_decoder(16#4e#));
reg_q1708_in <= (reg_q1708 AND symb_decoder(16#0a#)) OR
 					(reg_q1708 AND symb_decoder(16#0d#)) OR
 					(reg_q1708 AND symb_decoder(16#0c#)) OR
 					(reg_q1708 AND symb_decoder(16#09#)) OR
 					(reg_q1708 AND symb_decoder(16#20#)) OR
 					(reg_q1706 AND symb_decoder(16#0a#)) OR
 					(reg_q1706 AND symb_decoder(16#09#)) OR
 					(reg_q1706 AND symb_decoder(16#20#)) OR
 					(reg_q1706 AND symb_decoder(16#0d#)) OR
 					(reg_q1706 AND symb_decoder(16#0c#));
reg_q2258_in <= (reg_q2256 AND symb_decoder(16#21#));
reg_q2260_in <= (reg_q2258 AND symb_decoder(16#6f#)) OR
 					(reg_q2258 AND symb_decoder(16#4f#));
reg_q978_in <= (reg_q976 AND symb_decoder(16#45#)) OR
 					(reg_q976 AND symb_decoder(16#65#));
reg_q988_in <= (reg_q986 AND symb_decoder(16#45#)) OR
 					(reg_q986 AND symb_decoder(16#65#));
reg_q990_in <= (reg_q988 AND symb_decoder(16#56#)) OR
 					(reg_q988 AND symb_decoder(16#76#));
reg_q2565_in <= (reg_q2565 AND symb_decoder(16#0a#)) OR
 					(reg_q2565 AND symb_decoder(16#0d#)) OR
 					(reg_q2565 AND symb_decoder(16#0c#)) OR
 					(reg_q2565 AND symb_decoder(16#09#)) OR
 					(reg_q2565 AND symb_decoder(16#20#)) OR
 					(reg_q2563 AND symb_decoder(16#0d#)) OR
 					(reg_q2563 AND symb_decoder(16#0c#)) OR
 					(reg_q2563 AND symb_decoder(16#20#)) OR
 					(reg_q2563 AND symb_decoder(16#0a#)) OR
 					(reg_q2563 AND symb_decoder(16#09#));
reg_q2567_in <= (reg_q2565 AND symb_decoder(16#6f#)) OR
 					(reg_q2565 AND symb_decoder(16#4f#));
reg_q1325_in <= (reg_q1323 AND symb_decoder(16#52#)) OR
 					(reg_q1323 AND symb_decoder(16#72#));
reg_q1327_in <= (reg_q1325 AND symb_decoder(16#76#)) OR
 					(reg_q1325 AND symb_decoder(16#56#));
reg_q149_in <= (reg_q149 AND symb_decoder(16#0a#)) OR
 					(reg_q149 AND symb_decoder(16#0d#)) OR
 					(reg_q149 AND symb_decoder(16#0c#)) OR
 					(reg_q149 AND symb_decoder(16#09#)) OR
 					(reg_q149 AND symb_decoder(16#20#)) OR
 					(reg_q147 AND symb_decoder(16#0d#)) OR
 					(reg_q147 AND symb_decoder(16#09#)) OR
 					(reg_q147 AND symb_decoder(16#20#)) OR
 					(reg_q147 AND symb_decoder(16#0a#)) OR
 					(reg_q147 AND symb_decoder(16#0c#));
reg_q1088_in <= (reg_q1086 AND symb_decoder(16#2e#));
reg_q137_in <= (reg_q135 AND symb_decoder(16#6e#)) OR
 					(reg_q135 AND symb_decoder(16#4e#));
reg_q675_in <= (reg_q673 AND symb_decoder(16#3a#));
reg_q2136_in <= (reg_q2134 AND symb_decoder(16#74#)) OR
 					(reg_q2134 AND symb_decoder(16#54#));
reg_q2138_in <= (reg_q2136 AND symb_decoder(16#0c#)) OR
 					(reg_q2136 AND symb_decoder(16#09#)) OR
 					(reg_q2136 AND symb_decoder(16#0a#)) OR
 					(reg_q2136 AND symb_decoder(16#0d#)) OR
 					(reg_q2136 AND symb_decoder(16#20#)) OR
 					(reg_q2138 AND symb_decoder(16#20#)) OR
 					(reg_q2138 AND symb_decoder(16#0c#)) OR
 					(reg_q2138 AND symb_decoder(16#0a#)) OR
 					(reg_q2138 AND symb_decoder(16#09#)) OR
 					(reg_q2138 AND symb_decoder(16#0d#));
reg_q119_in <= (reg_q117 AND symb_decoder(16#0a#)) OR
 					(reg_q117 AND symb_decoder(16#0d#)) OR
 					(reg_q117 AND symb_decoder(16#20#)) OR
 					(reg_q117 AND symb_decoder(16#0c#)) OR
 					(reg_q117 AND symb_decoder(16#09#)) OR
 					(reg_q119 AND symb_decoder(16#0c#)) OR
 					(reg_q119 AND symb_decoder(16#09#)) OR
 					(reg_q119 AND symb_decoder(16#0a#)) OR
 					(reg_q119 AND symb_decoder(16#20#)) OR
 					(reg_q119 AND symb_decoder(16#0d#));
reg_q255_in <= (reg_q253 AND symb_decoder(16#ff#));
reg_q915_in <= (reg_q915 AND symb_decoder(16#09#)) OR
 					(reg_q915 AND symb_decoder(16#0a#)) OR
 					(reg_q915 AND symb_decoder(16#0c#)) OR
 					(reg_q915 AND symb_decoder(16#0d#)) OR
 					(reg_q915 AND symb_decoder(16#20#)) OR
 					(reg_q913 AND symb_decoder(16#0d#)) OR
 					(reg_q913 AND symb_decoder(16#0a#)) OR
 					(reg_q913 AND symb_decoder(16#09#)) OR
 					(reg_q913 AND symb_decoder(16#20#)) OR
 					(reg_q913 AND symb_decoder(16#0c#));
reg_q1008_in <= (reg_q1006 AND symb_decoder(16#0d#));
reg_q1010_in <= (reg_q1008 AND symb_decoder(16#0a#));
reg_q1672_in <= (reg_q1670 AND symb_decoder(16#3b#));
reg_q2642_in <= (reg_q2640 AND symb_decoder(16#76#)) OR
 					(reg_q2640 AND symb_decoder(16#56#));
reg_q2644_in <= (reg_q2642 AND symb_decoder(16#65#)) OR
 					(reg_q2642 AND symb_decoder(16#45#));
reg_q2599_in <= (reg_q2597 AND symb_decoder(16#74#)) OR
 					(reg_q2597 AND symb_decoder(16#54#));
reg_q2601_in <= (reg_q2599 AND symb_decoder(16#0d#)) OR
 					(reg_q2599 AND symb_decoder(16#20#)) OR
 					(reg_q2599 AND symb_decoder(16#0a#)) OR
 					(reg_q2599 AND symb_decoder(16#0c#)) OR
 					(reg_q2599 AND symb_decoder(16#09#)) OR
 					(reg_q2601 AND symb_decoder(16#20#)) OR
 					(reg_q2601 AND symb_decoder(16#09#)) OR
 					(reg_q2601 AND symb_decoder(16#0c#)) OR
 					(reg_q2601 AND symb_decoder(16#0a#)) OR
 					(reg_q2601 AND symb_decoder(16#0d#));
reg_q1637_in <= (reg_q1635 AND symb_decoder(16#4d#)) OR
 					(reg_q1635 AND symb_decoder(16#6d#));
reg_q1639_in <= (reg_q1637 AND symb_decoder(16#0d#));
reg_q107_in <= (reg_q105 AND symb_decoder(16#49#)) OR
 					(reg_q105 AND symb_decoder(16#69#));
reg_q109_in <= (reg_q107 AND symb_decoder(16#58#)) OR
 					(reg_q107 AND symb_decoder(16#78#));
reg_q783_in <= (reg_q781 AND symb_decoder(16#6d#)) OR
 					(reg_q781 AND symb_decoder(16#4d#));
reg_q785_in <= (reg_q783 AND symb_decoder(16#69#)) OR
 					(reg_q783 AND symb_decoder(16#49#));
reg_q1092_in <= (reg_q1090 AND symb_decoder(16#09#)) OR
 					(reg_q1090 AND symb_decoder(16#0a#)) OR
 					(reg_q1090 AND symb_decoder(16#0d#)) OR
 					(reg_q1090 AND symb_decoder(16#20#)) OR
 					(reg_q1090 AND symb_decoder(16#0c#)) OR
 					(reg_q1092 AND symb_decoder(16#09#)) OR
 					(reg_q1092 AND symb_decoder(16#0c#)) OR
 					(reg_q1092 AND symb_decoder(16#0a#)) OR
 					(reg_q1092 AND symb_decoder(16#20#)) OR
 					(reg_q1092 AND symb_decoder(16#0d#));
reg_q1347_in <= (reg_q1345 AND symb_decoder(16#70#)) OR
 					(reg_q1345 AND symb_decoder(16#50#));
reg_q1349_in <= (reg_q1347 AND symb_decoder(16#6f#)) OR
 					(reg_q1347 AND symb_decoder(16#4f#));
reg_q1115_in <= (reg_q1113 AND symb_decoder(16#6f#)) OR
 					(reg_q1113 AND symb_decoder(16#4f#));
reg_q1117_in <= (reg_q1115 AND symb_decoder(16#72#)) OR
 					(reg_q1115 AND symb_decoder(16#52#));
reg_q448_in <= (reg_q448 AND symb_decoder(16#0c#)) OR
 					(reg_q448 AND symb_decoder(16#0d#)) OR
 					(reg_q448 AND symb_decoder(16#09#)) OR
 					(reg_q448 AND symb_decoder(16#0a#)) OR
 					(reg_q448 AND symb_decoder(16#20#)) OR
 					(reg_q446 AND symb_decoder(16#0c#)) OR
 					(reg_q446 AND symb_decoder(16#0d#)) OR
 					(reg_q446 AND symb_decoder(16#0a#)) OR
 					(reg_q446 AND symb_decoder(16#20#)) OR
 					(reg_q446 AND symb_decoder(16#09#));
reg_q192_in <= (reg_q190 AND symb_decoder(16#61#)) OR
 					(reg_q190 AND symb_decoder(16#41#));
reg_q395_in <= (reg_q393 AND symb_decoder(16#22#));
reg_q397_in <= (reg_q395 AND symb_decoder(16#0a#)) OR
 					(reg_q395 AND symb_decoder(16#09#)) OR
 					(reg_q395 AND symb_decoder(16#0c#)) OR
 					(reg_q395 AND symb_decoder(16#0d#)) OR
 					(reg_q395 AND symb_decoder(16#20#)) OR
 					(reg_q397 AND symb_decoder(16#0c#)) OR
 					(reg_q397 AND symb_decoder(16#20#)) OR
 					(reg_q397 AND symb_decoder(16#09#)) OR
 					(reg_q397 AND symb_decoder(16#0d#)) OR
 					(reg_q397 AND symb_decoder(16#0a#));
reg_q84_in <= (reg_q82 AND symb_decoder(16#72#)) OR
 					(reg_q82 AND symb_decoder(16#52#));
reg_q86_in <= (reg_q84 AND symb_decoder(16#0d#)) OR
 					(reg_q84 AND symb_decoder(16#0c#)) OR
 					(reg_q84 AND symb_decoder(16#09#)) OR
 					(reg_q84 AND symb_decoder(16#20#)) OR
 					(reg_q84 AND symb_decoder(16#0a#)) OR
 					(reg_q86 AND symb_decoder(16#20#)) OR
 					(reg_q86 AND symb_decoder(16#09#)) OR
 					(reg_q86 AND symb_decoder(16#0c#)) OR
 					(reg_q86 AND symb_decoder(16#0a#)) OR
 					(reg_q86 AND symb_decoder(16#0d#));
reg_q365_in <= (reg_q363 AND symb_decoder(16#31#)) OR
 					(reg_q363 AND symb_decoder(16#35#)) OR
 					(reg_q363 AND symb_decoder(16#36#)) OR
 					(reg_q363 AND symb_decoder(16#30#)) OR
 					(reg_q363 AND symb_decoder(16#38#)) OR
 					(reg_q363 AND symb_decoder(16#32#)) OR
 					(reg_q363 AND symb_decoder(16#33#)) OR
 					(reg_q363 AND symb_decoder(16#39#)) OR
 					(reg_q363 AND symb_decoder(16#34#)) OR
 					(reg_q363 AND symb_decoder(16#37#)) OR
 					(reg_q365 AND symb_decoder(16#35#)) OR
 					(reg_q365 AND symb_decoder(16#30#)) OR
 					(reg_q365 AND symb_decoder(16#36#)) OR
 					(reg_q365 AND symb_decoder(16#37#)) OR
 					(reg_q365 AND symb_decoder(16#34#)) OR
 					(reg_q365 AND symb_decoder(16#32#)) OR
 					(reg_q365 AND symb_decoder(16#33#)) OR
 					(reg_q365 AND symb_decoder(16#38#)) OR
 					(reg_q365 AND symb_decoder(16#31#)) OR
 					(reg_q365 AND symb_decoder(16#39#));
reg_q698_in <= (reg_q696 AND symb_decoder(16#2e#));
reg_q1437_in <= (reg_q1437 AND symb_decoder(16#0c#)) OR
 					(reg_q1437 AND symb_decoder(16#09#)) OR
 					(reg_q1437 AND symb_decoder(16#0a#)) OR
 					(reg_q1437 AND symb_decoder(16#0d#)) OR
 					(reg_q1437 AND symb_decoder(16#20#)) OR
 					(reg_q1435 AND symb_decoder(16#09#)) OR
 					(reg_q1435 AND symb_decoder(16#20#)) OR
 					(reg_q1435 AND symb_decoder(16#0d#)) OR
 					(reg_q1435 AND symb_decoder(16#0c#)) OR
 					(reg_q1435 AND symb_decoder(16#0a#));
reg_q964_in <= (reg_q964 AND symb_decoder(16#09#)) OR
 					(reg_q964 AND symb_decoder(16#0a#)) OR
 					(reg_q964 AND symb_decoder(16#20#)) OR
 					(reg_q964 AND symb_decoder(16#0c#)) OR
 					(reg_q964 AND symb_decoder(16#0d#)) OR
 					(reg_q962 AND symb_decoder(16#0d#)) OR
 					(reg_q962 AND symb_decoder(16#20#)) OR
 					(reg_q962 AND symb_decoder(16#0c#)) OR
 					(reg_q962 AND symb_decoder(16#0a#)) OR
 					(reg_q962 AND symb_decoder(16#09#));
reg_q748_in <= (reg_q746 AND symb_decoder(16#74#)) OR
 					(reg_q746 AND symb_decoder(16#54#));
reg_q750_in <= (reg_q748 AND symb_decoder(16#0a#)) OR
 					(reg_q748 AND symb_decoder(16#09#)) OR
 					(reg_q748 AND symb_decoder(16#0c#)) OR
 					(reg_q748 AND symb_decoder(16#0d#)) OR
 					(reg_q748 AND symb_decoder(16#20#)) OR
 					(reg_q750 AND symb_decoder(16#09#)) OR
 					(reg_q750 AND symb_decoder(16#0a#)) OR
 					(reg_q750 AND symb_decoder(16#0d#)) OR
 					(reg_q750 AND symb_decoder(16#0c#)) OR
 					(reg_q750 AND symb_decoder(16#20#));
reg_q1435_in <= (reg_q1433 AND symb_decoder(16#67#)) OR
 					(reg_q1433 AND symb_decoder(16#47#));
reg_q1692_in <= (reg_q1690 AND symb_decoder(16#0c#)) OR
 					(reg_q1690 AND symb_decoder(16#09#)) OR
 					(reg_q1690 AND symb_decoder(16#0a#)) OR
 					(reg_q1690 AND symb_decoder(16#0d#)) OR
 					(reg_q1690 AND symb_decoder(16#20#)) OR
 					(reg_q1692 AND symb_decoder(16#0d#)) OR
 					(reg_q1692 AND symb_decoder(16#0c#)) OR
 					(reg_q1692 AND symb_decoder(16#09#)) OR
 					(reg_q1692 AND symb_decoder(16#20#)) OR
 					(reg_q1692 AND symb_decoder(16#0a#));
reg_q1262_in <= (reg_q1260 AND symb_decoder(16#53#)) OR
 					(reg_q1260 AND symb_decoder(16#73#));
reg_q1264_in <= (reg_q1262 AND symb_decoder(16#45#)) OR
 					(reg_q1262 AND symb_decoder(16#65#));
reg_q2686_in <= (reg_q2684 AND symb_decoder(16#45#)) OR
 					(reg_q2684 AND symb_decoder(16#65#));
reg_q2349_in <= (reg_q2347 AND symb_decoder(16#65#)) OR
 					(reg_q2347 AND symb_decoder(16#45#));
reg_q1023_in <= (reg_q1021 AND symb_decoder(16#45#)) OR
 					(reg_q1021 AND symb_decoder(16#65#));
reg_q1025_in <= (reg_q1023 AND symb_decoder(16#72#)) OR
 					(reg_q1023 AND symb_decoder(16#52#));
reg_q1133_in <= (reg_q1131 AND symb_decoder(16#52#)) OR
 					(reg_q1131 AND symb_decoder(16#72#));
reg_q2575_in <= (reg_q2573 AND symb_decoder(16#72#)) OR
 					(reg_q2573 AND symb_decoder(16#52#));
reg_q1272_in <= (reg_q1270 AND symb_decoder(16#72#)) OR
 					(reg_q1270 AND symb_decoder(16#52#));
reg_q1274_in <= (reg_q1272 AND symb_decoder(16#0a#)) OR
 					(reg_q1272 AND symb_decoder(16#0d#)) OR
 					(reg_q1272 AND symb_decoder(16#20#)) OR
 					(reg_q1272 AND symb_decoder(16#09#)) OR
 					(reg_q1272 AND symb_decoder(16#0c#)) OR
 					(reg_q1274 AND symb_decoder(16#0c#)) OR
 					(reg_q1274 AND symb_decoder(16#0a#)) OR
 					(reg_q1274 AND symb_decoder(16#09#)) OR
 					(reg_q1274 AND symb_decoder(16#0d#)) OR
 					(reg_q1274 AND symb_decoder(16#20#));
reg_q1504_in <= (reg_q1504 AND symb_decoder(16#0a#)) OR
 					(reg_q1504 AND symb_decoder(16#20#)) OR
 					(reg_q1504 AND symb_decoder(16#0c#)) OR
 					(reg_q1504 AND symb_decoder(16#09#)) OR
 					(reg_q1504 AND symb_decoder(16#0d#)) OR
 					(reg_q1502 AND symb_decoder(16#0a#)) OR
 					(reg_q1502 AND symb_decoder(16#09#)) OR
 					(reg_q1502 AND symb_decoder(16#0c#)) OR
 					(reg_q1502 AND symb_decoder(16#0d#)) OR
 					(reg_q1502 AND symb_decoder(16#20#));
reg_q1506_in <= (reg_q1504 AND symb_decoder(16#76#)) OR
 					(reg_q1504 AND symb_decoder(16#56#));
reg_q2497_in <= (reg_q2495 AND symb_decoder(16#2a#));
reg_q2499_in <= (reg_q2497 AND symb_decoder(16#38#)) OR
 					(reg_q2497 AND symb_decoder(16#30#)) OR
 					(reg_q2497 AND symb_decoder(16#31#)) OR
 					(reg_q2497 AND symb_decoder(16#37#)) OR
 					(reg_q2497 AND symb_decoder(16#34#)) OR
 					(reg_q2497 AND symb_decoder(16#32#)) OR
 					(reg_q2497 AND symb_decoder(16#36#)) OR
 					(reg_q2497 AND symb_decoder(16#33#)) OR
 					(reg_q2497 AND symb_decoder(16#35#)) OR
 					(reg_q2497 AND symb_decoder(16#39#)) OR
 					(reg_q2499 AND symb_decoder(16#31#)) OR
 					(reg_q2499 AND symb_decoder(16#32#)) OR
 					(reg_q2499 AND symb_decoder(16#34#)) OR
 					(reg_q2499 AND symb_decoder(16#37#)) OR
 					(reg_q2499 AND symb_decoder(16#33#)) OR
 					(reg_q2499 AND symb_decoder(16#30#)) OR
 					(reg_q2499 AND symb_decoder(16#35#)) OR
 					(reg_q2499 AND symb_decoder(16#38#)) OR
 					(reg_q2499 AND symb_decoder(16#36#)) OR
 					(reg_q2499 AND symb_decoder(16#39#));
reg_q923_in <= (reg_q921 AND symb_decoder(16#65#)) OR
 					(reg_q921 AND symb_decoder(16#45#));
reg_q925_in <= (reg_q923 AND symb_decoder(16#72#)) OR
 					(reg_q923 AND symb_decoder(16#52#));
reg_q1635_in <= (reg_q1633 AND symb_decoder(16#49#)) OR
 					(reg_q1633 AND symb_decoder(16#69#));
reg_q323_in <= (reg_q321 AND symb_decoder(16#00#));
reg_q325_in <= (reg_q323 AND symb_decoder(16#00#));
reg_q292_in <= (reg_q290 AND symb_decoder(16#6c#)) OR
 					(reg_q290 AND symb_decoder(16#4c#));
reg_q294_in <= (reg_q292 AND symb_decoder(16#63#)) OR
 					(reg_q292 AND symb_decoder(16#43#));
reg_q1664_in <= (reg_q1662 AND symb_decoder(16#2e#));
reg_q1666_in <= (reg_q1664 AND symb_decoder(16#39#)) OR
 					(reg_q1664 AND symb_decoder(16#30#)) OR
 					(reg_q1664 AND symb_decoder(16#34#)) OR
 					(reg_q1664 AND symb_decoder(16#36#)) OR
 					(reg_q1664 AND symb_decoder(16#33#)) OR
 					(reg_q1664 AND symb_decoder(16#37#)) OR
 					(reg_q1664 AND symb_decoder(16#32#)) OR
 					(reg_q1664 AND symb_decoder(16#31#)) OR
 					(reg_q1664 AND symb_decoder(16#38#)) OR
 					(reg_q1664 AND symb_decoder(16#35#)) OR
 					(reg_q1666 AND symb_decoder(16#32#)) OR
 					(reg_q1666 AND symb_decoder(16#38#)) OR
 					(reg_q1666 AND symb_decoder(16#34#)) OR
 					(reg_q1666 AND symb_decoder(16#37#)) OR
 					(reg_q1666 AND symb_decoder(16#30#)) OR
 					(reg_q1666 AND symb_decoder(16#36#)) OR
 					(reg_q1666 AND symb_decoder(16#39#)) OR
 					(reg_q1666 AND symb_decoder(16#31#)) OR
 					(reg_q1666 AND symb_decoder(16#35#)) OR
 					(reg_q1666 AND symb_decoder(16#33#));
reg_q377_in <= (reg_q375 AND symb_decoder(16#48#)) OR
 					(reg_q375 AND symb_decoder(16#68#));
reg_q1652_in <= (reg_q1652 AND symb_decoder(16#0d#)) OR
 					(reg_q1652 AND symb_decoder(16#0a#)) OR
 					(reg_q1652 AND symb_decoder(16#0c#)) OR
 					(reg_q1652 AND symb_decoder(16#09#)) OR
 					(reg_q1652 AND symb_decoder(16#20#)) OR
 					(reg_q1650 AND symb_decoder(16#0c#)) OR
 					(reg_q1650 AND symb_decoder(16#0a#)) OR
 					(reg_q1650 AND symb_decoder(16#09#)) OR
 					(reg_q1650 AND symb_decoder(16#20#)) OR
 					(reg_q1650 AND symb_decoder(16#0d#));
reg_q1728_in <= (reg_q1726 AND symb_decoder(16#72#)) OR
 					(reg_q1726 AND symb_decoder(16#52#));
reg_q1151_in <= (reg_q1149 AND symb_decoder(16#0a#));
reg_q1153_in <= (reg_q1151 AND symb_decoder(16#0d#));
reg_q1971_in <= (reg_q1969 AND symb_decoder(16#45#)) OR
 					(reg_q1969 AND symb_decoder(16#65#));
reg_q1973_in <= (reg_q1971 AND symb_decoder(16#52#)) OR
 					(reg_q1971 AND symb_decoder(16#72#));
reg_q1552_in <= (reg_q1550 AND symb_decoder(16#73#)) OR
 					(reg_q1550 AND symb_decoder(16#53#));
reg_q1179_in <= (reg_q1177 AND symb_decoder(16#6e#)) OR
 					(reg_q1177 AND symb_decoder(16#4e#));
reg_q1181_in <= (reg_q1179 AND symb_decoder(16#0d#)) OR
 					(reg_q1179 AND symb_decoder(16#0c#)) OR
 					(reg_q1179 AND symb_decoder(16#0a#)) OR
 					(reg_q1179 AND symb_decoder(16#09#)) OR
 					(reg_q1179 AND symb_decoder(16#20#)) OR
 					(reg_q1181 AND symb_decoder(16#20#)) OR
 					(reg_q1181 AND symb_decoder(16#0d#)) OR
 					(reg_q1181 AND symb_decoder(16#09#)) OR
 					(reg_q1181 AND symb_decoder(16#0c#)) OR
 					(reg_q1181 AND symb_decoder(16#0a#));
reg_q913_in <= (reg_q911 AND symb_decoder(16#74#)) OR
 					(reg_q911 AND symb_decoder(16#54#));
reg_q2304_in <= (reg_q2302 AND symb_decoder(16#4f#)) OR
 					(reg_q2302 AND symb_decoder(16#6f#));
reg_q2306_in <= (reg_q2304 AND symb_decoder(16#4e#)) OR
 					(reg_q2304 AND symb_decoder(16#6e#));
reg_q1319_in <= (reg_q1317 AND symb_decoder(16#0c#)) OR
 					(reg_q1317 AND symb_decoder(16#0d#)) OR
 					(reg_q1317 AND symb_decoder(16#0a#)) OR
 					(reg_q1317 AND symb_decoder(16#20#)) OR
 					(reg_q1317 AND symb_decoder(16#09#)) OR
 					(reg_q1319 AND symb_decoder(16#0a#)) OR
 					(reg_q1319 AND symb_decoder(16#09#)) OR
 					(reg_q1319 AND symb_decoder(16#0d#)) OR
 					(reg_q1319 AND symb_decoder(16#0c#)) OR
 					(reg_q1319 AND symb_decoder(16#20#));
reg_q986_in <= (reg_q984 AND symb_decoder(16#0d#)) OR
 					(reg_q984 AND symb_decoder(16#0c#)) OR
 					(reg_q984 AND symb_decoder(16#0a#)) OR
 					(reg_q984 AND symb_decoder(16#20#)) OR
 					(reg_q984 AND symb_decoder(16#09#)) OR
 					(reg_q986 AND symb_decoder(16#20#)) OR
 					(reg_q986 AND symb_decoder(16#09#)) OR
 					(reg_q986 AND symb_decoder(16#0d#)) OR
 					(reg_q986 AND symb_decoder(16#0a#)) OR
 					(reg_q986 AND symb_decoder(16#0c#));
reg_q82_in <= (reg_q80 AND symb_decoder(16#45#)) OR
 					(reg_q80 AND symb_decoder(16#65#));
reg_q280_in <= (reg_q278 AND symb_decoder(16#61#)) OR
 					(reg_q278 AND symb_decoder(16#41#));
reg_q282_in <= (reg_q280 AND symb_decoder(16#74#)) OR
 					(reg_q280 AND symb_decoder(16#54#));
reg_q2158_in <= (reg_q2156 AND symb_decoder(16#74#)) OR
 					(reg_q2156 AND symb_decoder(16#54#));
reg_q2160_in <= (reg_q2158 AND symb_decoder(16#09#)) OR
 					(reg_q2158 AND symb_decoder(16#0d#)) OR
 					(reg_q2158 AND symb_decoder(16#0a#)) OR
 					(reg_q2158 AND symb_decoder(16#20#)) OR
 					(reg_q2158 AND symb_decoder(16#0c#)) OR
 					(reg_q2160 AND symb_decoder(16#0d#)) OR
 					(reg_q2160 AND symb_decoder(16#09#)) OR
 					(reg_q2160 AND symb_decoder(16#20#)) OR
 					(reg_q2160 AND symb_decoder(16#0a#)) OR
 					(reg_q2160 AND symb_decoder(16#0c#));
reg_q1484_in <= (reg_q1482 AND symb_decoder(16#2d#));
reg_q2674_in <= (reg_q2672 AND symb_decoder(16#20#)) OR
 					(reg_q2672 AND symb_decoder(16#09#)) OR
 					(reg_q2672 AND symb_decoder(16#0c#)) OR
 					(reg_q2672 AND symb_decoder(16#0a#)) OR
 					(reg_q2672 AND symb_decoder(16#0d#));
reg_q2676_in <= (reg_q2674 AND symb_decoder(16#53#)) OR
 					(reg_q2674 AND symb_decoder(16#73#));
reg_q440_in <= (reg_q440 AND symb_decoder(16#20#)) OR
 					(reg_q440 AND symb_decoder(16#0d#)) OR
 					(reg_q440 AND symb_decoder(16#09#)) OR
 					(reg_q440 AND symb_decoder(16#0a#)) OR
 					(reg_q440 AND symb_decoder(16#0c#)) OR
 					(reg_q438 AND symb_decoder(16#0a#)) OR
 					(reg_q438 AND symb_decoder(16#20#)) OR
 					(reg_q438 AND symb_decoder(16#0c#)) OR
 					(reg_q438 AND symb_decoder(16#0d#)) OR
 					(reg_q438 AND symb_decoder(16#09#));
reg_q442_in <= (reg_q440 AND symb_decoder(16#56#)) OR
 					(reg_q440 AND symb_decoder(16#76#));
reg_q403_in <= (reg_q401 AND symb_decoder(16#6f#)) OR
 					(reg_q401 AND symb_decoder(16#4f#));
reg_q405_in <= (reg_q403 AND symb_decoder(16#6a#)) OR
 					(reg_q403 AND symb_decoder(16#4a#));
reg_q1246_in <= (reg_q1244 AND symb_decoder(16#72#)) OR
 					(reg_q1244 AND symb_decoder(16#52#));
reg_q752_in <= (reg_q750 AND symb_decoder(16#6f#)) OR
 					(reg_q750 AND symb_decoder(16#4f#));
reg_q1445_in <= (reg_q1443 AND symb_decoder(16#54#)) OR
 					(reg_q1443 AND symb_decoder(16#74#));
reg_q2288_in <= (reg_q2286 AND symb_decoder(16#20#)) OR
 					(reg_q2286 AND symb_decoder(16#0c#)) OR
 					(reg_q2286 AND symb_decoder(16#09#)) OR
 					(reg_q2286 AND symb_decoder(16#0a#)) OR
 					(reg_q2286 AND symb_decoder(16#0d#)) OR
 					(reg_q2288 AND symb_decoder(16#20#)) OR
 					(reg_q2288 AND symb_decoder(16#0d#)) OR
 					(reg_q2288 AND symb_decoder(16#0a#)) OR
 					(reg_q2288 AND symb_decoder(16#09#)) OR
 					(reg_q2288 AND symb_decoder(16#0c#));
reg_q1490_in <= (reg_q1490 AND symb_decoder(16#0a#)) OR
 					(reg_q1490 AND symb_decoder(16#0d#)) OR
 					(reg_q1490 AND symb_decoder(16#09#)) OR
 					(reg_q1490 AND symb_decoder(16#20#)) OR
 					(reg_q1490 AND symb_decoder(16#0c#)) OR
 					(reg_q1488 AND symb_decoder(16#0c#)) OR
 					(reg_q1488 AND symb_decoder(16#0d#)) OR
 					(reg_q1488 AND symb_decoder(16#20#)) OR
 					(reg_q1488 AND symb_decoder(16#0a#)) OR
 					(reg_q1488 AND symb_decoder(16#09#));
reg_q2130_in <= (reg_q2130 AND symb_decoder(16#0d#)) OR
 					(reg_q2130 AND symb_decoder(16#0c#)) OR
 					(reg_q2130 AND symb_decoder(16#0a#)) OR
 					(reg_q2130 AND symb_decoder(16#20#)) OR
 					(reg_q2130 AND symb_decoder(16#09#)) OR
 					(reg_q2128 AND symb_decoder(16#0d#)) OR
 					(reg_q2128 AND symb_decoder(16#0a#)) OR
 					(reg_q2128 AND symb_decoder(16#0c#)) OR
 					(reg_q2128 AND symb_decoder(16#09#)) OR
 					(reg_q2128 AND symb_decoder(16#20#));
reg_q2280_in <= (reg_q2278 AND symb_decoder(16#56#)) OR
 					(reg_q2278 AND symb_decoder(16#76#));
reg_q2282_in <= (reg_q2280 AND symb_decoder(16#36#)) OR
 					(reg_q2280 AND symb_decoder(16#35#)) OR
 					(reg_q2280 AND symb_decoder(16#32#)) OR
 					(reg_q2280 AND symb_decoder(16#31#)) OR
 					(reg_q2280 AND symb_decoder(16#37#)) OR
 					(reg_q2280 AND symb_decoder(16#30#)) OR
 					(reg_q2280 AND symb_decoder(16#34#)) OR
 					(reg_q2280 AND symb_decoder(16#38#)) OR
 					(reg_q2280 AND symb_decoder(16#33#)) OR
 					(reg_q2280 AND symb_decoder(16#39#)) OR
 					(reg_q2282 AND symb_decoder(16#31#)) OR
 					(reg_q2282 AND symb_decoder(16#39#)) OR
 					(reg_q2282 AND symb_decoder(16#30#)) OR
 					(reg_q2282 AND symb_decoder(16#33#)) OR
 					(reg_q2282 AND symb_decoder(16#35#)) OR
 					(reg_q2282 AND symb_decoder(16#38#)) OR
 					(reg_q2282 AND symb_decoder(16#34#)) OR
 					(reg_q2282 AND symb_decoder(16#37#)) OR
 					(reg_q2282 AND symb_decoder(16#32#)) OR
 					(reg_q2282 AND symb_decoder(16#36#));
reg_q1535_in <= (reg_q1535 AND symb_decoder(16#09#)) OR
 					(reg_q1535 AND symb_decoder(16#20#)) OR
 					(reg_q1535 AND symb_decoder(16#0a#)) OR
 					(reg_q1535 AND symb_decoder(16#0d#)) OR
 					(reg_q1535 AND symb_decoder(16#0c#)) OR
 					(reg_q1533 AND symb_decoder(16#0a#)) OR
 					(reg_q1533 AND symb_decoder(16#20#)) OR
 					(reg_q1533 AND symb_decoder(16#0c#)) OR
 					(reg_q1533 AND symb_decoder(16#09#)) OR
 					(reg_q1533 AND symb_decoder(16#0d#));
reg_q1537_in <= (reg_q1535 AND symb_decoder(16#31#)) OR
 					(reg_q1535 AND symb_decoder(16#34#)) OR
 					(reg_q1535 AND symb_decoder(16#33#)) OR
 					(reg_q1535 AND symb_decoder(16#38#)) OR
 					(reg_q1535 AND symb_decoder(16#32#)) OR
 					(reg_q1535 AND symb_decoder(16#35#)) OR
 					(reg_q1535 AND symb_decoder(16#37#)) OR
 					(reg_q1535 AND symb_decoder(16#30#)) OR
 					(reg_q1535 AND symb_decoder(16#39#)) OR
 					(reg_q1535 AND symb_decoder(16#36#)) OR
 					(reg_q1537 AND symb_decoder(16#38#)) OR
 					(reg_q1537 AND symb_decoder(16#35#)) OR
 					(reg_q1537 AND symb_decoder(16#32#)) OR
 					(reg_q1537 AND symb_decoder(16#31#)) OR
 					(reg_q1537 AND symb_decoder(16#36#)) OR
 					(reg_q1537 AND symb_decoder(16#34#)) OR
 					(reg_q1537 AND symb_decoder(16#39#)) OR
 					(reg_q1537 AND symb_decoder(16#37#)) OR
 					(reg_q1537 AND symb_decoder(16#33#)) OR
 					(reg_q1537 AND symb_decoder(16#30#));
reg_q313_in <= (reg_q311 AND symb_decoder(16#65#)) OR
 					(reg_q311 AND symb_decoder(16#45#));
reg_q315_in <= (reg_q313 AND symb_decoder(16#52#)) OR
 					(reg_q313 AND symb_decoder(16#72#));
reg_q1556_in <= (reg_q1554 AND symb_decoder(16#59#)) OR
 					(reg_q1554 AND symb_decoder(16#79#));
reg_q1558_in <= (reg_q1556 AND symb_decoder(16#0a#)) OR
 					(reg_q1556 AND symb_decoder(16#0d#)) OR
 					(reg_q1556 AND symb_decoder(16#0c#)) OR
 					(reg_q1556 AND symb_decoder(16#20#)) OR
 					(reg_q1556 AND symb_decoder(16#09#)) OR
 					(reg_q1558 AND symb_decoder(16#0c#)) OR
 					(reg_q1558 AND symb_decoder(16#09#)) OR
 					(reg_q1558 AND symb_decoder(16#20#)) OR
 					(reg_q1558 AND symb_decoder(16#0a#)) OR
 					(reg_q1558 AND symb_decoder(16#0d#));
reg_q1439_in <= (reg_q1437 AND symb_decoder(16#73#)) OR
 					(reg_q1437 AND symb_decoder(16#53#));
reg_q2357_in <= (reg_q2355 AND symb_decoder(16#6e#)) OR
 					(reg_q2355 AND symb_decoder(16#4e#));
reg_q2359_in <= (reg_q2357 AND symb_decoder(16#41#)) OR
 					(reg_q2357 AND symb_decoder(16#61#));
reg_q2105_in <= (reg_q2103 AND symb_decoder(16#58#)) OR
 					(reg_q2103 AND symb_decoder(16#78#));
reg_q2640_in <= (reg_q2638 AND symb_decoder(16#72#)) OR
 					(reg_q2638 AND symb_decoder(16#52#));
reg_q241_in <= (reg_q241 AND symb_decoder(16#36#)) OR
 					(reg_q241 AND symb_decoder(16#37#)) OR
 					(reg_q241 AND symb_decoder(16#32#)) OR
 					(reg_q241 AND symb_decoder(16#38#)) OR
 					(reg_q241 AND symb_decoder(16#31#)) OR
 					(reg_q241 AND symb_decoder(16#39#)) OR
 					(reg_q241 AND symb_decoder(16#35#)) OR
 					(reg_q241 AND symb_decoder(16#34#)) OR
 					(reg_q241 AND symb_decoder(16#30#)) OR
 					(reg_q241 AND symb_decoder(16#33#)) OR
 					(reg_q239 AND symb_decoder(16#39#)) OR
 					(reg_q239 AND symb_decoder(16#33#)) OR
 					(reg_q239 AND symb_decoder(16#35#)) OR
 					(reg_q239 AND symb_decoder(16#34#)) OR
 					(reg_q239 AND symb_decoder(16#31#)) OR
 					(reg_q239 AND symb_decoder(16#30#)) OR
 					(reg_q239 AND symb_decoder(16#36#)) OR
 					(reg_q239 AND symb_decoder(16#32#)) OR
 					(reg_q239 AND symb_decoder(16#38#)) OR
 					(reg_q239 AND symb_decoder(16#37#));
reg_q1313_in <= (reg_q1311 AND symb_decoder(16#45#)) OR
 					(reg_q1311 AND symb_decoder(16#65#));
reg_q1256_in <= (reg_q1256 AND symb_decoder(16#38#)) OR
 					(reg_q1256 AND symb_decoder(16#31#)) OR
 					(reg_q1256 AND symb_decoder(16#32#)) OR
 					(reg_q1256 AND symb_decoder(16#37#)) OR
 					(reg_q1256 AND symb_decoder(16#33#)) OR
 					(reg_q1256 AND symb_decoder(16#34#)) OR
 					(reg_q1256 AND symb_decoder(16#39#)) OR
 					(reg_q1256 AND symb_decoder(16#30#)) OR
 					(reg_q1256 AND symb_decoder(16#36#)) OR
 					(reg_q1256 AND symb_decoder(16#35#)) OR
 					(reg_q1254 AND symb_decoder(16#36#)) OR
 					(reg_q1254 AND symb_decoder(16#33#)) OR
 					(reg_q1254 AND symb_decoder(16#39#)) OR
 					(reg_q1254 AND symb_decoder(16#32#)) OR
 					(reg_q1254 AND symb_decoder(16#31#)) OR
 					(reg_q1254 AND symb_decoder(16#35#)) OR
 					(reg_q1254 AND symb_decoder(16#37#)) OR
 					(reg_q1254 AND symb_decoder(16#38#)) OR
 					(reg_q1254 AND symb_decoder(16#30#)) OR
 					(reg_q1254 AND symb_decoder(16#34#));
reg_q1033_in <= (reg_q1031 AND symb_decoder(16#6e#)) OR
 					(reg_q1031 AND symb_decoder(16#4e#));
reg_q2624_in <= (reg_q2622 AND symb_decoder(16#74#)) OR
 					(reg_q2622 AND symb_decoder(16#54#));
reg_q974_in <= (reg_q972 AND symb_decoder(16#6f#)) OR
 					(reg_q972 AND symb_decoder(16#4f#));
reg_q976_in <= (reg_q974 AND symb_decoder(16#6d#)) OR
 					(reg_q974 AND symb_decoder(16#4d#));
reg_q992_in <= (reg_q990 AND symb_decoder(16#69#)) OR
 					(reg_q990 AND symb_decoder(16#49#));
reg_q298_in <= (reg_q296 AND symb_decoder(16#4d#)) OR
 					(reg_q296 AND symb_decoder(16#6d#));
reg_q300_in <= (reg_q298 AND symb_decoder(16#45#)) OR
 					(reg_q298 AND symb_decoder(16#65#));
reg_q696_in <= (reg_q696 AND symb_decoder(16#39#)) OR
 					(reg_q696 AND symb_decoder(16#34#)) OR
 					(reg_q696 AND symb_decoder(16#38#)) OR
 					(reg_q696 AND symb_decoder(16#30#)) OR
 					(reg_q696 AND symb_decoder(16#31#)) OR
 					(reg_q696 AND symb_decoder(16#35#)) OR
 					(reg_q696 AND symb_decoder(16#36#)) OR
 					(reg_q696 AND symb_decoder(16#37#)) OR
 					(reg_q696 AND symb_decoder(16#32#)) OR
 					(reg_q696 AND symb_decoder(16#33#)) OR
 					(reg_q694 AND symb_decoder(16#37#)) OR
 					(reg_q694 AND symb_decoder(16#39#)) OR
 					(reg_q694 AND symb_decoder(16#35#)) OR
 					(reg_q694 AND symb_decoder(16#36#)) OR
 					(reg_q694 AND symb_decoder(16#33#)) OR
 					(reg_q694 AND symb_decoder(16#30#)) OR
 					(reg_q694 AND symb_decoder(16#38#)) OR
 					(reg_q694 AND symb_decoder(16#32#)) OR
 					(reg_q694 AND symb_decoder(16#34#)) OR
 					(reg_q694 AND symb_decoder(16#31#));
reg_q1539_in <= (reg_q1537 AND symb_decoder(16#2e#));
reg_q161_in <= (reg_q159 AND symb_decoder(16#53#)) OR
 					(reg_q159 AND symb_decoder(16#73#));
reg_q163_in <= (reg_q161 AND symb_decoder(16#53#)) OR
 					(reg_q161 AND symb_decoder(16#73#));
reg_q2547_in <= (reg_q2545 AND symb_decoder(16#45#)) OR
 					(reg_q2545 AND symb_decoder(16#65#));
reg_q2549_in <= (reg_q2547 AND symb_decoder(16#47#)) OR
 					(reg_q2547 AND symb_decoder(16#67#));
reg_q1070_in <= (reg_q1070 AND symb_decoder(16#20#)) OR
 					(reg_q1070 AND symb_decoder(16#0a#)) OR
 					(reg_q1070 AND symb_decoder(16#0c#)) OR
 					(reg_q1070 AND symb_decoder(16#0d#)) OR
 					(reg_q1070 AND symb_decoder(16#09#)) OR
 					(reg_q1068 AND symb_decoder(16#0d#)) OR
 					(reg_q1068 AND symb_decoder(16#09#)) OR
 					(reg_q1068 AND symb_decoder(16#0c#)) OR
 					(reg_q1068 AND symb_decoder(16#20#)) OR
 					(reg_q1068 AND symb_decoder(16#0a#));
reg_q438_in <= (reg_q436 AND symb_decoder(16#52#)) OR
 					(reg_q436 AND symb_decoder(16#72#));
reg_q1710_in <= (reg_q1708 AND symb_decoder(16#50#)) OR
 					(reg_q1708 AND symb_decoder(16#70#));
reg_q1712_in <= (reg_q1710 AND symb_decoder(16#4f#)) OR
 					(reg_q1710 AND symb_decoder(16#6f#));
reg_q407_in <= (reg_q405 AND symb_decoder(16#45#)) OR
 					(reg_q405 AND symb_decoder(16#65#));
reg_q409_in <= (reg_q407 AND symb_decoder(16#43#)) OR
 					(reg_q407 AND symb_decoder(16#63#));
reg_q2470_in <= (reg_q2468 AND symb_decoder(16#50#));
reg_q2472_in <= (reg_q2470 AND symb_decoder(16#4f#));
reg_q200_in <= (reg_q198 AND symb_decoder(16#54#)) OR
 					(reg_q198 AND symb_decoder(16#74#));
reg_q88_in <= (reg_q86 AND symb_decoder(16#3f#));
reg_q1230_in <= (reg_q1228 AND symb_decoder(16#54#)) OR
 					(reg_q1228 AND symb_decoder(16#74#));
reg_q1232_in <= (reg_q1230 AND symb_decoder(16#65#)) OR
 					(reg_q1230 AND symb_decoder(16#45#));
reg_q2646_in <= (reg_q2644 AND symb_decoder(16#72#)) OR
 					(reg_q2644 AND symb_decoder(16#52#));
reg_q2648_in <= (reg_q2646 AND symb_decoder(16#20#)) OR
 					(reg_q2646 AND symb_decoder(16#0a#)) OR
 					(reg_q2646 AND symb_decoder(16#0d#)) OR
 					(reg_q2646 AND symb_decoder(16#09#)) OR
 					(reg_q2646 AND symb_decoder(16#0c#));
reg_q1254_in <= (reg_q1252 AND symb_decoder(16#2e#));
reg_q1474_in <= (reg_q1472 AND symb_decoder(16#45#)) OR
 					(reg_q1472 AND symb_decoder(16#65#));
reg_q66_in <= (reg_q64 AND symb_decoder(16#74#)) OR
 					(reg_q64 AND symb_decoder(16#54#));
reg_q68_in <= (reg_q66 AND symb_decoder(16#65#)) OR
 					(reg_q66 AND symb_decoder(16#45#));
reg_q2300_in <= (reg_q2298 AND symb_decoder(16#72#)) OR
 					(reg_q2298 AND symb_decoder(16#52#));
reg_q2268_in <= (reg_q2266 AND symb_decoder(16#58#)) OR
 					(reg_q2266 AND symb_decoder(16#78#));
reg_q2270_in <= (reg_q2268 AND symb_decoder(16#09#)) OR
 					(reg_q2268 AND symb_decoder(16#0c#)) OR
 					(reg_q2268 AND symb_decoder(16#20#)) OR
 					(reg_q2268 AND symb_decoder(16#0d#)) OR
 					(reg_q2268 AND symb_decoder(16#0a#)) OR
 					(reg_q2270 AND symb_decoder(16#0c#)) OR
 					(reg_q2270 AND symb_decoder(16#0a#)) OR
 					(reg_q2270 AND symb_decoder(16#09#)) OR
 					(reg_q2270 AND symb_decoder(16#0d#)) OR
 					(reg_q2270 AND symb_decoder(16#20#));
reg_q2032_in <= (reg_q2030 AND symb_decoder(16#66#)) OR
 					(reg_q2030 AND symb_decoder(16#46#));
reg_q2034_in <= (reg_q2032 AND symb_decoder(16#49#)) OR
 					(reg_q2032 AND symb_decoder(16#69#));
reg_q430_in <= (reg_q428 AND symb_decoder(16#75#)) OR
 					(reg_q428 AND symb_decoder(16#55#));
reg_q766_in <= (reg_q764 AND symb_decoder(16#63#)) OR
 					(reg_q764 AND symb_decoder(16#43#));
reg_q768_in <= (reg_q766 AND symb_decoder(16#74#)) OR
 					(reg_q766 AND symb_decoder(16#54#));
reg_q2662_in <= (reg_q2660 AND symb_decoder(16#6f#)) OR
 					(reg_q2660 AND symb_decoder(16#4f#));
reg_q2664_in <= (reg_q2662 AND symb_decoder(16#47#)) OR
 					(reg_q2662 AND symb_decoder(16#67#));
reg_q139_in <= (reg_q137 AND symb_decoder(16#65#)) OR
 					(reg_q137 AND symb_decoder(16#45#));
reg_q1141_in <= (reg_q1139 AND symb_decoder(16#2e#));
reg_q2010_in <= (reg_q2008 AND symb_decoder(16#41#)) OR
 					(reg_q2008 AND symb_decoder(16#61#));
reg_q2012_in <= (reg_q2010 AND symb_decoder(16#4e#)) OR
 					(reg_q2010 AND symb_decoder(16#6e#));
reg_q1068_in <= (reg_q1066 AND symb_decoder(16#72#)) OR
 					(reg_q1066 AND symb_decoder(16#52#));
reg_q2557_in <= (reg_q2555 AND symb_decoder(16#65#)) OR
 					(reg_q2555 AND symb_decoder(16#45#));
reg_q2559_in <= (reg_q2557 AND symb_decoder(16#72#)) OR
 					(reg_q2557 AND symb_decoder(16#52#));
reg_q1617_in <= (reg_q1615 AND symb_decoder(16#52#)) OR
 					(reg_q1615 AND symb_decoder(16#72#));
reg_q1619_in <= (reg_q1617 AND symb_decoder(16#65#)) OR
 					(reg_q1617 AND symb_decoder(16#45#));
reg_q1258_in <= (reg_q1256 AND symb_decoder(16#2c#));
reg_q1260_in <= (reg_q1258 AND symb_decoder(16#09#)) OR
 					(reg_q1258 AND symb_decoder(16#0c#)) OR
 					(reg_q1258 AND symb_decoder(16#0d#)) OR
 					(reg_q1258 AND symb_decoder(16#0a#)) OR
 					(reg_q1258 AND symb_decoder(16#20#)) OR
 					(reg_q1260 AND symb_decoder(16#0a#)) OR
 					(reg_q1260 AND symb_decoder(16#09#)) OR
 					(reg_q1260 AND symb_decoder(16#0c#)) OR
 					(reg_q1260 AND symb_decoder(16#20#)) OR
 					(reg_q1260 AND symb_decoder(16#0d#));
reg_q734_in <= (reg_q734 AND symb_decoder(16#0d#)) OR
 					(reg_q734 AND symb_decoder(16#0a#)) OR
 					(reg_q734 AND symb_decoder(16#20#)) OR
 					(reg_q734 AND symb_decoder(16#09#)) OR
 					(reg_q734 AND symb_decoder(16#0c#)) OR
 					(reg_q732 AND symb_decoder(16#0d#)) OR
 					(reg_q732 AND symb_decoder(16#09#)) OR
 					(reg_q732 AND symb_decoder(16#20#)) OR
 					(reg_q732 AND symb_decoder(16#0c#)) OR
 					(reg_q732 AND symb_decoder(16#0a#));
reg_q1447_in <= (reg_q1445 AND symb_decoder(16#45#)) OR
 					(reg_q1445 AND symb_decoder(16#65#));
reg_q2014_in <= (reg_q2012 AND symb_decoder(16#53#)) OR
 					(reg_q2012 AND symb_decoder(16#73#));
reg_q2502_in <= (reg_q2695 AND symb_decoder(16#2a#));
reg_q2296_in <= (reg_q2294 AND symb_decoder(16#76#)) OR
 					(reg_q2294 AND symb_decoder(16#56#));
reg_q2298_in <= (reg_q2296 AND symb_decoder(16#65#)) OR
 					(reg_q2296 AND symb_decoder(16#45#));
reg_q1159_in <= (reg_q1157 AND symb_decoder(16#0a#));
reg_q444_in <= (reg_q442 AND symb_decoder(16#65#)) OR
 					(reg_q442 AND symb_decoder(16#45#));
reg_q446_in <= (reg_q444 AND symb_decoder(16#52#)) OR
 					(reg_q444 AND symb_decoder(16#72#));
reg_q1183_in <= (reg_q1181 AND symb_decoder(16#53#)) OR
 					(reg_q1181 AND symb_decoder(16#73#));
reg_q1185_in <= (reg_q1183 AND symb_decoder(16#54#)) OR
 					(reg_q1183 AND symb_decoder(16#74#));
reg_q962_in <= (reg_q960 AND symb_decoder(16#2d#));
reg_q2573_in <= (reg_q2571 AND symb_decoder(16#45#)) OR
 					(reg_q2571 AND symb_decoder(16#65#));
reg_q1123_in <= (reg_q1121 AND symb_decoder(16#44#)) OR
 					(reg_q1121 AND symb_decoder(16#64#));
reg_q1125_in <= (reg_q1123 AND symb_decoder(16#0a#)) OR
 					(reg_q1123 AND symb_decoder(16#0c#)) OR
 					(reg_q1123 AND symb_decoder(16#20#)) OR
 					(reg_q1123 AND symb_decoder(16#0d#)) OR
 					(reg_q1123 AND symb_decoder(16#09#)) OR
 					(reg_q1125 AND symb_decoder(16#0a#)) OR
 					(reg_q1125 AND symb_decoder(16#09#)) OR
 					(reg_q1125 AND symb_decoder(16#20#)) OR
 					(reg_q1125 AND symb_decoder(16#0d#)) OR
 					(reg_q1125 AND symb_decoder(16#0c#));
reg_q1613_in <= (reg_q1613 AND symb_decoder(16#09#)) OR
 					(reg_q1613 AND symb_decoder(16#20#)) OR
 					(reg_q1613 AND symb_decoder(16#0c#)) OR
 					(reg_q1613 AND symb_decoder(16#0a#)) OR
 					(reg_q1613 AND symb_decoder(16#0d#)) OR
 					(reg_q1611 AND symb_decoder(16#20#)) OR
 					(reg_q1611 AND symb_decoder(16#0d#)) OR
 					(reg_q1611 AND symb_decoder(16#09#)) OR
 					(reg_q1611 AND symb_decoder(16#0a#)) OR
 					(reg_q1611 AND symb_decoder(16#0c#));
reg_q2339_in <= (reg_q2337 AND symb_decoder(16#52#)) OR
 					(reg_q2337 AND symb_decoder(16#72#));
reg_q667_in <= (reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q666 AND symb_decoder(16#42#)) OR
 					(reg_q666 AND symb_decoder(16#62#));
reg_q60_in <= (reg_q58 AND symb_decoder(16#45#)) OR
 					(reg_q58 AND symb_decoder(16#65#));
reg_q399_in <= (reg_q397 AND symb_decoder(16#70#)) OR
 					(reg_q397 AND symb_decoder(16#50#));
reg_q2650_in <= (reg_q2648 AND symb_decoder(16#3a#));
reg_q1076_in <= (reg_q1074 AND symb_decoder(16#52#)) OR
 					(reg_q1074 AND symb_decoder(16#72#));
reg_q1078_in <= (reg_q1076 AND symb_decoder(16#56#)) OR
 					(reg_q1076 AND symb_decoder(16#76#));
reg_q284_in <= (reg_q282 AND symb_decoder(16#48#)) OR
 					(reg_q282 AND symb_decoder(16#68#));
reg_q2095_in <= (reg_q2093 AND symb_decoder(16#41#)) OR
 					(reg_q2093 AND symb_decoder(16#61#));
reg_q171_in <= (reg_q169 AND symb_decoder(16#6c#)) OR
 					(reg_q169 AND symb_decoder(16#4c#));
reg_q239_in <= (reg_q237 AND symb_decoder(16#ff#));
reg_q278_in <= (reg_q276 AND symb_decoder(16#45#)) OR
 					(reg_q276 AND symb_decoder(16#65#));
reg_q105_in <= (reg_q103 AND symb_decoder(16#74#)) OR
 					(reg_q103 AND symb_decoder(16#54#));
reg_q2148_in <= (reg_q2148 AND symb_decoder(16#0a#)) OR
 					(reg_q2148 AND symb_decoder(16#09#)) OR
 					(reg_q2148 AND symb_decoder(16#0d#)) OR
 					(reg_q2148 AND symb_decoder(16#0c#)) OR
 					(reg_q2148 AND symb_decoder(16#20#)) OR
 					(reg_q2146 AND symb_decoder(16#0a#)) OR
 					(reg_q2146 AND symb_decoder(16#0c#)) OR
 					(reg_q2146 AND symb_decoder(16#09#)) OR
 					(reg_q2146 AND symb_decoder(16#20#)) OR
 					(reg_q2146 AND symb_decoder(16#0d#));
reg_q1343_in <= (reg_q1341 AND symb_decoder(16#2e#));
reg_q1625_in <= (reg_q1623 AND symb_decoder(16#5f#));
reg_q1627_in <= (reg_q1625 AND symb_decoder(16#56#)) OR
 					(reg_q1625 AND symb_decoder(16#76#));
reg_q349_in <= (reg_q347 AND symb_decoder(16#2e#));
reg_q351_in <= (reg_q349 AND symb_decoder(16#73#)) OR
 					(reg_q349 AND symb_decoder(16#53#));
reg_q1648_in <= (reg_q1646 AND symb_decoder(16#74#)) OR
 					(reg_q1646 AND symb_decoder(16#54#));
reg_q307_in <= (reg_q305 AND symb_decoder(16#4e#)) OR
 					(reg_q305 AND symb_decoder(16#6e#));
reg_q2290_in <= (reg_q2288 AND symb_decoder(16#73#)) OR
 					(reg_q2288 AND symb_decoder(16#53#));
reg_q1533_in <= (reg_q1531 AND symb_decoder(16#53#)) OR
 					(reg_q1531 AND symb_decoder(16#73#));
reg_q2237_in <= (reg_q2235 AND symb_decoder(16#76#)) OR
 					(reg_q2235 AND symb_decoder(16#56#));
reg_q2239_in <= (reg_q2237 AND symb_decoder(16#45#)) OR
 					(reg_q2237 AND symb_decoder(16#65#));
reg_q1242_in <= (reg_q1240 AND symb_decoder(16#68#)) OR
 					(reg_q1240 AND symb_decoder(16#48#));
reg_q1244_in <= (reg_q1242 AND symb_decoder(16#45#)) OR
 					(reg_q1242 AND symb_decoder(16#65#));
reg_q1282_in <= (reg_q1280 AND symb_decoder(16#6c#)) OR
 					(reg_q1280 AND symb_decoder(16#4c#));
reg_q1284_in <= (reg_q1282 AND symb_decoder(16#49#)) OR
 					(reg_q1282 AND symb_decoder(16#69#));
reg_q1570_in <= (reg_q1568 AND symb_decoder(16#6f#)) OR
 					(reg_q1568 AND symb_decoder(16#4f#));
reg_q1572_in <= (reg_q1570 AND symb_decoder(16#4e#)) OR
 					(reg_q1570 AND symb_decoder(16#6e#));
reg_q1706_in <= (reg_q1704 AND symb_decoder(16#44#)) OR
 					(reg_q1704 AND symb_decoder(16#64#));
reg_q436_in <= (reg_q434 AND symb_decoder(16#65#)) OR
 					(reg_q434 AND symb_decoder(16#45#));
reg_q220_in <= (reg_q218 AND symb_decoder(16#69#)) OR
 					(reg_q218 AND symb_decoder(16#49#));
reg_q222_in <= (reg_q220 AND symb_decoder(16#4e#)) OR
 					(reg_q220 AND symb_decoder(16#6e#));
reg_q210_in <= (reg_q208 AND symb_decoder(16#5e#));
reg_q212_in <= (reg_q210 AND symb_decoder(16#4d#)) OR
 					(reg_q210 AND symb_decoder(16#6d#));
reg_q78_in <= (reg_q76 AND symb_decoder(16#72#)) OR
 					(reg_q76 AND symb_decoder(16#52#));
reg_q80_in <= (reg_q78 AND symb_decoder(16#56#)) OR
 					(reg_q78 AND symb_decoder(16#76#));
reg_q684_in <= (reg_q682 AND symb_decoder(16#31#));
reg_q1039_in <= (reg_q1037 AND symb_decoder(16#65#)) OR
 					(reg_q1037 AND symb_decoder(16#45#));
reg_q1041_in <= (reg_q1039 AND symb_decoder(16#72#)) OR
 					(reg_q1039 AND symb_decoder(16#52#));
reg_q2241_in <= (reg_q2239 AND symb_decoder(16#52#)) OR
 					(reg_q2239 AND symb_decoder(16#72#));
reg_q2233_in <= (reg_q2231 AND symb_decoder(16#45#)) OR
 					(reg_q2231 AND symb_decoder(16#65#));
reg_q2235_in <= (reg_q2233 AND symb_decoder(16#52#)) OR
 					(reg_q2233 AND symb_decoder(16#72#));
reg_q972_in <= (reg_q970 AND symb_decoder(16#63#)) OR
 					(reg_q970 AND symb_decoder(16#43#));
reg_q2219_in <= (reg_q2217 AND symb_decoder(16#63#)) OR
 					(reg_q2217 AND symb_decoder(16#43#));
reg_q1492_in <= (reg_q1490 AND symb_decoder(16#73#)) OR
 					(reg_q1490 AND symb_decoder(16#53#));
reg_q1554_in <= (reg_q1552 AND symb_decoder(16#70#)) OR
 					(reg_q1552 AND symb_decoder(16#50#));
reg_q2495_in <= (reg_q2493 AND symb_decoder(16#32#));
reg_q2231_in <= (reg_q2229 AND symb_decoder(16#53#)) OR
 					(reg_q2229 AND symb_decoder(16#73#));
reg_q724_in <= (reg_q722 AND symb_decoder(16#74#)) OR
 					(reg_q722 AND symb_decoder(16#54#));
reg_q726_in <= (reg_q724 AND symb_decoder(16#54#)) OR
 					(reg_q724 AND symb_decoder(16#74#));
reg_q2113_in <= (reg_q2111 AND symb_decoder(16#59#)) OR
 					(reg_q2111 AND symb_decoder(16#79#));
reg_q2144_in <= (reg_q2142 AND symb_decoder(16#69#)) OR
 					(reg_q2142 AND symb_decoder(16#49#));
reg_q2146_in <= (reg_q2144 AND symb_decoder(16#73#)) OR
 					(reg_q2144 AND symb_decoder(16#53#));
reg_q1228_in <= (reg_q1226 AND symb_decoder(16#61#)) OR
 					(reg_q1226 AND symb_decoder(16#41#));
reg_q1650_in <= (reg_q1648 AND symb_decoder(16#62#)) OR
 					(reg_q1648 AND symb_decoder(16#42#));
reg_q147_in <= (reg_q145 AND symb_decoder(16#44#)) OR
 					(reg_q145 AND symb_decoder(16#64#));
reg_q296_in <= (reg_q294 AND symb_decoder(16#6f#)) OR
 					(reg_q294 AND symb_decoder(16#4f#));
reg_q1611_in <= (reg_q1609 AND symb_decoder(16#6b#)) OR
 					(reg_q1609 AND symb_decoder(16#4b#));
reg_q1169_in <= (reg_q1167 AND symb_decoder(16#65#)) OR
 					(reg_q1167 AND symb_decoder(16#45#));
reg_q1171_in <= (reg_q1169 AND symb_decoder(16#63#)) OR
 					(reg_q1169 AND symb_decoder(16#43#));
reg_q1017_in <= (reg_q1015 AND symb_decoder(16#72#)) OR
 					(reg_q1015 AND symb_decoder(16#52#));
reg_q1019_in <= (reg_q1017 AND symb_decoder(16#41#)) OR
 					(reg_q1017 AND symb_decoder(16#61#));
reg_q2571_in <= (reg_q2569 AND symb_decoder(16#6e#)) OR
 					(reg_q2569 AND symb_decoder(16#4e#));
reg_q1615_in <= (reg_q1613 AND symb_decoder(16#66#)) OR
 					(reg_q1613 AND symb_decoder(16#46#));
reg_q2561_in <= (reg_q2559 AND symb_decoder(16#65#)) OR
 					(reg_q2559 AND symb_decoder(16#45#));
reg_q1353_in <= (reg_q1351 AND symb_decoder(16#54#)) OR
 					(reg_q1351 AND symb_decoder(16#74#));
reg_q1127_in <= (reg_q1125 AND symb_decoder(16#45#)) OR
 					(reg_q1125 AND symb_decoder(16#65#));
reg_q1129_in <= (reg_q1127 AND symb_decoder(16#4e#)) OR
 					(reg_q1127 AND symb_decoder(16#6e#));
reg_q1351_in <= (reg_q1349 AND symb_decoder(16#52#)) OR
 					(reg_q1349 AND symb_decoder(16#72#));
reg_q385_in <= (reg_q383 AND symb_decoder(16#4e#)) OR
 					(reg_q383 AND symb_decoder(16#6e#));
reg_q387_in <= (reg_q385 AND symb_decoder(16#73#)) OR
 					(reg_q385 AND symb_decoder(16#53#));
reg_q432_in <= (reg_q430 AND symb_decoder(16#6e#)) OR
 					(reg_q430 AND symb_decoder(16#4e#));
reg_q2318_in <= (reg_q2316 AND symb_decoder(16#21#));
reg_q2320_in <= (reg_q2318 AND symb_decoder(16#21#));
reg_q2682_in <= (reg_q2680 AND symb_decoder(16#72#)) OR
 					(reg_q2680 AND symb_decoder(16#52#));
reg_q2684_in <= (reg_q2682 AND symb_decoder(16#74#)) OR
 					(reg_q2682 AND symb_decoder(16#54#));
reg_q1514_in <= (reg_q1512 AND symb_decoder(16#69#)) OR
 					(reg_q1512 AND symb_decoder(16#49#));
reg_q1516_in <= (reg_q1514 AND symb_decoder(16#4f#)) OR
 					(reg_q1514 AND symb_decoder(16#6f#));
reg_q2107_in <= (reg_q2105 AND symb_decoder(16#68#)) OR
 					(reg_q2105 AND symb_decoder(16#48#));
reg_q728_in <= (reg_q726 AND symb_decoder(16#49#)) OR
 					(reg_q726 AND symb_decoder(16#69#));
reg_q2329_in <= (reg_q2327 AND symb_decoder(16#6f#)) OR
 					(reg_q2327 AND symb_decoder(16#4f#));
reg_q2331_in <= (reg_q2329 AND symb_decoder(16#4c#)) OR
 					(reg_q2329 AND symb_decoder(16#6c#));
reg_q1157_in <= (reg_q1155 AND symb_decoder(16#0d#));
reg_q2654_in <= (reg_q2652 AND symb_decoder(16#6b#)) OR
 					(reg_q2652 AND symb_decoder(16#4b#));
reg_q2656_in <= (reg_q2654 AND symb_decoder(16#45#)) OR
 					(reg_q2654 AND symb_decoder(16#65#));
reg_q2607_in <= (reg_q2605 AND symb_decoder(16#45#)) OR
 					(reg_q2605 AND symb_decoder(16#65#));
reg_q1345_in <= (reg_q1343 AND symb_decoder(16#0d#)) OR
 					(reg_q1343 AND symb_decoder(16#0a#)) OR
 					(reg_q1343 AND symb_decoder(16#0c#)) OR
 					(reg_q1343 AND symb_decoder(16#09#)) OR
 					(reg_q1343 AND symb_decoder(16#20#)) OR
 					(reg_q1345 AND symb_decoder(16#0c#)) OR
 					(reg_q1345 AND symb_decoder(16#20#)) OR
 					(reg_q1345 AND symb_decoder(16#0a#)) OR
 					(reg_q1345 AND symb_decoder(16#09#)) OR
 					(reg_q1345 AND symb_decoder(16#0d#));
reg_q347_in <= (reg_q345 AND symb_decoder(16#4c#)) OR
 					(reg_q345 AND symb_decoder(16#6c#));
reg_q1488_in <= (reg_q1486 AND symb_decoder(16#3e#));
reg_q1286_in <= (reg_q1284 AND symb_decoder(16#4e#)) OR
 					(reg_q1284 AND symb_decoder(16#6e#));
reg_q321_in <= (reg_q319 AND symb_decoder(16#00#));
reg_q1508_in <= (reg_q1506 AND symb_decoder(16#45#)) OR
 					(reg_q1506 AND symb_decoder(16#65#));
reg_q1510_in <= (reg_q1508 AND symb_decoder(16#52#)) OR
 					(reg_q1508 AND symb_decoder(16#72#));
reg_q2099_in <= (reg_q2097 AND symb_decoder(16#49#)) OR
 					(reg_q2097 AND symb_decoder(16#69#));
reg_q70_in <= (reg_q68 AND symb_decoder(16#72#)) OR
 					(reg_q68 AND symb_decoder(16#52#));
reg_q970_in <= (reg_q968 AND symb_decoder(16#4c#)) OR
 					(reg_q968 AND symb_decoder(16#6c#));
reg_q760_in <= (reg_q758 AND symb_decoder(16#49#)) OR
 					(reg_q758 AND symb_decoder(16#69#));
reg_q762_in <= (reg_q760 AND symb_decoder(16#72#)) OR
 					(reg_q760 AND symb_decoder(16#52#));
reg_q707_in <= (reg_q705 AND symb_decoder(16#32#));
reg_q1234_in <= (reg_q1232 AND symb_decoder(16#63#)) OR
 					(reg_q1232 AND symb_decoder(16#43#));
reg_q1173_in <= (reg_q1171 AND symb_decoder(16#54#)) OR
 					(reg_q1171 AND symb_decoder(16#74#));
reg_q1175_in <= (reg_q1173 AND symb_decoder(16#49#)) OR
 					(reg_q1173 AND symb_decoder(16#69#));
reg_q2512_in <= (reg_q2510 AND symb_decoder(16#33#));
reg_q2652_in <= (reg_q2650 AND symb_decoder(16#0d#)) OR
 					(reg_q2650 AND symb_decoder(16#20#)) OR
 					(reg_q2650 AND symb_decoder(16#0c#)) OR
 					(reg_q2650 AND symb_decoder(16#0a#)) OR
 					(reg_q2650 AND symb_decoder(16#09#));
reg_q1584_in <= (reg_q1582 AND symb_decoder(16#0a#));
reg_q1006_in <= (reg_q1004 AND symb_decoder(16#29#));
reg_q1486_in <= (reg_q1484 AND symb_decoder(16#5c#));
reg_q331_in <= (reg_q329 AND symb_decoder(16#65#)) OR
 					(reg_q329 AND symb_decoder(16#45#));
reg_q1270_in <= (reg_q1268 AND symb_decoder(16#65#)) OR
 					(reg_q1268 AND symb_decoder(16#45#));
reg_q141_in <= (reg_q139 AND symb_decoder(16#43#)) OR
 					(reg_q139 AND symb_decoder(16#63#));
reg_q143_in <= (reg_q141 AND symb_decoder(16#74#)) OR
 					(reg_q141 AND symb_decoder(16#54#));
reg_q353_in <= (reg_q351 AND symb_decoder(16#65#)) OR
 					(reg_q351 AND symb_decoder(16#45#));
reg_q355_in <= (reg_q353 AND symb_decoder(16#52#)) OR
 					(reg_q353 AND symb_decoder(16#72#));
reg_q2668_in <= (reg_q2666 AND symb_decoder(16#49#)) OR
 					(reg_q2666 AND symb_decoder(16#69#));
reg_q72_in <= (reg_q70 AND symb_decoder(16#0d#)) OR
 					(reg_q70 AND symb_decoder(16#20#)) OR
 					(reg_q70 AND symb_decoder(16#0c#)) OR
 					(reg_q70 AND symb_decoder(16#0a#)) OR
 					(reg_q70 AND symb_decoder(16#09#)) OR
 					(reg_q72 AND symb_decoder(16#0c#)) OR
 					(reg_q72 AND symb_decoder(16#0a#)) OR
 					(reg_q72 AND symb_decoder(16#09#)) OR
 					(reg_q72 AND symb_decoder(16#20#)) OR
 					(reg_q72 AND symb_decoder(16#0d#));
reg_q165_in <= (reg_q163 AND symb_decoder(16#66#)) OR
 					(reg_q163 AND symb_decoder(16#46#));
reg_q1454_in <= (reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q1453 AND symb_decoder(16#48#)) OR
 					(reg_q1453 AND symb_decoder(16#68#));
reg_q1456_in <= (reg_q1454 AND symb_decoder(16#52#)) OR
 					(reg_q1454 AND symb_decoder(16#72#));
reg_q1607_in <= (reg_q1605 AND symb_decoder(16#49#)) OR
 					(reg_q1605 AND symb_decoder(16#69#));
reg_q1131_in <= (reg_q1129 AND symb_decoder(16#74#)) OR
 					(reg_q1129 AND symb_decoder(16#54#));
reg_q907_in <= (reg_q905 AND symb_decoder(16#6a#)) OR
 					(reg_q905 AND symb_decoder(16#4a#));
reg_q2254_in <= (reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2253 AND symb_decoder(16#21#));
reg_q2256_in <= (reg_q2254 AND symb_decoder(16#21#));
reg_q1629_in <= (reg_q1627 AND symb_decoder(16#49#)) OR
 					(reg_q1627 AND symb_decoder(16#69#));
reg_q1631_in <= (reg_q1629 AND symb_decoder(16#63#)) OR
 					(reg_q1629 AND symb_decoder(16#43#));
reg_q157_in <= (reg_q155 AND symb_decoder(16#43#)) OR
 					(reg_q155 AND symb_decoder(16#63#));
reg_q159_in <= (reg_q157 AND symb_decoder(16#45#)) OR
 					(reg_q157 AND symb_decoder(16#65#));
reg_q1590_in <= (reg_q1588 AND symb_decoder(16#52#)) OR
 					(reg_q1588 AND symb_decoder(16#72#));
reg_q1592_in <= (reg_q1590 AND symb_decoder(16#76#)) OR
 					(reg_q1590 AND symb_decoder(16#56#));
reg_q1564_in <= (reg_q1562 AND symb_decoder(16#72#)) OR
 					(reg_q1562 AND symb_decoder(16#52#));
reg_q1566_in <= (reg_q1564 AND symb_decoder(16#53#)) OR
 					(reg_q1564 AND symb_decoder(16#73#));
reg_q1720_in <= (reg_q1720 AND symb_decoder(16#0a#)) OR
 					(reg_q1720 AND symb_decoder(16#0d#)) OR
 					(reg_q1720 AND symb_decoder(16#09#)) OR
 					(reg_q1720 AND symb_decoder(16#20#)) OR
 					(reg_q1720 AND symb_decoder(16#0c#)) OR
 					(reg_q1718 AND symb_decoder(16#0c#)) OR
 					(reg_q1718 AND symb_decoder(16#0d#)) OR
 					(reg_q1718 AND symb_decoder(16#09#)) OR
 					(reg_q1718 AND symb_decoder(16#0a#)) OR
 					(reg_q1718 AND symb_decoder(16#20#));
reg_q1722_in <= (reg_q1720 AND symb_decoder(16#59#)) OR
 					(reg_q1720 AND symb_decoder(16#79#));
reg_q2006_in <= (reg_q2004 AND symb_decoder(16#54#)) OR
 					(reg_q2004 AND symb_decoder(16#74#));
reg_q1965_in <= (reg_q1963 AND symb_decoder(16#65#)) OR
 					(reg_q1963 AND symb_decoder(16#45#));
reg_q1967_in <= (reg_q1965 AND symb_decoder(16#52#)) OR
 					(reg_q1965 AND symb_decoder(16#72#));
reg_q272_in <= (reg_q270 AND symb_decoder(16#31#));
reg_q274_in <= (reg_q272 AND symb_decoder(16#20#));
reg_q2264_in <= (reg_q2262 AND symb_decoder(16#74#)) OR
 					(reg_q2262 AND symb_decoder(16#54#));
reg_q2266_in <= (reg_q2264 AND symb_decoder(16#69#)) OR
 					(reg_q2264 AND symb_decoder(16#49#));
reg_q204_in <= (reg_q202 AND symb_decoder(16#76#)) OR
 					(reg_q202 AND symb_decoder(16#56#));
reg_q206_in <= (reg_q204 AND symb_decoder(16#72#)) OR
 					(reg_q204 AND symb_decoder(16#52#));
reg_q1311_in <= (reg_q1309 AND symb_decoder(16#69#)) OR
 					(reg_q1309 AND symb_decoder(16#49#));
reg_q909_in <= (reg_q907 AND symb_decoder(16#55#)) OR
 					(reg_q907 AND symb_decoder(16#75#));
reg_q911_in <= (reg_q909 AND symb_decoder(16#73#)) OR
 					(reg_q909 AND symb_decoder(16#53#));
reg_q2164_in <= (reg_q2162 AND symb_decoder(16#41#)) OR
 					(reg_q2162 AND symb_decoder(16#61#));
reg_q2166_in <= (reg_q2164 AND symb_decoder(16#45#)) OR
 					(reg_q2164 AND symb_decoder(16#65#));
reg_q1098_in <= (reg_q1096 AND symb_decoder(16#70#)) OR
 					(reg_q1096 AND symb_decoder(16#50#));
reg_q2563_in <= (reg_q2561 AND symb_decoder(16#64#)) OR
 					(reg_q2561 AND symb_decoder(16#44#));
reg_q2121_in <= (reg_q2119 AND symb_decoder(16#72#)) OR
 					(reg_q2119 AND symb_decoder(16#52#));
reg_q151_in <= (reg_q149 AND symb_decoder(16#53#)) OR
 					(reg_q149 AND symb_decoder(16#73#));
reg_q1121_in <= (reg_q1119 AND symb_decoder(16#45#)) OR
 					(reg_q1119 AND symb_decoder(16#65#));
reg_q243_in <= (reg_q241 AND symb_decoder(16#ff#));
reg_q1043_in <= (reg_q1041 AND symb_decoder(16#56#)) OR
 					(reg_q1041 AND symb_decoder(16#76#));
reg_q1045_in <= (reg_q1043 AND symb_decoder(16#65#)) OR
 					(reg_q1043 AND symb_decoder(16#45#));
reg_q276_in <= (reg_q274 AND symb_decoder(16#64#)) OR
 					(reg_q274 AND symb_decoder(16#44#));
reg_q1047_in <= (reg_q1045 AND symb_decoder(16#52#)) OR
 					(reg_q1045 AND symb_decoder(16#72#));
reg_q2367_in <= (reg_q2365 AND symb_decoder(16#22#));
reg_q1066_in <= (reg_q1064 AND symb_decoder(16#45#)) OR
 					(reg_q1064 AND symb_decoder(16#65#));
reg_q1496_in <= (reg_q1494 AND symb_decoder(16#72#)) OR
 					(reg_q1494 AND symb_decoder(16#52#));
reg_q1498_in <= (reg_q1496 AND symb_decoder(16#76#)) OR
 					(reg_q1496 AND symb_decoder(16#56#));
reg_q1696_in <= (reg_q1694 AND symb_decoder(16#55#)) OR
 					(reg_q1694 AND symb_decoder(16#75#));
reg_q1494_in <= (reg_q1492 AND symb_decoder(16#45#)) OR
 					(reg_q1492 AND symb_decoder(16#65#));
reg_q2036_in <= (reg_q2034 AND symb_decoder(16#4c#)) OR
 					(reg_q2034 AND symb_decoder(16#6c#));
reg_q1684_in <= (reg_q1682 AND symb_decoder(16#77#)) OR
 					(reg_q1682 AND symb_decoder(16#57#));
reg_q337_in <= (reg_q335 AND symb_decoder(16#6f#)) OR
 					(reg_q335 AND symb_decoder(16#4f#));
reg_q339_in <= (reg_q337 AND symb_decoder(16#6e#)) OR
 					(reg_q337 AND symb_decoder(16#4e#));
reg_q1959_in <= (reg_q1957 AND symb_decoder(16#49#)) OR
 					(reg_q1957 AND symb_decoder(16#69#));
reg_q1961_in <= (reg_q1959 AND symb_decoder(16#23#));
reg_q1518_in <= (reg_q1516 AND symb_decoder(16#4e#)) OR
 					(reg_q1516 AND symb_decoder(16#6e#));
reg_q1656_in <= (reg_q1654 AND symb_decoder(16#36#));
reg_q1658_in <= (reg_q1656 AND symb_decoder(16#36#));
reg_q2314_in <= (reg_q2312 AND symb_decoder(16#45#)) OR
 					(reg_q2312 AND symb_decoder(16#65#));
reg_q2316_in <= (reg_q2314 AND symb_decoder(16#21#));
reg_q2638_in <= (reg_q2636 AND symb_decoder(16#65#)) OR
 					(reg_q2636 AND symb_decoder(16#45#));
reg_q2142_in <= (reg_q2140 AND symb_decoder(16#68#)) OR
 					(reg_q2140 AND symb_decoder(16#48#));
reg_q2660_in <= (reg_q2658 AND symb_decoder(16#6c#)) OR
 					(reg_q2658 AND symb_decoder(16#4c#));
reg_q1568_in <= (reg_q1566 AND symb_decoder(16#69#)) OR
 					(reg_q1566 AND symb_decoder(16#49#));
reg_q1062_in <= (reg_q1060 AND symb_decoder(16#69#)) OR
 					(reg_q1060 AND symb_decoder(16#49#));
reg_q1064_in <= (reg_q1062 AND symb_decoder(16#54#)) OR
 					(reg_q1062 AND symb_decoder(16#74#));
reg_q1686_in <= (reg_q1684 AND symb_decoder(16#61#)) OR
 					(reg_q1684 AND symb_decoder(16#41#));
reg_q1240_in <= (reg_q1238 AND symb_decoder(16#53#)) OR
 					(reg_q1238 AND symb_decoder(16#73#));
reg_q764_in <= (reg_q762 AND symb_decoder(16#45#)) OR
 					(reg_q762 AND symb_decoder(16#65#));
reg_q1119_in <= (reg_q1117 AND symb_decoder(16#63#)) OR
 					(reg_q1117 AND symb_decoder(16#43#));
reg_q1476_in <= (reg_q1474 AND symb_decoder(16#41#)) OR
 					(reg_q1474 AND symb_decoder(16#61#));
reg_q62_in <= (reg_q60 AND symb_decoder(16#43#)) OR
 					(reg_q60 AND symb_decoder(16#63#));
reg_q2678_in <= (reg_q2676 AND symb_decoder(16#54#)) OR
 					(reg_q2676 AND symb_decoder(16#74#));
reg_q327_in <= (reg_q325 AND symb_decoder(16#00#));
reg_q329_in <= (reg_q327 AND symb_decoder(16#4e#)) OR
 					(reg_q327 AND symb_decoder(16#6e#));
reg_q1718_in <= (reg_q1716 AND symb_decoder(16#2e#));
reg_q1054_in <= (reg_q1052 AND symb_decoder(16#58#)) OR
 					(reg_q1052 AND symb_decoder(16#78#));
reg_q1056_in <= (reg_q1054 AND symb_decoder(16#50#)) OR
 					(reg_q1054 AND symb_decoder(16#70#));
reg_q1512_in <= (reg_q1510 AND symb_decoder(16#53#)) OR
 					(reg_q1510 AND symb_decoder(16#73#));
reg_q2262_in <= (reg_q2260 AND symb_decoder(16#50#)) OR
 					(reg_q2260 AND symb_decoder(16#70#));
reg_q1167_in <= (reg_q1165 AND symb_decoder(16#6e#)) OR
 					(reg_q1165 AND symb_decoder(16#4e#));
reg_q2379_in <= (reg_q2377 AND symb_decoder(16#0d#));
reg_q2016_in <= (reg_q2014 AND symb_decoder(16#46#)) OR
 					(reg_q2014 AND symb_decoder(16#66#));
reg_q64_in <= (reg_q62 AND symb_decoder(16#48#)) OR
 					(reg_q62 AND symb_decoder(16#68#));
reg_q1623_in <= (reg_q1621 AND symb_decoder(16#6b#)) OR
 					(reg_q1621 AND symb_decoder(16#4b#));
reg_q145_in <= (reg_q143 AND symb_decoder(16#65#)) OR
 					(reg_q143 AND symb_decoder(16#45#));
reg_q1594_in <= (reg_q1592 AND symb_decoder(16#69#)) OR
 					(reg_q1592 AND symb_decoder(16#49#));
reg_q1596_in <= (reg_q1594 AND symb_decoder(16#63#)) OR
 					(reg_q1594 AND symb_decoder(16#43#));
reg_q2626_in <= (reg_q2624 AND symb_decoder(16#61#)) OR
 					(reg_q2624 AND symb_decoder(16#41#));
reg_q2365_in <= (reg_q2363 AND symb_decoder(16#72#)) OR
 					(reg_q2363 AND symb_decoder(16#52#));
reg_q1609_in <= (reg_q1607 AND symb_decoder(16#63#)) OR
 					(reg_q1607 AND symb_decoder(16#43#));
reg_q1058_in <= (reg_q1056 AND symb_decoder(16#4c#)) OR
 					(reg_q1056 AND symb_decoder(16#6c#));
reg_q1060_in <= (reg_q1058 AND symb_decoder(16#6f#)) OR
 					(reg_q1058 AND symb_decoder(16#4f#));
reg_q208_in <= (reg_q206 AND symb_decoder(16#5e#));
reg_q1621_in <= (reg_q1619 AND symb_decoder(16#61#)) OR
 					(reg_q1619 AND symb_decoder(16#41#));
reg_q694_in <= (reg_q692 AND symb_decoder(16#2e#));
reg_q214_in <= (reg_q212 AND symb_decoder(16#45#)) OR
 					(reg_q212 AND symb_decoder(16#65#));
reg_q2555_in <= (reg_q2553 AND symb_decoder(16#74#)) OR
 					(reg_q2553 AND symb_decoder(16#54#));
reg_q2152_in <= (reg_q2150 AND symb_decoder(16#72#)) OR
 					(reg_q2150 AND symb_decoder(16#52#));
reg_q2154_in <= (reg_q2152 AND symb_decoder(16#45#)) OR
 					(reg_q2152 AND symb_decoder(16#65#));
reg_q2312_in <= (reg_q2310 AND symb_decoder(16#6e#)) OR
 					(reg_q2310 AND symb_decoder(16#4e#));
reg_q311_in <= (reg_q309 AND symb_decoder(16#77#)) OR
 					(reg_q309 AND symb_decoder(16#57#));
reg_q1500_in <= (reg_q1498 AND symb_decoder(16#45#)) OR
 					(reg_q1498 AND symb_decoder(16#65#));
reg_q317_in <= (reg_q315 AND symb_decoder(16#00#));
reg_q2680_in <= (reg_q2678 AND symb_decoder(16#61#)) OR
 					(reg_q2678 AND symb_decoder(16#41#));
reg_q1266_in <= (reg_q1264 AND symb_decoder(16#52#)) OR
 					(reg_q1264 AND symb_decoder(16#72#));
reg_q1268_in <= (reg_q1266 AND symb_decoder(16#56#)) OR
 					(reg_q1266 AND symb_decoder(16#76#));
reg_q2628_in <= (reg_q2626 AND symb_decoder(16#74#)) OR
 					(reg_q2626 AND symb_decoder(16#54#));
reg_q2630_in <= (reg_q2628 AND symb_decoder(16#75#)) OR
 					(reg_q2628 AND symb_decoder(16#55#));
reg_q1429_in <= (reg_q1427 AND symb_decoder(16#54#)) OR
 					(reg_q1427 AND symb_decoder(16#74#));
reg_q1236_in <= (reg_q1234 AND symb_decoder(16#72#)) OR
 					(reg_q1234 AND symb_decoder(16#52#));
reg_q1238_in <= (reg_q1236 AND symb_decoder(16#61#)) OR
 					(reg_q1236 AND symb_decoder(16#41#));
reg_q2478_in <= (reg_q2476 AND symb_decoder(16#31#));
reg_q722_in <= (reg_q720 AND symb_decoder(16#65#)) OR
 					(reg_q720 AND symb_decoder(16#45#));
reg_q391_in <= (reg_q389 AND symb_decoder(16#45#)) OR
 					(reg_q389 AND symb_decoder(16#65#));
reg_q393_in <= (reg_q391 AND symb_decoder(16#4e#)) OR
 					(reg_q391 AND symb_decoder(16#6e#));
reg_q1280_in <= (reg_q1278 AND symb_decoder(16#2d#));
reg_q2569_in <= (reg_q2567 AND symb_decoder(16#57#)) OR
 					(reg_q2567 AND symb_decoder(16#77#));
reg_q202_in <= (reg_q200 AND symb_decoder(16#73#)) OR
 					(reg_q200 AND symb_decoder(16#53#));
reg_q268_in <= (reg_q266 AND symb_decoder(16#33#));
reg_q270_in <= (reg_q268 AND symb_decoder(16#31#));
reg_q173_in <= (reg_q171 AND symb_decoder(16#79#)) OR
 					(reg_q171 AND symb_decoder(16#59#));
reg_q175_in <= (reg_q173 AND symb_decoder(16#21#));
reg_q669_in <= (reg_q667 AND symb_decoder(16#6f#)) OR
 					(reg_q667 AND symb_decoder(16#4f#));
reg_q1502_in <= (reg_q1500 AND symb_decoder(16#52#)) OR
 					(reg_q1500 AND symb_decoder(16#72#));
reg_q738_in <= (reg_q736 AND symb_decoder(16#6f#)) OR
 					(reg_q736 AND symb_decoder(16#4f#));
reg_q54_in <= (reg_q52 AND symb_decoder(16#4f#)) OR
 					(reg_q52 AND symb_decoder(16#6f#));
reg_q1963_in <= (reg_q1961 AND symb_decoder(16#73#)) OR
 					(reg_q1961 AND symb_decoder(16#53#));
reg_q2381_in <= (reg_q2379 AND symb_decoder(16#0a#));
reg_q2345_in <= (reg_q2343 AND symb_decoder(16#4f#)) OR
 					(reg_q2343 AND symb_decoder(16#6f#));
reg_q2008_in <= (reg_q2006 AND symb_decoder(16#72#)) OR
 					(reg_q2006 AND symb_decoder(16#52#));
reg_q730_in <= (reg_q728 AND symb_decoder(16#4e#)) OR
 					(reg_q728 AND symb_decoder(16#6e#));
reg_q1321_in <= (reg_q1319 AND symb_decoder(16#53#)) OR
 					(reg_q1319 AND symb_decoder(16#73#));
reg_q1323_in <= (reg_q1321 AND symb_decoder(16#45#)) OR
 					(reg_q1321 AND symb_decoder(16#65#));
reg_q1309_in <= (reg_q1307 AND symb_decoder(16#72#)) OR
 					(reg_q1307 AND symb_decoder(16#52#));
reg_q99_in <= (reg_q97 AND symb_decoder(16#ac#));
reg_q1586_in <= (reg_q1584 AND symb_decoder(16#73#)) OR
 					(reg_q1584 AND symb_decoder(16#53#));
reg_q2156_in <= (reg_q2154 AND symb_decoder(16#61#)) OR
 					(reg_q2154 AND symb_decoder(16#41#));
reg_q319_in <= (reg_q317 AND symb_decoder(16#00#));
reg_q2026_in <= (reg_q2024 AND symb_decoder(16#6e#)) OR
 					(reg_q2024 AND symb_decoder(16#4e#));
reg_q401_in <= (reg_q399 AND symb_decoder(16#52#)) OR
 					(reg_q399 AND symb_decoder(16#72#));
reg_q2666_in <= (reg_q2664 AND symb_decoder(16#47#)) OR
 					(reg_q2664 AND symb_decoder(16#67#));
reg_q286_in <= (reg_q284 AND symb_decoder(16#20#));
reg_q2658_in <= (reg_q2656 AND symb_decoder(16#59#)) OR
 					(reg_q2656 AND symb_decoder(16#79#));
reg_q754_in <= (reg_q752 AND symb_decoder(16#46#)) OR
 					(reg_q752 AND symb_decoder(16#66#));
reg_q345_in <= (reg_q343 AND symb_decoder(16#6f#)) OR
 					(reg_q343 AND symb_decoder(16#4f#));
reg_q1021_in <= (reg_q1019 AND symb_decoder(16#7a#)) OR
 					(reg_q1019 AND symb_decoder(16#5a#));
reg_q2539_in <= (reg_q2537 AND symb_decoder(16#66#)) OR
 					(reg_q2537 AND symb_decoder(16#46#));
reg_q1163_in <= (reg_q1161 AND symb_decoder(16#4f#)) OR
 					(reg_q1161 AND symb_decoder(16#6f#));
reg_q1165_in <= (reg_q1163 AND symb_decoder(16#4e#)) OR
 					(reg_q1163 AND symb_decoder(16#6e#));
reg_q411_in <= (reg_q409 AND symb_decoder(16#54#)) OR
 					(reg_q409 AND symb_decoder(16#74#));
reg_q720_in <= (reg_q718 AND symb_decoder(16#47#)) OR
 					(reg_q718 AND symb_decoder(16#67#));
reg_q1292_in <= (reg_q1290 AND symb_decoder(16#2e#));
reg_q1294_in <= (reg_q1292 AND symb_decoder(16#2e#));
reg_q2553_in <= (reg_q2551 AND symb_decoder(16#73#)) OR
 					(reg_q2551 AND symb_decoder(16#53#));
reg_q1449_in <= (reg_q1447 AND symb_decoder(16#6d#)) OR
 					(reg_q1447 AND symb_decoder(16#4d#));
reg_q1100_in <= (reg_q1098 AND symb_decoder(16#4f#)) OR
 					(reg_q1098 AND symb_decoder(16#6f#));
reg_q424_in <= (reg_q422 AND symb_decoder(16#65#)) OR
 					(reg_q422 AND symb_decoder(16#45#));
reg_q1177_in <= (reg_q1175 AND symb_decoder(16#6f#)) OR
 					(reg_q1175 AND symb_decoder(16#4f#));
reg_q2355_in <= (reg_q2353 AND symb_decoder(16#41#)) OR
 					(reg_q2353 AND symb_decoder(16#61#));
reg_q732_in <= (reg_q730 AND symb_decoder(16#67#)) OR
 					(reg_q730 AND symb_decoder(16#47#));
reg_q434_in <= (reg_q432 AND symb_decoder(16#4e#)) OR
 					(reg_q432 AND symb_decoder(16#6e#));
reg_q2551_in <= (reg_q2549 AND symb_decoder(16#69#)) OR
 					(reg_q2549 AND symb_decoder(16#49#));
reg_q2044_in <= (reg_q2042 AND symb_decoder(16#72#)) OR
 					(reg_q2042 AND symb_decoder(16#52#));
reg_q2046_in <= (reg_q2044 AND symb_decoder(16#6f#)) OR
 					(reg_q2044 AND symb_decoder(16#4f#));
reg_q2541_in <= (reg_q2539 AND symb_decoder(16#6f#)) OR
 					(reg_q2539 AND symb_decoder(16#4f#));
reg_q1588_in <= (reg_q1586 AND symb_decoder(16#45#)) OR
 					(reg_q1586 AND symb_decoder(16#65#));
reg_q2693_in <= (reg_q2692 AND symb_decoder(16#0d#));
reg_q2543_in <= (reg_q2541 AND symb_decoder(16#2c#));
reg_q2545_in <= (reg_q2543 AND symb_decoder(16#72#)) OR
 					(reg_q2543 AND symb_decoder(16#52#));
reg_q2347_in <= (reg_q2345 AND symb_decoder(16#54#)) OR
 					(reg_q2345 AND symb_decoder(16#74#));
reg_q1740_in <= (reg_q1738 AND symb_decoder(16#73#)) OR
 					(reg_q1738 AND symb_decoder(16#53#));
reg_q1329_in <= (reg_q1327 AND symb_decoder(16#45#)) OR
 					(reg_q1327 AND symb_decoder(16#65#));
reg_q2632_in <= (reg_q2630 AND symb_decoder(16#73#)) OR
 					(reg_q2630 AND symb_decoder(16#53#));
reg_q1303_in <= (reg_q1301 AND symb_decoder(16#52#)) OR
 					(reg_q1301 AND symb_decoder(16#72#));
reg_q309_in <= (reg_q307 AND symb_decoder(16#53#)) OR
 					(reg_q307 AND symb_decoder(16#73#));
reg_q216_in <= (reg_q214 AND symb_decoder(16#72#)) OR
 					(reg_q214 AND symb_decoder(16#52#));
reg_q2134_in <= (reg_q2132 AND symb_decoder(16#4f#)) OR
 					(reg_q2132 AND symb_decoder(16#6f#));
reg_q770_in <= (reg_q768 AND symb_decoder(16#6f#)) OR
 					(reg_q768 AND symb_decoder(16#4f#));
reg_q155_in <= (reg_q153 AND symb_decoder(16#63#)) OR
 					(reg_q153 AND symb_decoder(16#43#));
reg_q2140_in <= (reg_q2138 AND symb_decoder(16#54#)) OR
 					(reg_q2138 AND symb_decoder(16#74#));
reg_q383_in <= (reg_q381 AND symb_decoder(16#75#)) OR
 					(reg_q381 AND symb_decoder(16#55#));
reg_q1633_in <= (reg_q1631 AND symb_decoder(16#74#)) OR
 					(reg_q1631 AND symb_decoder(16#54#));
reg_q772_in <= (reg_q770 AND symb_decoder(16#72#)) OR
 					(reg_q770 AND symb_decoder(16#52#));
reg_q1155_in <= (reg_q1153 AND symb_decoder(16#0a#));
reg_q927_in <= (reg_q925 AND symb_decoder(16#76#)) OR
 					(reg_q925 AND symb_decoder(16#56#));
reg_q929_in <= (reg_q927 AND symb_decoder(16#65#)) OR
 					(reg_q927 AND symb_decoder(16#45#));
reg_q1969_in <= (reg_q1967 AND symb_decoder(16#56#)) OR
 					(reg_q1967 AND symb_decoder(16#76#));
reg_q1415_in <= (reg_q1413 AND symb_decoder(16#0d#));
reg_q1417_in <= (reg_q1415 AND symb_decoder(16#0a#));
reg_q153_in <= (reg_q151 AND symb_decoder(16#55#)) OR
 					(reg_q151 AND symb_decoder(16#75#));
reg_q1288_in <= (reg_q1286 AND symb_decoder(16#65#)) OR
 					(reg_q1286 AND symb_decoder(16#45#));
reg_q1276_in <= (reg_q1274 AND symb_decoder(16#4f#)) OR
 					(reg_q1274 AND symb_decoder(16#6f#));
reg_q2048_in <= (reg_q2046 AND symb_decoder(16#6d#)) OR
 					(reg_q2046 AND symb_decoder(16#4d#));
reg_q218_in <= (reg_q216 AND symb_decoder(16#4c#)) OR
 					(reg_q216 AND symb_decoder(16#6c#));
reg_q1149_in <= (reg_q1147 AND symb_decoder(16#0d#));
reg_q259_in <= (reg_q257 AND symb_decoder(16#ff#));
reg_q2327_in <= (reg_q2325 AND symb_decoder(16#57#)) OR
 					(reg_q2325 AND symb_decoder(16#77#));
reg_q266_in <= (reg_q264 AND symb_decoder(16#2d#));
reg_q746_in <= (reg_q744 AND symb_decoder(16#6e#)) OR
 					(reg_q744 AND symb_decoder(16#4e#));
reg_q774_in <= (reg_q772 AND symb_decoder(16#79#)) OR
 					(reg_q772 AND symb_decoder(16#59#));
reg_q776_in <= (reg_q774 AND symb_decoder(16#3a#));
reg_q389_in <= (reg_q387 AND symb_decoder(16#45#)) OR
 					(reg_q387 AND symb_decoder(16#65#));
reg_q1598_in <= (reg_q1596 AND symb_decoder(16#65#)) OR
 					(reg_q1596 AND symb_decoder(16#45#));
reg_q1004_in <= (reg_q1002 AND symb_decoder(16#3a#));
reg_q1419_in <= (reg_q1417 AND symb_decoder(16#6f#)) OR
 					(reg_q1417 AND symb_decoder(16#4f#));
reg_q1278_in <= (reg_q1276 AND symb_decoder(16#6e#)) OR
 					(reg_q1276 AND symb_decoder(16#4e#));
reg_q1654_in <= (reg_q1652 AND symb_decoder(16#36#));
reg_q1458_in <= (reg_q1456 AND symb_decoder(16#41#)) OR
 					(reg_q1456 AND symb_decoder(16#61#));
reg_q1641_in <= (reg_q1639 AND symb_decoder(16#0a#));
reg_q1600_in <= (reg_q1598 AND symb_decoder(16#3a#));
reg_q2097_in <= (reg_q2095 AND symb_decoder(16#49#)) OR
 					(reg_q2095 AND symb_decoder(16#69#));
reg_q1290_in <= (reg_q1288 AND symb_decoder(16#2e#));
reg_q740_in <= (reg_q738 AND symb_decoder(16#6e#)) OR
 					(reg_q738 AND symb_decoder(16#4e#));
reg_q677_in <= (reg_q675 AND symb_decoder(16#5c#));
reg_q2050_in <= (reg_q2048 AND symb_decoder(16#3a#));
reg_fullgraph2_init <= "0000000000";

reg_fullgraph2_sel <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & reg_q2050_in & reg_q677_in & reg_q740_in & reg_q1290_in & reg_q2097_in & reg_q1600_in & reg_q1641_in & reg_q1458_in & reg_q1654_in & reg_q1278_in & reg_q1419_in & reg_q1004_in & reg_q1598_in & reg_q389_in & reg_q776_in & reg_q774_in & reg_q746_in & reg_q266_in & reg_q2327_in & reg_q259_in & reg_q1149_in & reg_q218_in & reg_q2048_in & reg_q1276_in & reg_q1288_in & reg_q153_in & reg_q1417_in & reg_q1415_in & reg_q1969_in & reg_q929_in & reg_q927_in & reg_q1155_in & reg_q772_in & reg_q1633_in & reg_q383_in & reg_q2140_in & reg_q155_in & reg_q770_in & reg_q2134_in & reg_q216_in & reg_q309_in & reg_q1303_in & reg_q2632_in & reg_q1329_in & reg_q1740_in & reg_q2347_in & reg_q2545_in & reg_q2543_in & reg_q2693_in & reg_q1588_in & reg_q2541_in & reg_q2046_in & reg_q2044_in & reg_q2551_in & reg_q434_in & reg_q732_in & reg_q2355_in & reg_q1177_in & reg_q424_in & reg_q1100_in & reg_q1449_in & reg_q2553_in & reg_q1294_in & reg_q1292_in & reg_q720_in & reg_q411_in & reg_q1165_in & reg_q1163_in & reg_q2539_in & reg_q1021_in & reg_q345_in & reg_q754_in & reg_q2658_in & reg_q286_in & reg_q2666_in & reg_q401_in & reg_q2026_in & reg_q319_in & reg_q2156_in & reg_q1586_in & reg_q99_in & reg_q1309_in & reg_q1323_in & reg_q1321_in & reg_q730_in & reg_q2008_in & reg_q2345_in & reg_q2381_in & reg_q1963_in & reg_q54_in & reg_q738_in & reg_q1502_in & reg_q669_in & reg_q175_in & reg_q173_in & reg_q270_in & reg_q268_in & reg_q202_in & reg_q2569_in & reg_q1280_in & reg_q393_in & reg_q391_in & reg_q722_in & reg_q2478_in & reg_q1238_in & reg_q1236_in & reg_q1429_in & reg_q2630_in & reg_q2628_in & reg_q1268_in & reg_q1266_in & reg_q2680_in & reg_q317_in & reg_q1500_in & reg_q311_in & reg_q2312_in & reg_q2154_in & reg_q2152_in & reg_q2555_in & reg_q214_in & reg_q694_in & reg_q1621_in & reg_q208_in & reg_q1060_in & reg_q1058_in & reg_q1609_in & reg_q2365_in & reg_q2626_in & reg_q1596_in & reg_q1594_in & reg_q145_in & reg_q1623_in & reg_q64_in & reg_q2016_in & reg_q2379_in & reg_q1167_in & reg_q2262_in & reg_q1512_in & reg_q1056_in & reg_q1054_in & reg_q1718_in & reg_q329_in & reg_q327_in & reg_q2678_in & reg_q62_in & reg_q1476_in & reg_q1119_in & reg_q764_in & reg_q1240_in & reg_q1686_in & reg_q1064_in & reg_q1062_in & reg_q1568_in & reg_q2660_in & reg_q2142_in & reg_q2638_in & reg_q2316_in & reg_q2314_in & reg_q1658_in & reg_q1656_in & reg_q1518_in & reg_q1961_in & reg_q1959_in & reg_q339_in & reg_q337_in & reg_q1684_in & reg_q2036_in & reg_q1494_in & reg_q1696_in & reg_q1498_in & reg_q1496_in & reg_q1066_in & reg_q2367_in & reg_q1047_in & reg_q276_in & reg_q1045_in & reg_q1043_in & reg_q243_in & reg_q1121_in & reg_q151_in & reg_q2121_in & reg_q2563_in & reg_q1098_in & reg_q2166_in & reg_q2164_in & reg_q911_in & reg_q909_in & reg_q1311_in & reg_q206_in & reg_q204_in & reg_q2266_in & reg_q2264_in & reg_q274_in & reg_q272_in & reg_q1967_in & reg_q1965_in & reg_q2006_in & reg_q1722_in & reg_q1720_in & reg_q1566_in & reg_q1564_in & reg_q1592_in & reg_q1590_in & reg_q159_in & reg_q157_in & reg_q1631_in & reg_q1629_in & reg_q2256_in & reg_q2254_in & reg_q907_in & reg_q1131_in & reg_q1607_in & reg_q1456_in & reg_q1454_in & reg_q165_in & reg_q72_in & reg_q2668_in & reg_q355_in & reg_q353_in & reg_q143_in & reg_q141_in & reg_q1270_in & reg_q331_in & reg_q1486_in & reg_q1006_in & reg_q1584_in & reg_q2652_in & reg_q2512_in & reg_q1175_in & reg_q1173_in & reg_q1234_in & reg_q707_in & reg_q762_in & reg_q760_in & reg_q970_in & reg_q70_in & reg_q2099_in & reg_q1510_in & reg_q1508_in & reg_q321_in & reg_q1286_in & reg_q1488_in & reg_q347_in & reg_q1345_in & reg_q2607_in & reg_q2656_in & reg_q2654_in & reg_q1157_in & reg_q2331_in & reg_q2329_in & reg_q728_in & reg_q2107_in & reg_q1516_in & reg_q1514_in & reg_q2684_in & reg_q2682_in & reg_q2320_in & reg_q2318_in & reg_q432_in & reg_q387_in & reg_q385_in & reg_q1351_in & reg_q1129_in & reg_q1127_in & reg_q1353_in & reg_q2561_in & reg_q1615_in & reg_q2571_in & reg_q1019_in & reg_q1017_in & reg_q1171_in & reg_q1169_in & reg_q1611_in & reg_q296_in & reg_q147_in & reg_q1650_in & reg_q1228_in & reg_q2146_in & reg_q2144_in & reg_q2113_in & reg_q726_in & reg_q724_in & reg_q2231_in & reg_q2495_in & reg_q1554_in & reg_q1492_in & reg_q2219_in & reg_q972_in & reg_q2235_in & reg_q2233_in & reg_q2241_in & reg_q1041_in & reg_q1039_in & reg_q684_in & reg_q80_in & reg_q78_in & reg_q212_in & reg_q210_in & reg_q222_in & reg_q220_in & reg_q436_in & reg_q1706_in & reg_q1572_in & reg_q1570_in & reg_q1284_in & reg_q1282_in & reg_q1244_in & reg_q1242_in & reg_q2239_in & reg_q2237_in & reg_q1533_in & reg_q2290_in & reg_q307_in & reg_q1648_in & reg_q351_in & reg_q349_in & reg_q1627_in & reg_q1625_in & reg_q1343_in & reg_q2148_in & reg_q105_in & reg_q278_in & reg_q239_in & reg_q171_in & reg_q2095_in & reg_q284_in & reg_q1078_in & reg_q1076_in & reg_q2650_in & reg_q399_in & reg_q60_in & reg_q667_in & reg_q2339_in & reg_q1613_in & reg_q1125_in & reg_q1123_in & reg_q2573_in & reg_q962_in & reg_q1185_in & reg_q1183_in & reg_q446_in & reg_q444_in & reg_q1159_in & reg_q2298_in & reg_q2296_in & reg_q2502_in & reg_q2014_in & reg_q1447_in & reg_q734_in & reg_q1260_in & reg_q1258_in & reg_q1619_in & reg_q1617_in & reg_q2559_in & reg_q2557_in & reg_q1068_in & reg_q2012_in & reg_q2010_in & reg_q1141_in & reg_q139_in & reg_q2664_in & reg_q2662_in & reg_q768_in & reg_q766_in & reg_q430_in & reg_q2034_in & reg_q2032_in & reg_q2270_in & reg_q2268_in & reg_q2300_in & reg_q68_in & reg_q66_in & reg_q1474_in & reg_q1254_in & reg_q2648_in & reg_q2646_in & reg_q1232_in & reg_q1230_in & reg_q88_in & reg_q200_in & reg_q2472_in & reg_q2470_in & reg_q409_in & reg_q407_in & reg_q1712_in & reg_q1710_in & reg_q438_in & reg_q1070_in & reg_q2549_in & reg_q2547_in & reg_q163_in & reg_q161_in & reg_q1539_in & reg_q696_in & reg_q300_in & reg_q298_in & reg_q992_in & reg_q976_in & reg_q974_in & reg_q2624_in & reg_q1033_in & reg_q1256_in & reg_q1313_in & reg_q241_in & reg_q2640_in & reg_q2105_in & reg_q2359_in & reg_q2357_in & reg_q1439_in & reg_q1558_in & reg_q1556_in & reg_q315_in & reg_q313_in & reg_q1537_in & reg_q1535_in & reg_q2282_in & reg_q2280_in & reg_q2130_in & reg_q1490_in & reg_q2288_in & reg_q1445_in & reg_q752_in & reg_q1246_in & reg_q405_in & reg_q403_in & reg_q442_in & reg_q440_in & reg_q2676_in & reg_q2674_in & reg_q1484_in & reg_q2160_in & reg_q2158_in & reg_q282_in & reg_q280_in & reg_q82_in & reg_q986_in & reg_q1319_in & reg_q2306_in & reg_q2304_in & reg_q913_in & reg_q1181_in & reg_q1179_in & reg_q1552_in & reg_q1973_in & reg_q1971_in & reg_q1153_in & reg_q1151_in & reg_q1728_in & reg_q1652_in & reg_q377_in & reg_q1666_in & reg_q1664_in & reg_q294_in & reg_q292_in & reg_q325_in & reg_q323_in & reg_q1635_in & reg_q925_in & reg_q923_in & reg_q2499_in & reg_q2497_in & reg_q1506_in & reg_q1504_in & reg_q1274_in & reg_q1272_in & reg_q2575_in & reg_q1133_in & reg_q1025_in & reg_q1023_in & reg_q2349_in & reg_q2686_in & reg_q1264_in & reg_q1262_in & reg_q1692_in & reg_q1435_in & reg_q750_in & reg_q748_in & reg_q964_in & reg_q1437_in & reg_q698_in & reg_q365_in & reg_q86_in & reg_q84_in & reg_q397_in & reg_q395_in & reg_q192_in & reg_q448_in & reg_q1117_in & reg_q1115_in & reg_q1349_in & reg_q1347_in & reg_q1092_in & reg_q785_in & reg_q783_in & reg_q109_in & reg_q107_in & reg_q1639_in & reg_q1637_in & reg_q2601_in & reg_q2599_in & reg_q2644_in & reg_q2642_in & reg_q1672_in & reg_q1010_in & reg_q1008_in & reg_q915_in & reg_q255_in & reg_q119_in & reg_q2138_in & reg_q2136_in & reg_q675_in & reg_q137_in & reg_q1088_in & reg_q149_in & reg_q1327_in & reg_q1325_in & reg_q2567_in & reg_q2565_in & reg_q990_in & reg_q988_in & reg_q978_in & reg_q2260_in & reg_q2258_in & reg_q1708_in & reg_q2597_in & reg_q2310_in & reg_q2308_in & reg_q1433_in & reg_q1431_in & reg_q1137_in & reg_q1135_in & reg_q129_in & reg_q1090_in & reg_q744_in & reg_q742_in & reg_q245_in & reg_q2249_in & reg_q2247_in & reg_q1082_in & reg_q1080_in & reg_q2294_in & reg_q2292_in & reg_q135_in & reg_q133_in & reg_q111_in & reg_q1472_in & reg_q1470_in & reg_q2225_in & reg_q1732_in & reg_q1730_in & reg_q2024_in & reg_q2022_in & reg_q1548_in & reg_q1546_in & reg_q1541_in & reg_q1143_in & reg_q235_in & reg_q2028_in & reg_q305_in & reg_q1704_in & reg_q1734_in & reg_q688_in & reg_q686_in & reg_q1562_in & reg_q1560_in & reg_q2476_in & reg_q2474_in & reg_q1074_in & reg_q1072_in & reg_q1468_in & reg_q1466_in & reg_q2229_in & reg_q2227_in & reg_q2335_in & reg_q2333_in & reg_q1462_in & reg_q1460_in & reg_q335_in & reg_q333_in & reg_q2115_in & reg_q2272_in & reg_q2636_in & reg_q2634_in & reg_q2223_in & reg_q2221_in & reg_q450_in & reg_q169_in & reg_q167_in & reg_q1341_in & reg_q1339_in & reg_q2030_in & reg_q2591_in & reg_q2589_in & reg_q2373_in & reg_q2371_in & reg_q2692_in & reg_q1102_in & reg_q1317_in & reg_q1315_in & reg_q931_in & reg_q1582_in & reg_q921_in & reg_q919_in & reg_q371_in & reg_q1702_in & reg_q980_in & reg_q1002_in & reg_q125_in & reg_q290_in & reg_q288_in & reg_q2672_in & reg_q2670_in & reg_q1738_in & reg_q1736_in & reg_q1145_in & reg_q1578_in & reg_q2245_in & reg_q2243_in & reg_q1700_in & reg_q1698_in & reg_q1000_in & reg_q998_in & reg_q682_in & reg_q2286_in & reg_q2284_in & reg_q2537_in & reg_q2535_in & reg_q257_in & reg_q237_in & reg_q996_in & reg_q994_in & reg_q2170_in & reg_q2168_in & reg_q2611_in & reg_q2609_in & reg_q2217_in & reg_q2215_in & reg_q1576_in & reg_q1574_in & reg_q2119_in & reg_q2117_in & reg_q343_in & reg_q341_in & reg_q1716_in & reg_q1714_in & reg_q1189_in & reg_q1187_in & reg_q113_in & reg_q76_in & reg_q74_in & reg_q1682_in & reg_q1680_in & reg_q1423_in & reg_q1421_in & reg_q2042_in & reg_q2622_in & reg_q2620_in & reg_q1252_in & reg_q1250_in & reg_q117_in & reg_q115_in & reg_q194_in & reg_q1427_in & reg_q1425_in & reg_q1307_in & reg_q1305_in & reg_q756_in & reg_q1674_in & reg_q1531_in & reg_q2690_in & reg_q2688_in & reg_q2577_in & reg_q381_in & reg_q379_in & reg_q1678_in & reg_q1676_in & reg_q968_in & reg_q966_in & reg_q2343_in & reg_q2341_in & reg_q1337_in & reg_q127_in & reg_q2337_in & reg_q428_in & reg_q426_in & reg_q2595_in & reg_q2593_in & reg_q818_in & reg_q2613_in & reg_q123_in & reg_q121_in & reg_q2363_in & reg_q2361_in & reg_q2377_in & reg_q2375_in & reg_q2103_in & reg_q2101_in & reg_q359_in & reg_q357_in & reg_q1690_in & reg_q1688_in & reg_q418_in & reg_q198_in & reg_q196_in & reg_q700_in & reg_q369_in & reg_q367_in & reg_q1482_in & reg_q2482_in & reg_q2480_in & reg_q103_in & reg_q101_in & reg_q58_in & reg_q56_in & reg_q1108_in & reg_q1096_in & reg_q1094_in & reg_q2369_in & reg_q1248_in & reg_q1975_in & reg_q2040_in & reg_q2038_in & reg_q249_in & reg_q247_in & reg_q375_in & reg_q373_in & reg_q711_in & reg_q709_in & reg_q692_in & reg_q690_in & reg_q826_in & reg_q824_in & reg_q1580_in & reg_q1193_in & reg_q1191_in & reg_q2004_in & reg_q1357_in & reg_q1355_in & reg_q2111_in & reg_q2109_in & reg_q1335_in & reg_q1726_in & reg_q1724_in & reg_q2516_in & reg_q2514_in & reg_q1086_in & reg_q1084_in & reg_q1029_in & reg_q1027_in & reg_q2278_in & reg_q2353_in & reg_q1443_in & reg_q1441_in & reg_q1662_in & reg_q1660_in & reg_q1301_in & reg_q1529_in & reg_q1527_in & reg_q2020_in & reg_q2018_in & reg_q1480_in & reg_q1478_in & reg_q673_in & reg_q671_in & reg_q1037_in & reg_q1035_in & reg_q2276_in & reg_q2274_in & reg_q2172_in & reg_q2605_in & reg_q2603_in & reg_q1299_in & reg_q984_in & reg_q982_in & reg_q1147_in & reg_q422_in & reg_q420_in & reg_q2351_in & reg_q1670_in & reg_q1668_in & reg_q1106_in & reg_q1104_in & reg_q363_in & reg_q361_in & reg_q2302_in & reg_q1997_in & reg_q1333_in & reg_q1331_in & reg_q253_in & reg_q251_in & reg_q933_in & reg_q955_in & reg_q2579_in & reg_q848_in & reg_q828_in & reg_q1139_in;

	--coder fullgraph2
with reg_fullgraph2_sel select
reg_fullgraph2_in <=
	"0000000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001",
	"0000000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010",
	"0000000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100",
	"0000000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000",
	"0000000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000",
	"0000000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000",
	"0000000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000",
	"0000001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000",
	"0000001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
	"0000001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000",
	"0000001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000",
	"0000001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000",
	"0000001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000",
	"0000001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000",
	"0000001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000",
	"0000010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000",
	"0000010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000",
	"0000010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000",
	"0000010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000",
	"0000010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000",
	"0000010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000",
	"0000010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000",
	"0000010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000",
	"0000011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000",
	"0000011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000",
	"0000011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000",
	"0000011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000",
	"0000011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000",
	"0000011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000",
	"0000011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000",
	"0000011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000",
	"0000100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000",
	"0000100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000",
	"0000100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000",
	"0000100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000",
	"0000100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000",
	"0000100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000",
	"0000100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000",
	"0000100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000",
	"0000101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000",
	"0000101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000",
	"0000101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000",
	"0000101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000",
	"0000101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000",
	"0000101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"0000101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000",
	"0000101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000",
	"0000110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000",
	"0000110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000",
	"0000110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000",
	"0000110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000",
	"0000110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000",
	"0000110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000",
	"0000110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000",
	"0000110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000",
	"0000111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000",
	"0000111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000",
	"0000111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000",
	"0000111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000",
	"0000111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000",
	"0000111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000",
	"0000111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000",
	"0000111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000",
	"0001000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000",
	"0001000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000",
	"0001000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000",
	"0001000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000",
	"0001000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000",
	"0001000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000",
	"0001000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000",
	"0001000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0001111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0010111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0011111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0100111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0101111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0110111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0111111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1000111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1001111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1010111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011011101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011011110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011011111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011100000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011100001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011100010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011100011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011100100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011100101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011100110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011100111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011101000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011101001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011101010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011101011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011101100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011101101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011101110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011101111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011110000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011110001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011110010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011110011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011110100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011110101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011110110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011110111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011111000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011111001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011111010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011111011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011111100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011111101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011111110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1011111111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100000000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100000001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100000010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100000011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100000100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100000101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100000110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100000111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100001000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100001001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100001010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100001011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100001100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100001101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100001110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100001111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100010000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100010001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100010010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100010011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100010100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100010101" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100010110" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100010111" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100011000" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100011001" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100011010" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100011011" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"1100011100" when "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"0000000000" when others;
 --end coder

	p_reg_fullgraph2: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph2 <= reg_fullgraph2_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph2 <= reg_fullgraph2_init;
        else
          reg_fullgraph2 <= reg_fullgraph2_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph2

		reg_q1139 <= '1' when reg_fullgraph2 = "0000000001" else '0'; 
		reg_q828 <= '1' when reg_fullgraph2 = "0000000010" else '0'; 
		reg_q848 <= '1' when reg_fullgraph2 = "0000000011" else '0'; 
		reg_q2579 <= '1' when reg_fullgraph2 = "0000000100" else '0'; 
		reg_q955 <= '1' when reg_fullgraph2 = "0000000101" else '0'; 
		reg_q933 <= '1' when reg_fullgraph2 = "0000000110" else '0'; 
		reg_q251 <= '1' when reg_fullgraph2 = "0000000111" else '0'; 
		reg_q253 <= '1' when reg_fullgraph2 = "0000001000" else '0'; 
		reg_q1331 <= '1' when reg_fullgraph2 = "0000001001" else '0'; 
		reg_q1333 <= '1' when reg_fullgraph2 = "0000001010" else '0'; 
		reg_q1997 <= '1' when reg_fullgraph2 = "0000001011" else '0'; 
		reg_q2302 <= '1' when reg_fullgraph2 = "0000001100" else '0'; 
		reg_q361 <= '1' when reg_fullgraph2 = "0000001101" else '0'; 
		reg_q363 <= '1' when reg_fullgraph2 = "0000001110" else '0'; 
		reg_q1104 <= '1' when reg_fullgraph2 = "0000001111" else '0'; 
		reg_q1106 <= '1' when reg_fullgraph2 = "0000010000" else '0'; 
		reg_q1668 <= '1' when reg_fullgraph2 = "0000010001" else '0'; 
		reg_q1670 <= '1' when reg_fullgraph2 = "0000010010" else '0'; 
		reg_q2351 <= '1' when reg_fullgraph2 = "0000010011" else '0'; 
		reg_q420 <= '1' when reg_fullgraph2 = "0000010100" else '0'; 
		reg_q422 <= '1' when reg_fullgraph2 = "0000010101" else '0'; 
		reg_q1147 <= '1' when reg_fullgraph2 = "0000010110" else '0'; 
		reg_q982 <= '1' when reg_fullgraph2 = "0000010111" else '0'; 
		reg_q984 <= '1' when reg_fullgraph2 = "0000011000" else '0'; 
		reg_q1299 <= '1' when reg_fullgraph2 = "0000011001" else '0'; 
		reg_q2603 <= '1' when reg_fullgraph2 = "0000011010" else '0'; 
		reg_q2605 <= '1' when reg_fullgraph2 = "0000011011" else '0'; 
		reg_q2172 <= '1' when reg_fullgraph2 = "0000011100" else '0'; 
		reg_q2274 <= '1' when reg_fullgraph2 = "0000011101" else '0'; 
		reg_q2276 <= '1' when reg_fullgraph2 = "0000011110" else '0'; 
		reg_q1035 <= '1' when reg_fullgraph2 = "0000011111" else '0'; 
		reg_q1037 <= '1' when reg_fullgraph2 = "0000100000" else '0'; 
		reg_q671 <= '1' when reg_fullgraph2 = "0000100001" else '0'; 
		reg_q673 <= '1' when reg_fullgraph2 = "0000100010" else '0'; 
		reg_q1478 <= '1' when reg_fullgraph2 = "0000100011" else '0'; 
		reg_q1480 <= '1' when reg_fullgraph2 = "0000100100" else '0'; 
		reg_q2018 <= '1' when reg_fullgraph2 = "0000100101" else '0'; 
		reg_q2020 <= '1' when reg_fullgraph2 = "0000100110" else '0'; 
		reg_q1527 <= '1' when reg_fullgraph2 = "0000100111" else '0'; 
		reg_q1529 <= '1' when reg_fullgraph2 = "0000101000" else '0'; 
		reg_q1301 <= '1' when reg_fullgraph2 = "0000101001" else '0'; 
		reg_q1660 <= '1' when reg_fullgraph2 = "0000101010" else '0'; 
		reg_q1662 <= '1' when reg_fullgraph2 = "0000101011" else '0'; 
		reg_q1441 <= '1' when reg_fullgraph2 = "0000101100" else '0'; 
		reg_q1443 <= '1' when reg_fullgraph2 = "0000101101" else '0'; 
		reg_q2353 <= '1' when reg_fullgraph2 = "0000101110" else '0'; 
		reg_q2278 <= '1' when reg_fullgraph2 = "0000101111" else '0'; 
		reg_q1027 <= '1' when reg_fullgraph2 = "0000110000" else '0'; 
		reg_q1029 <= '1' when reg_fullgraph2 = "0000110001" else '0'; 
		reg_q1084 <= '1' when reg_fullgraph2 = "0000110010" else '0'; 
		reg_q1086 <= '1' when reg_fullgraph2 = "0000110011" else '0'; 
		reg_q2514 <= '1' when reg_fullgraph2 = "0000110100" else '0'; 
		reg_q2516 <= '1' when reg_fullgraph2 = "0000110101" else '0'; 
		reg_q1724 <= '1' when reg_fullgraph2 = "0000110110" else '0'; 
		reg_q1726 <= '1' when reg_fullgraph2 = "0000110111" else '0'; 
		reg_q1335 <= '1' when reg_fullgraph2 = "0000111000" else '0'; 
		reg_q2109 <= '1' when reg_fullgraph2 = "0000111001" else '0'; 
		reg_q2111 <= '1' when reg_fullgraph2 = "0000111010" else '0'; 
		reg_q1355 <= '1' when reg_fullgraph2 = "0000111011" else '0'; 
		reg_q1357 <= '1' when reg_fullgraph2 = "0000111100" else '0'; 
		reg_q2004 <= '1' when reg_fullgraph2 = "0000111101" else '0'; 
		reg_q1191 <= '1' when reg_fullgraph2 = "0000111110" else '0'; 
		reg_q1193 <= '1' when reg_fullgraph2 = "0000111111" else '0'; 
		reg_q1580 <= '1' when reg_fullgraph2 = "0001000000" else '0'; 
		reg_q824 <= '1' when reg_fullgraph2 = "0001000001" else '0'; 
		reg_q826 <= '1' when reg_fullgraph2 = "0001000010" else '0'; 
		reg_q690 <= '1' when reg_fullgraph2 = "0001000011" else '0'; 
		reg_q692 <= '1' when reg_fullgraph2 = "0001000100" else '0'; 
		reg_q709 <= '1' when reg_fullgraph2 = "0001000101" else '0'; 
		reg_q711 <= '1' when reg_fullgraph2 = "0001000110" else '0'; 
		reg_q373 <= '1' when reg_fullgraph2 = "0001000111" else '0'; 
		reg_q375 <= '1' when reg_fullgraph2 = "0001001000" else '0'; 
		reg_q247 <= '1' when reg_fullgraph2 = "0001001001" else '0'; 
		reg_q249 <= '1' when reg_fullgraph2 = "0001001010" else '0'; 
		reg_q2038 <= '1' when reg_fullgraph2 = "0001001011" else '0'; 
		reg_q2040 <= '1' when reg_fullgraph2 = "0001001100" else '0'; 
		reg_q1975 <= '1' when reg_fullgraph2 = "0001001101" else '0'; 
		reg_q1248 <= '1' when reg_fullgraph2 = "0001001110" else '0'; 
		reg_q2369 <= '1' when reg_fullgraph2 = "0001001111" else '0'; 
		reg_q1094 <= '1' when reg_fullgraph2 = "0001010000" else '0'; 
		reg_q1096 <= '1' when reg_fullgraph2 = "0001010001" else '0'; 
		reg_q1108 <= '1' when reg_fullgraph2 = "0001010010" else '0'; 
		reg_q56 <= '1' when reg_fullgraph2 = "0001010011" else '0'; 
		reg_q58 <= '1' when reg_fullgraph2 = "0001010100" else '0'; 
		reg_q101 <= '1' when reg_fullgraph2 = "0001010101" else '0'; 
		reg_q103 <= '1' when reg_fullgraph2 = "0001010110" else '0'; 
		reg_q2480 <= '1' when reg_fullgraph2 = "0001010111" else '0'; 
		reg_q2482 <= '1' when reg_fullgraph2 = "0001011000" else '0'; 
		reg_q1482 <= '1' when reg_fullgraph2 = "0001011001" else '0'; 
		reg_q367 <= '1' when reg_fullgraph2 = "0001011010" else '0'; 
		reg_q369 <= '1' when reg_fullgraph2 = "0001011011" else '0'; 
		reg_q700 <= '1' when reg_fullgraph2 = "0001011100" else '0'; 
		reg_q196 <= '1' when reg_fullgraph2 = "0001011101" else '0'; 
		reg_q198 <= '1' when reg_fullgraph2 = "0001011110" else '0'; 
		reg_q418 <= '1' when reg_fullgraph2 = "0001011111" else '0'; 
		reg_q1688 <= '1' when reg_fullgraph2 = "0001100000" else '0'; 
		reg_q1690 <= '1' when reg_fullgraph2 = "0001100001" else '0'; 
		reg_q357 <= '1' when reg_fullgraph2 = "0001100010" else '0'; 
		reg_q359 <= '1' when reg_fullgraph2 = "0001100011" else '0'; 
		reg_q2101 <= '1' when reg_fullgraph2 = "0001100100" else '0'; 
		reg_q2103 <= '1' when reg_fullgraph2 = "0001100101" else '0'; 
		reg_q2375 <= '1' when reg_fullgraph2 = "0001100110" else '0'; 
		reg_q2377 <= '1' when reg_fullgraph2 = "0001100111" else '0'; 
		reg_q2361 <= '1' when reg_fullgraph2 = "0001101000" else '0'; 
		reg_q2363 <= '1' when reg_fullgraph2 = "0001101001" else '0'; 
		reg_q121 <= '1' when reg_fullgraph2 = "0001101010" else '0'; 
		reg_q123 <= '1' when reg_fullgraph2 = "0001101011" else '0'; 
		reg_q2613 <= '1' when reg_fullgraph2 = "0001101100" else '0'; 
		reg_q818 <= '1' when reg_fullgraph2 = "0001101101" else '0'; 
		reg_q2593 <= '1' when reg_fullgraph2 = "0001101110" else '0'; 
		reg_q2595 <= '1' when reg_fullgraph2 = "0001101111" else '0'; 
		reg_q426 <= '1' when reg_fullgraph2 = "0001110000" else '0'; 
		reg_q428 <= '1' when reg_fullgraph2 = "0001110001" else '0'; 
		reg_q2337 <= '1' when reg_fullgraph2 = "0001110010" else '0'; 
		reg_q127 <= '1' when reg_fullgraph2 = "0001110011" else '0'; 
		reg_q1337 <= '1' when reg_fullgraph2 = "0001110100" else '0'; 
		reg_q2341 <= '1' when reg_fullgraph2 = "0001110101" else '0'; 
		reg_q2343 <= '1' when reg_fullgraph2 = "0001110110" else '0'; 
		reg_q966 <= '1' when reg_fullgraph2 = "0001110111" else '0'; 
		reg_q968 <= '1' when reg_fullgraph2 = "0001111000" else '0'; 
		reg_q1676 <= '1' when reg_fullgraph2 = "0001111001" else '0'; 
		reg_q1678 <= '1' when reg_fullgraph2 = "0001111010" else '0'; 
		reg_q379 <= '1' when reg_fullgraph2 = "0001111011" else '0'; 
		reg_q381 <= '1' when reg_fullgraph2 = "0001111100" else '0'; 
		reg_q2577 <= '1' when reg_fullgraph2 = "0001111101" else '0'; 
		reg_q2688 <= '1' when reg_fullgraph2 = "0001111110" else '0'; 
		reg_q2690 <= '1' when reg_fullgraph2 = "0001111111" else '0'; 
		reg_q1531 <= '1' when reg_fullgraph2 = "0010000000" else '0'; 
		reg_q1674 <= '1' when reg_fullgraph2 = "0010000001" else '0'; 
		reg_q756 <= '1' when reg_fullgraph2 = "0010000010" else '0'; 
		reg_q1305 <= '1' when reg_fullgraph2 = "0010000011" else '0'; 
		reg_q1307 <= '1' when reg_fullgraph2 = "0010000100" else '0'; 
		reg_q1425 <= '1' when reg_fullgraph2 = "0010000101" else '0'; 
		reg_q1427 <= '1' when reg_fullgraph2 = "0010000110" else '0'; 
		reg_q194 <= '1' when reg_fullgraph2 = "0010000111" else '0'; 
		reg_q115 <= '1' when reg_fullgraph2 = "0010001000" else '0'; 
		reg_q117 <= '1' when reg_fullgraph2 = "0010001001" else '0'; 
		reg_q1250 <= '1' when reg_fullgraph2 = "0010001010" else '0'; 
		reg_q1252 <= '1' when reg_fullgraph2 = "0010001011" else '0'; 
		reg_q2620 <= '1' when reg_fullgraph2 = "0010001100" else '0'; 
		reg_q2622 <= '1' when reg_fullgraph2 = "0010001101" else '0'; 
		reg_q2042 <= '1' when reg_fullgraph2 = "0010001110" else '0'; 
		reg_q1421 <= '1' when reg_fullgraph2 = "0010001111" else '0'; 
		reg_q1423 <= '1' when reg_fullgraph2 = "0010010000" else '0'; 
		reg_q1680 <= '1' when reg_fullgraph2 = "0010010001" else '0'; 
		reg_q1682 <= '1' when reg_fullgraph2 = "0010010010" else '0'; 
		reg_q74 <= '1' when reg_fullgraph2 = "0010010011" else '0'; 
		reg_q76 <= '1' when reg_fullgraph2 = "0010010100" else '0'; 
		reg_q113 <= '1' when reg_fullgraph2 = "0010010101" else '0'; 
		reg_q1187 <= '1' when reg_fullgraph2 = "0010010110" else '0'; 
		reg_q1189 <= '1' when reg_fullgraph2 = "0010010111" else '0'; 
		reg_q1714 <= '1' when reg_fullgraph2 = "0010011000" else '0'; 
		reg_q1716 <= '1' when reg_fullgraph2 = "0010011001" else '0'; 
		reg_q341 <= '1' when reg_fullgraph2 = "0010011010" else '0'; 
		reg_q343 <= '1' when reg_fullgraph2 = "0010011011" else '0'; 
		reg_q2117 <= '1' when reg_fullgraph2 = "0010011100" else '0'; 
		reg_q2119 <= '1' when reg_fullgraph2 = "0010011101" else '0'; 
		reg_q1574 <= '1' when reg_fullgraph2 = "0010011110" else '0'; 
		reg_q1576 <= '1' when reg_fullgraph2 = "0010011111" else '0'; 
		reg_q2215 <= '1' when reg_fullgraph2 = "0010100000" else '0'; 
		reg_q2217 <= '1' when reg_fullgraph2 = "0010100001" else '0'; 
		reg_q2609 <= '1' when reg_fullgraph2 = "0010100010" else '0'; 
		reg_q2611 <= '1' when reg_fullgraph2 = "0010100011" else '0'; 
		reg_q2168 <= '1' when reg_fullgraph2 = "0010100100" else '0'; 
		reg_q2170 <= '1' when reg_fullgraph2 = "0010100101" else '0'; 
		reg_q994 <= '1' when reg_fullgraph2 = "0010100110" else '0'; 
		reg_q996 <= '1' when reg_fullgraph2 = "0010100111" else '0'; 
		reg_q237 <= '1' when reg_fullgraph2 = "0010101000" else '0'; 
		reg_q257 <= '1' when reg_fullgraph2 = "0010101001" else '0'; 
		reg_q2535 <= '1' when reg_fullgraph2 = "0010101010" else '0'; 
		reg_q2537 <= '1' when reg_fullgraph2 = "0010101011" else '0'; 
		reg_q2284 <= '1' when reg_fullgraph2 = "0010101100" else '0'; 
		reg_q2286 <= '1' when reg_fullgraph2 = "0010101101" else '0'; 
		reg_q682 <= '1' when reg_fullgraph2 = "0010101110" else '0'; 
		reg_q998 <= '1' when reg_fullgraph2 = "0010101111" else '0'; 
		reg_q1000 <= '1' when reg_fullgraph2 = "0010110000" else '0'; 
		reg_q1698 <= '1' when reg_fullgraph2 = "0010110001" else '0'; 
		reg_q1700 <= '1' when reg_fullgraph2 = "0010110010" else '0'; 
		reg_q2243 <= '1' when reg_fullgraph2 = "0010110011" else '0'; 
		reg_q2245 <= '1' when reg_fullgraph2 = "0010110100" else '0'; 
		reg_q1578 <= '1' when reg_fullgraph2 = "0010110101" else '0'; 
		reg_q1145 <= '1' when reg_fullgraph2 = "0010110110" else '0'; 
		reg_q1736 <= '1' when reg_fullgraph2 = "0010110111" else '0'; 
		reg_q1738 <= '1' when reg_fullgraph2 = "0010111000" else '0'; 
		reg_q2670 <= '1' when reg_fullgraph2 = "0010111001" else '0'; 
		reg_q2672 <= '1' when reg_fullgraph2 = "0010111010" else '0'; 
		reg_q288 <= '1' when reg_fullgraph2 = "0010111011" else '0'; 
		reg_q290 <= '1' when reg_fullgraph2 = "0010111100" else '0'; 
		reg_q125 <= '1' when reg_fullgraph2 = "0010111101" else '0'; 
		reg_q1002 <= '1' when reg_fullgraph2 = "0010111110" else '0'; 
		reg_q980 <= '1' when reg_fullgraph2 = "0010111111" else '0'; 
		reg_q1702 <= '1' when reg_fullgraph2 = "0011000000" else '0'; 
		reg_q371 <= '1' when reg_fullgraph2 = "0011000001" else '0'; 
		reg_q919 <= '1' when reg_fullgraph2 = "0011000010" else '0'; 
		reg_q921 <= '1' when reg_fullgraph2 = "0011000011" else '0'; 
		reg_q1582 <= '1' when reg_fullgraph2 = "0011000100" else '0'; 
		reg_q931 <= '1' when reg_fullgraph2 = "0011000101" else '0'; 
		reg_q1315 <= '1' when reg_fullgraph2 = "0011000110" else '0'; 
		reg_q1317 <= '1' when reg_fullgraph2 = "0011000111" else '0'; 
		reg_q1102 <= '1' when reg_fullgraph2 = "0011001000" else '0'; 
		reg_q2692 <= '1' when reg_fullgraph2 = "0011001001" else '0'; 
		reg_q2371 <= '1' when reg_fullgraph2 = "0011001010" else '0'; 
		reg_q2373 <= '1' when reg_fullgraph2 = "0011001011" else '0'; 
		reg_q2589 <= '1' when reg_fullgraph2 = "0011001100" else '0'; 
		reg_q2591 <= '1' when reg_fullgraph2 = "0011001101" else '0'; 
		reg_q2030 <= '1' when reg_fullgraph2 = "0011001110" else '0'; 
		reg_q1339 <= '1' when reg_fullgraph2 = "0011001111" else '0'; 
		reg_q1341 <= '1' when reg_fullgraph2 = "0011010000" else '0'; 
		reg_q167 <= '1' when reg_fullgraph2 = "0011010001" else '0'; 
		reg_q169 <= '1' when reg_fullgraph2 = "0011010010" else '0'; 
		reg_q450 <= '1' when reg_fullgraph2 = "0011010011" else '0'; 
		reg_q2221 <= '1' when reg_fullgraph2 = "0011010100" else '0'; 
		reg_q2223 <= '1' when reg_fullgraph2 = "0011010101" else '0'; 
		reg_q2634 <= '1' when reg_fullgraph2 = "0011010110" else '0'; 
		reg_q2636 <= '1' when reg_fullgraph2 = "0011010111" else '0'; 
		reg_q2272 <= '1' when reg_fullgraph2 = "0011011000" else '0'; 
		reg_q2115 <= '1' when reg_fullgraph2 = "0011011001" else '0'; 
		reg_q333 <= '1' when reg_fullgraph2 = "0011011010" else '0'; 
		reg_q335 <= '1' when reg_fullgraph2 = "0011011011" else '0'; 
		reg_q1460 <= '1' when reg_fullgraph2 = "0011011100" else '0'; 
		reg_q1462 <= '1' when reg_fullgraph2 = "0011011101" else '0'; 
		reg_q2333 <= '1' when reg_fullgraph2 = "0011011110" else '0'; 
		reg_q2335 <= '1' when reg_fullgraph2 = "0011011111" else '0'; 
		reg_q2227 <= '1' when reg_fullgraph2 = "0011100000" else '0'; 
		reg_q2229 <= '1' when reg_fullgraph2 = "0011100001" else '0'; 
		reg_q1466 <= '1' when reg_fullgraph2 = "0011100010" else '0'; 
		reg_q1468 <= '1' when reg_fullgraph2 = "0011100011" else '0'; 
		reg_q1072 <= '1' when reg_fullgraph2 = "0011100100" else '0'; 
		reg_q1074 <= '1' when reg_fullgraph2 = "0011100101" else '0'; 
		reg_q2474 <= '1' when reg_fullgraph2 = "0011100110" else '0'; 
		reg_q2476 <= '1' when reg_fullgraph2 = "0011100111" else '0'; 
		reg_q1560 <= '1' when reg_fullgraph2 = "0011101000" else '0'; 
		reg_q1562 <= '1' when reg_fullgraph2 = "0011101001" else '0'; 
		reg_q686 <= '1' when reg_fullgraph2 = "0011101010" else '0'; 
		reg_q688 <= '1' when reg_fullgraph2 = "0011101011" else '0'; 
		reg_q1734 <= '1' when reg_fullgraph2 = "0011101100" else '0'; 
		reg_q1704 <= '1' when reg_fullgraph2 = "0011101101" else '0'; 
		reg_q305 <= '1' when reg_fullgraph2 = "0011101110" else '0'; 
		reg_q2028 <= '1' when reg_fullgraph2 = "0011101111" else '0'; 
		reg_q235 <= '1' when reg_fullgraph2 = "0011110000" else '0'; 
		reg_q1143 <= '1' when reg_fullgraph2 = "0011110001" else '0'; 
		reg_q1541 <= '1' when reg_fullgraph2 = "0011110010" else '0'; 
		reg_q1546 <= '1' when reg_fullgraph2 = "0011110011" else '0'; 
		reg_q1548 <= '1' when reg_fullgraph2 = "0011110100" else '0'; 
		reg_q2022 <= '1' when reg_fullgraph2 = "0011110101" else '0'; 
		reg_q2024 <= '1' when reg_fullgraph2 = "0011110110" else '0'; 
		reg_q1730 <= '1' when reg_fullgraph2 = "0011110111" else '0'; 
		reg_q1732 <= '1' when reg_fullgraph2 = "0011111000" else '0'; 
		reg_q2225 <= '1' when reg_fullgraph2 = "0011111001" else '0'; 
		reg_q1470 <= '1' when reg_fullgraph2 = "0011111010" else '0'; 
		reg_q1472 <= '1' when reg_fullgraph2 = "0011111011" else '0'; 
		reg_q111 <= '1' when reg_fullgraph2 = "0011111100" else '0'; 
		reg_q133 <= '1' when reg_fullgraph2 = "0011111101" else '0'; 
		reg_q135 <= '1' when reg_fullgraph2 = "0011111110" else '0'; 
		reg_q2292 <= '1' when reg_fullgraph2 = "0011111111" else '0'; 
		reg_q2294 <= '1' when reg_fullgraph2 = "0100000000" else '0'; 
		reg_q1080 <= '1' when reg_fullgraph2 = "0100000001" else '0'; 
		reg_q1082 <= '1' when reg_fullgraph2 = "0100000010" else '0'; 
		reg_q2247 <= '1' when reg_fullgraph2 = "0100000011" else '0'; 
		reg_q2249 <= '1' when reg_fullgraph2 = "0100000100" else '0'; 
		reg_q245 <= '1' when reg_fullgraph2 = "0100000101" else '0'; 
		reg_q742 <= '1' when reg_fullgraph2 = "0100000110" else '0'; 
		reg_q744 <= '1' when reg_fullgraph2 = "0100000111" else '0'; 
		reg_q1090 <= '1' when reg_fullgraph2 = "0100001000" else '0'; 
		reg_q129 <= '1' when reg_fullgraph2 = "0100001001" else '0'; 
		reg_q1135 <= '1' when reg_fullgraph2 = "0100001010" else '0'; 
		reg_q1137 <= '1' when reg_fullgraph2 = "0100001011" else '0'; 
		reg_q1431 <= '1' when reg_fullgraph2 = "0100001100" else '0'; 
		reg_q1433 <= '1' when reg_fullgraph2 = "0100001101" else '0'; 
		reg_q2308 <= '1' when reg_fullgraph2 = "0100001110" else '0'; 
		reg_q2310 <= '1' when reg_fullgraph2 = "0100001111" else '0'; 
		reg_q2597 <= '1' when reg_fullgraph2 = "0100010000" else '0'; 
		reg_q1708 <= '1' when reg_fullgraph2 = "0100010001" else '0'; 
		reg_q2258 <= '1' when reg_fullgraph2 = "0100010010" else '0'; 
		reg_q2260 <= '1' when reg_fullgraph2 = "0100010011" else '0'; 
		reg_q978 <= '1' when reg_fullgraph2 = "0100010100" else '0'; 
		reg_q988 <= '1' when reg_fullgraph2 = "0100010101" else '0'; 
		reg_q990 <= '1' when reg_fullgraph2 = "0100010110" else '0'; 
		reg_q2565 <= '1' when reg_fullgraph2 = "0100010111" else '0'; 
		reg_q2567 <= '1' when reg_fullgraph2 = "0100011000" else '0'; 
		reg_q1325 <= '1' when reg_fullgraph2 = "0100011001" else '0'; 
		reg_q1327 <= '1' when reg_fullgraph2 = "0100011010" else '0'; 
		reg_q149 <= '1' when reg_fullgraph2 = "0100011011" else '0'; 
		reg_q1088 <= '1' when reg_fullgraph2 = "0100011100" else '0'; 
		reg_q137 <= '1' when reg_fullgraph2 = "0100011101" else '0'; 
		reg_q675 <= '1' when reg_fullgraph2 = "0100011110" else '0'; 
		reg_q2136 <= '1' when reg_fullgraph2 = "0100011111" else '0'; 
		reg_q2138 <= '1' when reg_fullgraph2 = "0100100000" else '0'; 
		reg_q119 <= '1' when reg_fullgraph2 = "0100100001" else '0'; 
		reg_q255 <= '1' when reg_fullgraph2 = "0100100010" else '0'; 
		reg_q915 <= '1' when reg_fullgraph2 = "0100100011" else '0'; 
		reg_q1008 <= '1' when reg_fullgraph2 = "0100100100" else '0'; 
		reg_q1010 <= '1' when reg_fullgraph2 = "0100100101" else '0'; 
		reg_q1672 <= '1' when reg_fullgraph2 = "0100100110" else '0'; 
		reg_q2642 <= '1' when reg_fullgraph2 = "0100100111" else '0'; 
		reg_q2644 <= '1' when reg_fullgraph2 = "0100101000" else '0'; 
		reg_q2599 <= '1' when reg_fullgraph2 = "0100101001" else '0'; 
		reg_q2601 <= '1' when reg_fullgraph2 = "0100101010" else '0'; 
		reg_q1637 <= '1' when reg_fullgraph2 = "0100101011" else '0'; 
		reg_q1639 <= '1' when reg_fullgraph2 = "0100101100" else '0'; 
		reg_q107 <= '1' when reg_fullgraph2 = "0100101101" else '0'; 
		reg_q109 <= '1' when reg_fullgraph2 = "0100101110" else '0'; 
		reg_q783 <= '1' when reg_fullgraph2 = "0100101111" else '0'; 
		reg_q785 <= '1' when reg_fullgraph2 = "0100110000" else '0'; 
		reg_q1092 <= '1' when reg_fullgraph2 = "0100110001" else '0'; 
		reg_q1347 <= '1' when reg_fullgraph2 = "0100110010" else '0'; 
		reg_q1349 <= '1' when reg_fullgraph2 = "0100110011" else '0'; 
		reg_q1115 <= '1' when reg_fullgraph2 = "0100110100" else '0'; 
		reg_q1117 <= '1' when reg_fullgraph2 = "0100110101" else '0'; 
		reg_q448 <= '1' when reg_fullgraph2 = "0100110110" else '0'; 
		reg_q192 <= '1' when reg_fullgraph2 = "0100110111" else '0'; 
		reg_q395 <= '1' when reg_fullgraph2 = "0100111000" else '0'; 
		reg_q397 <= '1' when reg_fullgraph2 = "0100111001" else '0'; 
		reg_q84 <= '1' when reg_fullgraph2 = "0100111010" else '0'; 
		reg_q86 <= '1' when reg_fullgraph2 = "0100111011" else '0'; 
		reg_q365 <= '1' when reg_fullgraph2 = "0100111100" else '0'; 
		reg_q698 <= '1' when reg_fullgraph2 = "0100111101" else '0'; 
		reg_q1437 <= '1' when reg_fullgraph2 = "0100111110" else '0'; 
		reg_q964 <= '1' when reg_fullgraph2 = "0100111111" else '0'; 
		reg_q748 <= '1' when reg_fullgraph2 = "0101000000" else '0'; 
		reg_q750 <= '1' when reg_fullgraph2 = "0101000001" else '0'; 
		reg_q1435 <= '1' when reg_fullgraph2 = "0101000010" else '0'; 
		reg_q1692 <= '1' when reg_fullgraph2 = "0101000011" else '0'; 
		reg_q1262 <= '1' when reg_fullgraph2 = "0101000100" else '0'; 
		reg_q1264 <= '1' when reg_fullgraph2 = "0101000101" else '0'; 
		reg_q2686 <= '1' when reg_fullgraph2 = "0101000110" else '0'; 
		reg_q2349 <= '1' when reg_fullgraph2 = "0101000111" else '0'; 
		reg_q1023 <= '1' when reg_fullgraph2 = "0101001000" else '0'; 
		reg_q1025 <= '1' when reg_fullgraph2 = "0101001001" else '0'; 
		reg_q1133 <= '1' when reg_fullgraph2 = "0101001010" else '0'; 
		reg_q2575 <= '1' when reg_fullgraph2 = "0101001011" else '0'; 
		reg_q1272 <= '1' when reg_fullgraph2 = "0101001100" else '0'; 
		reg_q1274 <= '1' when reg_fullgraph2 = "0101001101" else '0'; 
		reg_q1504 <= '1' when reg_fullgraph2 = "0101001110" else '0'; 
		reg_q1506 <= '1' when reg_fullgraph2 = "0101001111" else '0'; 
		reg_q2497 <= '1' when reg_fullgraph2 = "0101010000" else '0'; 
		reg_q2499 <= '1' when reg_fullgraph2 = "0101010001" else '0'; 
		reg_q923 <= '1' when reg_fullgraph2 = "0101010010" else '0'; 
		reg_q925 <= '1' when reg_fullgraph2 = "0101010011" else '0'; 
		reg_q1635 <= '1' when reg_fullgraph2 = "0101010100" else '0'; 
		reg_q323 <= '1' when reg_fullgraph2 = "0101010101" else '0'; 
		reg_q325 <= '1' when reg_fullgraph2 = "0101010110" else '0'; 
		reg_q292 <= '1' when reg_fullgraph2 = "0101010111" else '0'; 
		reg_q294 <= '1' when reg_fullgraph2 = "0101011000" else '0'; 
		reg_q1664 <= '1' when reg_fullgraph2 = "0101011001" else '0'; 
		reg_q1666 <= '1' when reg_fullgraph2 = "0101011010" else '0'; 
		reg_q377 <= '1' when reg_fullgraph2 = "0101011011" else '0'; 
		reg_q1652 <= '1' when reg_fullgraph2 = "0101011100" else '0'; 
		reg_q1728 <= '1' when reg_fullgraph2 = "0101011101" else '0'; 
		reg_q1151 <= '1' when reg_fullgraph2 = "0101011110" else '0'; 
		reg_q1153 <= '1' when reg_fullgraph2 = "0101011111" else '0'; 
		reg_q1971 <= '1' when reg_fullgraph2 = "0101100000" else '0'; 
		reg_q1973 <= '1' when reg_fullgraph2 = "0101100001" else '0'; 
		reg_q1552 <= '1' when reg_fullgraph2 = "0101100010" else '0'; 
		reg_q1179 <= '1' when reg_fullgraph2 = "0101100011" else '0'; 
		reg_q1181 <= '1' when reg_fullgraph2 = "0101100100" else '0'; 
		reg_q913 <= '1' when reg_fullgraph2 = "0101100101" else '0'; 
		reg_q2304 <= '1' when reg_fullgraph2 = "0101100110" else '0'; 
		reg_q2306 <= '1' when reg_fullgraph2 = "0101100111" else '0'; 
		reg_q1319 <= '1' when reg_fullgraph2 = "0101101000" else '0'; 
		reg_q986 <= '1' when reg_fullgraph2 = "0101101001" else '0'; 
		reg_q82 <= '1' when reg_fullgraph2 = "0101101010" else '0'; 
		reg_q280 <= '1' when reg_fullgraph2 = "0101101011" else '0'; 
		reg_q282 <= '1' when reg_fullgraph2 = "0101101100" else '0'; 
		reg_q2158 <= '1' when reg_fullgraph2 = "0101101101" else '0'; 
		reg_q2160 <= '1' when reg_fullgraph2 = "0101101110" else '0'; 
		reg_q1484 <= '1' when reg_fullgraph2 = "0101101111" else '0'; 
		reg_q2674 <= '1' when reg_fullgraph2 = "0101110000" else '0'; 
		reg_q2676 <= '1' when reg_fullgraph2 = "0101110001" else '0'; 
		reg_q440 <= '1' when reg_fullgraph2 = "0101110010" else '0'; 
		reg_q442 <= '1' when reg_fullgraph2 = "0101110011" else '0'; 
		reg_q403 <= '1' when reg_fullgraph2 = "0101110100" else '0'; 
		reg_q405 <= '1' when reg_fullgraph2 = "0101110101" else '0'; 
		reg_q1246 <= '1' when reg_fullgraph2 = "0101110110" else '0'; 
		reg_q752 <= '1' when reg_fullgraph2 = "0101110111" else '0'; 
		reg_q1445 <= '1' when reg_fullgraph2 = "0101111000" else '0'; 
		reg_q2288 <= '1' when reg_fullgraph2 = "0101111001" else '0'; 
		reg_q1490 <= '1' when reg_fullgraph2 = "0101111010" else '0'; 
		reg_q2130 <= '1' when reg_fullgraph2 = "0101111011" else '0'; 
		reg_q2280 <= '1' when reg_fullgraph2 = "0101111100" else '0'; 
		reg_q2282 <= '1' when reg_fullgraph2 = "0101111101" else '0'; 
		reg_q1535 <= '1' when reg_fullgraph2 = "0101111110" else '0'; 
		reg_q1537 <= '1' when reg_fullgraph2 = "0101111111" else '0'; 
		reg_q313 <= '1' when reg_fullgraph2 = "0110000000" else '0'; 
		reg_q315 <= '1' when reg_fullgraph2 = "0110000001" else '0'; 
		reg_q1556 <= '1' when reg_fullgraph2 = "0110000010" else '0'; 
		reg_q1558 <= '1' when reg_fullgraph2 = "0110000011" else '0'; 
		reg_q1439 <= '1' when reg_fullgraph2 = "0110000100" else '0'; 
		reg_q2357 <= '1' when reg_fullgraph2 = "0110000101" else '0'; 
		reg_q2359 <= '1' when reg_fullgraph2 = "0110000110" else '0'; 
		reg_q2105 <= '1' when reg_fullgraph2 = "0110000111" else '0'; 
		reg_q2640 <= '1' when reg_fullgraph2 = "0110001000" else '0'; 
		reg_q241 <= '1' when reg_fullgraph2 = "0110001001" else '0'; 
		reg_q1313 <= '1' when reg_fullgraph2 = "0110001010" else '0'; 
		reg_q1256 <= '1' when reg_fullgraph2 = "0110001011" else '0'; 
		reg_q1033 <= '1' when reg_fullgraph2 = "0110001100" else '0'; 
		reg_q2624 <= '1' when reg_fullgraph2 = "0110001101" else '0'; 
		reg_q974 <= '1' when reg_fullgraph2 = "0110001110" else '0'; 
		reg_q976 <= '1' when reg_fullgraph2 = "0110001111" else '0'; 
		reg_q992 <= '1' when reg_fullgraph2 = "0110010000" else '0'; 
		reg_q298 <= '1' when reg_fullgraph2 = "0110010001" else '0'; 
		reg_q300 <= '1' when reg_fullgraph2 = "0110010010" else '0'; 
		reg_q696 <= '1' when reg_fullgraph2 = "0110010011" else '0'; 
		reg_q1539 <= '1' when reg_fullgraph2 = "0110010100" else '0'; 
		reg_q161 <= '1' when reg_fullgraph2 = "0110010101" else '0'; 
		reg_q163 <= '1' when reg_fullgraph2 = "0110010110" else '0'; 
		reg_q2547 <= '1' when reg_fullgraph2 = "0110010111" else '0'; 
		reg_q2549 <= '1' when reg_fullgraph2 = "0110011000" else '0'; 
		reg_q1070 <= '1' when reg_fullgraph2 = "0110011001" else '0'; 
		reg_q438 <= '1' when reg_fullgraph2 = "0110011010" else '0'; 
		reg_q1710 <= '1' when reg_fullgraph2 = "0110011011" else '0'; 
		reg_q1712 <= '1' when reg_fullgraph2 = "0110011100" else '0'; 
		reg_q407 <= '1' when reg_fullgraph2 = "0110011101" else '0'; 
		reg_q409 <= '1' when reg_fullgraph2 = "0110011110" else '0'; 
		reg_q2470 <= '1' when reg_fullgraph2 = "0110011111" else '0'; 
		reg_q2472 <= '1' when reg_fullgraph2 = "0110100000" else '0'; 
		reg_q200 <= '1' when reg_fullgraph2 = "0110100001" else '0'; 
		reg_q88 <= '1' when reg_fullgraph2 = "0110100010" else '0'; 
		reg_q1230 <= '1' when reg_fullgraph2 = "0110100011" else '0'; 
		reg_q1232 <= '1' when reg_fullgraph2 = "0110100100" else '0'; 
		reg_q2646 <= '1' when reg_fullgraph2 = "0110100101" else '0'; 
		reg_q2648 <= '1' when reg_fullgraph2 = "0110100110" else '0'; 
		reg_q1254 <= '1' when reg_fullgraph2 = "0110100111" else '0'; 
		reg_q1474 <= '1' when reg_fullgraph2 = "0110101000" else '0'; 
		reg_q66 <= '1' when reg_fullgraph2 = "0110101001" else '0'; 
		reg_q68 <= '1' when reg_fullgraph2 = "0110101010" else '0'; 
		reg_q2300 <= '1' when reg_fullgraph2 = "0110101011" else '0'; 
		reg_q2268 <= '1' when reg_fullgraph2 = "0110101100" else '0'; 
		reg_q2270 <= '1' when reg_fullgraph2 = "0110101101" else '0'; 
		reg_q2032 <= '1' when reg_fullgraph2 = "0110101110" else '0'; 
		reg_q2034 <= '1' when reg_fullgraph2 = "0110101111" else '0'; 
		reg_q430 <= '1' when reg_fullgraph2 = "0110110000" else '0'; 
		reg_q766 <= '1' when reg_fullgraph2 = "0110110001" else '0'; 
		reg_q768 <= '1' when reg_fullgraph2 = "0110110010" else '0'; 
		reg_q2662 <= '1' when reg_fullgraph2 = "0110110011" else '0'; 
		reg_q2664 <= '1' when reg_fullgraph2 = "0110110100" else '0'; 
		reg_q139 <= '1' when reg_fullgraph2 = "0110110101" else '0'; 
		reg_q1141 <= '1' when reg_fullgraph2 = "0110110110" else '0'; 
		reg_q2010 <= '1' when reg_fullgraph2 = "0110110111" else '0'; 
		reg_q2012 <= '1' when reg_fullgraph2 = "0110111000" else '0'; 
		reg_q1068 <= '1' when reg_fullgraph2 = "0110111001" else '0'; 
		reg_q2557 <= '1' when reg_fullgraph2 = "0110111010" else '0'; 
		reg_q2559 <= '1' when reg_fullgraph2 = "0110111011" else '0'; 
		reg_q1617 <= '1' when reg_fullgraph2 = "0110111100" else '0'; 
		reg_q1619 <= '1' when reg_fullgraph2 = "0110111101" else '0'; 
		reg_q1258 <= '1' when reg_fullgraph2 = "0110111110" else '0'; 
		reg_q1260 <= '1' when reg_fullgraph2 = "0110111111" else '0'; 
		reg_q734 <= '1' when reg_fullgraph2 = "0111000000" else '0'; 
		reg_q1447 <= '1' when reg_fullgraph2 = "0111000001" else '0'; 
		reg_q2014 <= '1' when reg_fullgraph2 = "0111000010" else '0'; 
		reg_q2502 <= '1' when reg_fullgraph2 = "0111000011" else '0'; 
		reg_q2296 <= '1' when reg_fullgraph2 = "0111000100" else '0'; 
		reg_q2298 <= '1' when reg_fullgraph2 = "0111000101" else '0'; 
		reg_q1159 <= '1' when reg_fullgraph2 = "0111000110" else '0'; 
		reg_q444 <= '1' when reg_fullgraph2 = "0111000111" else '0'; 
		reg_q446 <= '1' when reg_fullgraph2 = "0111001000" else '0'; 
		reg_q1183 <= '1' when reg_fullgraph2 = "0111001001" else '0'; 
		reg_q1185 <= '1' when reg_fullgraph2 = "0111001010" else '0'; 
		reg_q962 <= '1' when reg_fullgraph2 = "0111001011" else '0'; 
		reg_q2573 <= '1' when reg_fullgraph2 = "0111001100" else '0'; 
		reg_q1123 <= '1' when reg_fullgraph2 = "0111001101" else '0'; 
		reg_q1125 <= '1' when reg_fullgraph2 = "0111001110" else '0'; 
		reg_q1613 <= '1' when reg_fullgraph2 = "0111001111" else '0'; 
		reg_q2339 <= '1' when reg_fullgraph2 = "0111010000" else '0'; 
		reg_q667 <= '1' when reg_fullgraph2 = "0111010001" else '0'; 
		reg_q60 <= '1' when reg_fullgraph2 = "0111010010" else '0'; 
		reg_q399 <= '1' when reg_fullgraph2 = "0111010011" else '0'; 
		reg_q2650 <= '1' when reg_fullgraph2 = "0111010100" else '0'; 
		reg_q1076 <= '1' when reg_fullgraph2 = "0111010101" else '0'; 
		reg_q1078 <= '1' when reg_fullgraph2 = "0111010110" else '0'; 
		reg_q284 <= '1' when reg_fullgraph2 = "0111010111" else '0'; 
		reg_q2095 <= '1' when reg_fullgraph2 = "0111011000" else '0'; 
		reg_q171 <= '1' when reg_fullgraph2 = "0111011001" else '0'; 
		reg_q239 <= '1' when reg_fullgraph2 = "0111011010" else '0'; 
		reg_q278 <= '1' when reg_fullgraph2 = "0111011011" else '0'; 
		reg_q105 <= '1' when reg_fullgraph2 = "0111011100" else '0'; 
		reg_q2148 <= '1' when reg_fullgraph2 = "0111011101" else '0'; 
		reg_q1343 <= '1' when reg_fullgraph2 = "0111011110" else '0'; 
		reg_q1625 <= '1' when reg_fullgraph2 = "0111011111" else '0'; 
		reg_q1627 <= '1' when reg_fullgraph2 = "0111100000" else '0'; 
		reg_q349 <= '1' when reg_fullgraph2 = "0111100001" else '0'; 
		reg_q351 <= '1' when reg_fullgraph2 = "0111100010" else '0'; 
		reg_q1648 <= '1' when reg_fullgraph2 = "0111100011" else '0'; 
		reg_q307 <= '1' when reg_fullgraph2 = "0111100100" else '0'; 
		reg_q2290 <= '1' when reg_fullgraph2 = "0111100101" else '0'; 
		reg_q1533 <= '1' when reg_fullgraph2 = "0111100110" else '0'; 
		reg_q2237 <= '1' when reg_fullgraph2 = "0111100111" else '0'; 
		reg_q2239 <= '1' when reg_fullgraph2 = "0111101000" else '0'; 
		reg_q1242 <= '1' when reg_fullgraph2 = "0111101001" else '0'; 
		reg_q1244 <= '1' when reg_fullgraph2 = "0111101010" else '0'; 
		reg_q1282 <= '1' when reg_fullgraph2 = "0111101011" else '0'; 
		reg_q1284 <= '1' when reg_fullgraph2 = "0111101100" else '0'; 
		reg_q1570 <= '1' when reg_fullgraph2 = "0111101101" else '0'; 
		reg_q1572 <= '1' when reg_fullgraph2 = "0111101110" else '0'; 
		reg_q1706 <= '1' when reg_fullgraph2 = "0111101111" else '0'; 
		reg_q436 <= '1' when reg_fullgraph2 = "0111110000" else '0'; 
		reg_q220 <= '1' when reg_fullgraph2 = "0111110001" else '0'; 
		reg_q222 <= '1' when reg_fullgraph2 = "0111110010" else '0'; 
		reg_q210 <= '1' when reg_fullgraph2 = "0111110011" else '0'; 
		reg_q212 <= '1' when reg_fullgraph2 = "0111110100" else '0'; 
		reg_q78 <= '1' when reg_fullgraph2 = "0111110101" else '0'; 
		reg_q80 <= '1' when reg_fullgraph2 = "0111110110" else '0'; 
		reg_q684 <= '1' when reg_fullgraph2 = "0111110111" else '0'; 
		reg_q1039 <= '1' when reg_fullgraph2 = "0111111000" else '0'; 
		reg_q1041 <= '1' when reg_fullgraph2 = "0111111001" else '0'; 
		reg_q2241 <= '1' when reg_fullgraph2 = "0111111010" else '0'; 
		reg_q2233 <= '1' when reg_fullgraph2 = "0111111011" else '0'; 
		reg_q2235 <= '1' when reg_fullgraph2 = "0111111100" else '0'; 
		reg_q972 <= '1' when reg_fullgraph2 = "0111111101" else '0'; 
		reg_q2219 <= '1' when reg_fullgraph2 = "0111111110" else '0'; 
		reg_q1492 <= '1' when reg_fullgraph2 = "0111111111" else '0'; 
		reg_q1554 <= '1' when reg_fullgraph2 = "1000000000" else '0'; 
		reg_q2495 <= '1' when reg_fullgraph2 = "1000000001" else '0'; 
		reg_q2231 <= '1' when reg_fullgraph2 = "1000000010" else '0'; 
		reg_q724 <= '1' when reg_fullgraph2 = "1000000011" else '0'; 
		reg_q726 <= '1' when reg_fullgraph2 = "1000000100" else '0'; 
		reg_q2113 <= '1' when reg_fullgraph2 = "1000000101" else '0'; 
		reg_q2144 <= '1' when reg_fullgraph2 = "1000000110" else '0'; 
		reg_q2146 <= '1' when reg_fullgraph2 = "1000000111" else '0'; 
		reg_q1228 <= '1' when reg_fullgraph2 = "1000001000" else '0'; 
		reg_q1650 <= '1' when reg_fullgraph2 = "1000001001" else '0'; 
		reg_q147 <= '1' when reg_fullgraph2 = "1000001010" else '0'; 
		reg_q296 <= '1' when reg_fullgraph2 = "1000001011" else '0'; 
		reg_q1611 <= '1' when reg_fullgraph2 = "1000001100" else '0'; 
		reg_q1169 <= '1' when reg_fullgraph2 = "1000001101" else '0'; 
		reg_q1171 <= '1' when reg_fullgraph2 = "1000001110" else '0'; 
		reg_q1017 <= '1' when reg_fullgraph2 = "1000001111" else '0'; 
		reg_q1019 <= '1' when reg_fullgraph2 = "1000010000" else '0'; 
		reg_q2571 <= '1' when reg_fullgraph2 = "1000010001" else '0'; 
		reg_q1615 <= '1' when reg_fullgraph2 = "1000010010" else '0'; 
		reg_q2561 <= '1' when reg_fullgraph2 = "1000010011" else '0'; 
		reg_q1353 <= '1' when reg_fullgraph2 = "1000010100" else '0'; 
		reg_q1127 <= '1' when reg_fullgraph2 = "1000010101" else '0'; 
		reg_q1129 <= '1' when reg_fullgraph2 = "1000010110" else '0'; 
		reg_q1351 <= '1' when reg_fullgraph2 = "1000010111" else '0'; 
		reg_q385 <= '1' when reg_fullgraph2 = "1000011000" else '0'; 
		reg_q387 <= '1' when reg_fullgraph2 = "1000011001" else '0'; 
		reg_q432 <= '1' when reg_fullgraph2 = "1000011010" else '0'; 
		reg_q2318 <= '1' when reg_fullgraph2 = "1000011011" else '0'; 
		reg_q2320 <= '1' when reg_fullgraph2 = "1000011100" else '0'; 
		reg_q2682 <= '1' when reg_fullgraph2 = "1000011101" else '0'; 
		reg_q2684 <= '1' when reg_fullgraph2 = "1000011110" else '0'; 
		reg_q1514 <= '1' when reg_fullgraph2 = "1000011111" else '0'; 
		reg_q1516 <= '1' when reg_fullgraph2 = "1000100000" else '0'; 
		reg_q2107 <= '1' when reg_fullgraph2 = "1000100001" else '0'; 
		reg_q728 <= '1' when reg_fullgraph2 = "1000100010" else '0'; 
		reg_q2329 <= '1' when reg_fullgraph2 = "1000100011" else '0'; 
		reg_q2331 <= '1' when reg_fullgraph2 = "1000100100" else '0'; 
		reg_q1157 <= '1' when reg_fullgraph2 = "1000100101" else '0'; 
		reg_q2654 <= '1' when reg_fullgraph2 = "1000100110" else '0'; 
		reg_q2656 <= '1' when reg_fullgraph2 = "1000100111" else '0'; 
		reg_q2607 <= '1' when reg_fullgraph2 = "1000101000" else '0'; 
		reg_q1345 <= '1' when reg_fullgraph2 = "1000101001" else '0'; 
		reg_q347 <= '1' when reg_fullgraph2 = "1000101010" else '0'; 
		reg_q1488 <= '1' when reg_fullgraph2 = "1000101011" else '0'; 
		reg_q1286 <= '1' when reg_fullgraph2 = "1000101100" else '0'; 
		reg_q321 <= '1' when reg_fullgraph2 = "1000101101" else '0'; 
		reg_q1508 <= '1' when reg_fullgraph2 = "1000101110" else '0'; 
		reg_q1510 <= '1' when reg_fullgraph2 = "1000101111" else '0'; 
		reg_q2099 <= '1' when reg_fullgraph2 = "1000110000" else '0'; 
		reg_q70 <= '1' when reg_fullgraph2 = "1000110001" else '0'; 
		reg_q970 <= '1' when reg_fullgraph2 = "1000110010" else '0'; 
		reg_q760 <= '1' when reg_fullgraph2 = "1000110011" else '0'; 
		reg_q762 <= '1' when reg_fullgraph2 = "1000110100" else '0'; 
		reg_q707 <= '1' when reg_fullgraph2 = "1000110101" else '0'; 
		reg_q1234 <= '1' when reg_fullgraph2 = "1000110110" else '0'; 
		reg_q1173 <= '1' when reg_fullgraph2 = "1000110111" else '0'; 
		reg_q1175 <= '1' when reg_fullgraph2 = "1000111000" else '0'; 
		reg_q2512 <= '1' when reg_fullgraph2 = "1000111001" else '0'; 
		reg_q2652 <= '1' when reg_fullgraph2 = "1000111010" else '0'; 
		reg_q1584 <= '1' when reg_fullgraph2 = "1000111011" else '0'; 
		reg_q1006 <= '1' when reg_fullgraph2 = "1000111100" else '0'; 
		reg_q1486 <= '1' when reg_fullgraph2 = "1000111101" else '0'; 
		reg_q331 <= '1' when reg_fullgraph2 = "1000111110" else '0'; 
		reg_q1270 <= '1' when reg_fullgraph2 = "1000111111" else '0'; 
		reg_q141 <= '1' when reg_fullgraph2 = "1001000000" else '0'; 
		reg_q143 <= '1' when reg_fullgraph2 = "1001000001" else '0'; 
		reg_q353 <= '1' when reg_fullgraph2 = "1001000010" else '0'; 
		reg_q355 <= '1' when reg_fullgraph2 = "1001000011" else '0'; 
		reg_q2668 <= '1' when reg_fullgraph2 = "1001000100" else '0'; 
		reg_q72 <= '1' when reg_fullgraph2 = "1001000101" else '0'; 
		reg_q165 <= '1' when reg_fullgraph2 = "1001000110" else '0'; 
		reg_q1454 <= '1' when reg_fullgraph2 = "1001000111" else '0'; 
		reg_q1456 <= '1' when reg_fullgraph2 = "1001001000" else '0'; 
		reg_q1607 <= '1' when reg_fullgraph2 = "1001001001" else '0'; 
		reg_q1131 <= '1' when reg_fullgraph2 = "1001001010" else '0'; 
		reg_q907 <= '1' when reg_fullgraph2 = "1001001011" else '0'; 
		reg_q2254 <= '1' when reg_fullgraph2 = "1001001100" else '0'; 
		reg_q2256 <= '1' when reg_fullgraph2 = "1001001101" else '0'; 
		reg_q1629 <= '1' when reg_fullgraph2 = "1001001110" else '0'; 
		reg_q1631 <= '1' when reg_fullgraph2 = "1001001111" else '0'; 
		reg_q157 <= '1' when reg_fullgraph2 = "1001010000" else '0'; 
		reg_q159 <= '1' when reg_fullgraph2 = "1001010001" else '0'; 
		reg_q1590 <= '1' when reg_fullgraph2 = "1001010010" else '0'; 
		reg_q1592 <= '1' when reg_fullgraph2 = "1001010011" else '0'; 
		reg_q1564 <= '1' when reg_fullgraph2 = "1001010100" else '0'; 
		reg_q1566 <= '1' when reg_fullgraph2 = "1001010101" else '0'; 
		reg_q1720 <= '1' when reg_fullgraph2 = "1001010110" else '0'; 
		reg_q1722 <= '1' when reg_fullgraph2 = "1001010111" else '0'; 
		reg_q2006 <= '1' when reg_fullgraph2 = "1001011000" else '0'; 
		reg_q1965 <= '1' when reg_fullgraph2 = "1001011001" else '0'; 
		reg_q1967 <= '1' when reg_fullgraph2 = "1001011010" else '0'; 
		reg_q272 <= '1' when reg_fullgraph2 = "1001011011" else '0'; 
		reg_q274 <= '1' when reg_fullgraph2 = "1001011100" else '0'; 
		reg_q2264 <= '1' when reg_fullgraph2 = "1001011101" else '0'; 
		reg_q2266 <= '1' when reg_fullgraph2 = "1001011110" else '0'; 
		reg_q204 <= '1' when reg_fullgraph2 = "1001011111" else '0'; 
		reg_q206 <= '1' when reg_fullgraph2 = "1001100000" else '0'; 
		reg_q1311 <= '1' when reg_fullgraph2 = "1001100001" else '0'; 
		reg_q909 <= '1' when reg_fullgraph2 = "1001100010" else '0'; 
		reg_q911 <= '1' when reg_fullgraph2 = "1001100011" else '0'; 
		reg_q2164 <= '1' when reg_fullgraph2 = "1001100100" else '0'; 
		reg_q2166 <= '1' when reg_fullgraph2 = "1001100101" else '0'; 
		reg_q1098 <= '1' when reg_fullgraph2 = "1001100110" else '0'; 
		reg_q2563 <= '1' when reg_fullgraph2 = "1001100111" else '0'; 
		reg_q2121 <= '1' when reg_fullgraph2 = "1001101000" else '0'; 
		reg_q151 <= '1' when reg_fullgraph2 = "1001101001" else '0'; 
		reg_q1121 <= '1' when reg_fullgraph2 = "1001101010" else '0'; 
		reg_q243 <= '1' when reg_fullgraph2 = "1001101011" else '0'; 
		reg_q1043 <= '1' when reg_fullgraph2 = "1001101100" else '0'; 
		reg_q1045 <= '1' when reg_fullgraph2 = "1001101101" else '0'; 
		reg_q276 <= '1' when reg_fullgraph2 = "1001101110" else '0'; 
		reg_q1047 <= '1' when reg_fullgraph2 = "1001101111" else '0'; 
		reg_q2367 <= '1' when reg_fullgraph2 = "1001110000" else '0'; 
		reg_q1066 <= '1' when reg_fullgraph2 = "1001110001" else '0'; 
		reg_q1496 <= '1' when reg_fullgraph2 = "1001110010" else '0'; 
		reg_q1498 <= '1' when reg_fullgraph2 = "1001110011" else '0'; 
		reg_q1696 <= '1' when reg_fullgraph2 = "1001110100" else '0'; 
		reg_q1494 <= '1' when reg_fullgraph2 = "1001110101" else '0'; 
		reg_q2036 <= '1' when reg_fullgraph2 = "1001110110" else '0'; 
		reg_q1684 <= '1' when reg_fullgraph2 = "1001110111" else '0'; 
		reg_q337 <= '1' when reg_fullgraph2 = "1001111000" else '0'; 
		reg_q339 <= '1' when reg_fullgraph2 = "1001111001" else '0'; 
		reg_q1959 <= '1' when reg_fullgraph2 = "1001111010" else '0'; 
		reg_q1961 <= '1' when reg_fullgraph2 = "1001111011" else '0'; 
		reg_q1518 <= '1' when reg_fullgraph2 = "1001111100" else '0'; 
		reg_q1656 <= '1' when reg_fullgraph2 = "1001111101" else '0'; 
		reg_q1658 <= '1' when reg_fullgraph2 = "1001111110" else '0'; 
		reg_q2314 <= '1' when reg_fullgraph2 = "1001111111" else '0'; 
		reg_q2316 <= '1' when reg_fullgraph2 = "1010000000" else '0'; 
		reg_q2638 <= '1' when reg_fullgraph2 = "1010000001" else '0'; 
		reg_q2142 <= '1' when reg_fullgraph2 = "1010000010" else '0'; 
		reg_q2660 <= '1' when reg_fullgraph2 = "1010000011" else '0'; 
		reg_q1568 <= '1' when reg_fullgraph2 = "1010000100" else '0'; 
		reg_q1062 <= '1' when reg_fullgraph2 = "1010000101" else '0'; 
		reg_q1064 <= '1' when reg_fullgraph2 = "1010000110" else '0'; 
		reg_q1686 <= '1' when reg_fullgraph2 = "1010000111" else '0'; 
		reg_q1240 <= '1' when reg_fullgraph2 = "1010001000" else '0'; 
		reg_q764 <= '1' when reg_fullgraph2 = "1010001001" else '0'; 
		reg_q1119 <= '1' when reg_fullgraph2 = "1010001010" else '0'; 
		reg_q1476 <= '1' when reg_fullgraph2 = "1010001011" else '0'; 
		reg_q62 <= '1' when reg_fullgraph2 = "1010001100" else '0'; 
		reg_q2678 <= '1' when reg_fullgraph2 = "1010001101" else '0'; 
		reg_q327 <= '1' when reg_fullgraph2 = "1010001110" else '0'; 
		reg_q329 <= '1' when reg_fullgraph2 = "1010001111" else '0'; 
		reg_q1718 <= '1' when reg_fullgraph2 = "1010010000" else '0'; 
		reg_q1054 <= '1' when reg_fullgraph2 = "1010010001" else '0'; 
		reg_q1056 <= '1' when reg_fullgraph2 = "1010010010" else '0'; 
		reg_q1512 <= '1' when reg_fullgraph2 = "1010010011" else '0'; 
		reg_q2262 <= '1' when reg_fullgraph2 = "1010010100" else '0'; 
		reg_q1167 <= '1' when reg_fullgraph2 = "1010010101" else '0'; 
		reg_q2379 <= '1' when reg_fullgraph2 = "1010010110" else '0'; 
		reg_q2016 <= '1' when reg_fullgraph2 = "1010010111" else '0'; 
		reg_q64 <= '1' when reg_fullgraph2 = "1010011000" else '0'; 
		reg_q1623 <= '1' when reg_fullgraph2 = "1010011001" else '0'; 
		reg_q145 <= '1' when reg_fullgraph2 = "1010011010" else '0'; 
		reg_q1594 <= '1' when reg_fullgraph2 = "1010011011" else '0'; 
		reg_q1596 <= '1' when reg_fullgraph2 = "1010011100" else '0'; 
		reg_q2626 <= '1' when reg_fullgraph2 = "1010011101" else '0'; 
		reg_q2365 <= '1' when reg_fullgraph2 = "1010011110" else '0'; 
		reg_q1609 <= '1' when reg_fullgraph2 = "1010011111" else '0'; 
		reg_q1058 <= '1' when reg_fullgraph2 = "1010100000" else '0'; 
		reg_q1060 <= '1' when reg_fullgraph2 = "1010100001" else '0'; 
		reg_q208 <= '1' when reg_fullgraph2 = "1010100010" else '0'; 
		reg_q1621 <= '1' when reg_fullgraph2 = "1010100011" else '0'; 
		reg_q694 <= '1' when reg_fullgraph2 = "1010100100" else '0'; 
		reg_q214 <= '1' when reg_fullgraph2 = "1010100101" else '0'; 
		reg_q2555 <= '1' when reg_fullgraph2 = "1010100110" else '0'; 
		reg_q2152 <= '1' when reg_fullgraph2 = "1010100111" else '0'; 
		reg_q2154 <= '1' when reg_fullgraph2 = "1010101000" else '0'; 
		reg_q2312 <= '1' when reg_fullgraph2 = "1010101001" else '0'; 
		reg_q311 <= '1' when reg_fullgraph2 = "1010101010" else '0'; 
		reg_q1500 <= '1' when reg_fullgraph2 = "1010101011" else '0'; 
		reg_q317 <= '1' when reg_fullgraph2 = "1010101100" else '0'; 
		reg_q2680 <= '1' when reg_fullgraph2 = "1010101101" else '0'; 
		reg_q1266 <= '1' when reg_fullgraph2 = "1010101110" else '0'; 
		reg_q1268 <= '1' when reg_fullgraph2 = "1010101111" else '0'; 
		reg_q2628 <= '1' when reg_fullgraph2 = "1010110000" else '0'; 
		reg_q2630 <= '1' when reg_fullgraph2 = "1010110001" else '0'; 
		reg_q1429 <= '1' when reg_fullgraph2 = "1010110010" else '0'; 
		reg_q1236 <= '1' when reg_fullgraph2 = "1010110011" else '0'; 
		reg_q1238 <= '1' when reg_fullgraph2 = "1010110100" else '0'; 
		reg_q2478 <= '1' when reg_fullgraph2 = "1010110101" else '0'; 
		reg_q722 <= '1' when reg_fullgraph2 = "1010110110" else '0'; 
		reg_q391 <= '1' when reg_fullgraph2 = "1010110111" else '0'; 
		reg_q393 <= '1' when reg_fullgraph2 = "1010111000" else '0'; 
		reg_q1280 <= '1' when reg_fullgraph2 = "1010111001" else '0'; 
		reg_q2569 <= '1' when reg_fullgraph2 = "1010111010" else '0'; 
		reg_q202 <= '1' when reg_fullgraph2 = "1010111011" else '0'; 
		reg_q268 <= '1' when reg_fullgraph2 = "1010111100" else '0'; 
		reg_q270 <= '1' when reg_fullgraph2 = "1010111101" else '0'; 
		reg_q173 <= '1' when reg_fullgraph2 = "1010111110" else '0'; 
		reg_q175 <= '1' when reg_fullgraph2 = "1010111111" else '0'; 
		reg_q669 <= '1' when reg_fullgraph2 = "1011000000" else '0'; 
		reg_q1502 <= '1' when reg_fullgraph2 = "1011000001" else '0'; 
		reg_q738 <= '1' when reg_fullgraph2 = "1011000010" else '0'; 
		reg_q54 <= '1' when reg_fullgraph2 = "1011000011" else '0'; 
		reg_q1963 <= '1' when reg_fullgraph2 = "1011000100" else '0'; 
		reg_q2381 <= '1' when reg_fullgraph2 = "1011000101" else '0'; 
		reg_q2345 <= '1' when reg_fullgraph2 = "1011000110" else '0'; 
		reg_q2008 <= '1' when reg_fullgraph2 = "1011000111" else '0'; 
		reg_q730 <= '1' when reg_fullgraph2 = "1011001000" else '0'; 
		reg_q1321 <= '1' when reg_fullgraph2 = "1011001001" else '0'; 
		reg_q1323 <= '1' when reg_fullgraph2 = "1011001010" else '0'; 
		reg_q1309 <= '1' when reg_fullgraph2 = "1011001011" else '0'; 
		reg_q99 <= '1' when reg_fullgraph2 = "1011001100" else '0'; 
		reg_q1586 <= '1' when reg_fullgraph2 = "1011001101" else '0'; 
		reg_q2156 <= '1' when reg_fullgraph2 = "1011001110" else '0'; 
		reg_q319 <= '1' when reg_fullgraph2 = "1011001111" else '0'; 
		reg_q2026 <= '1' when reg_fullgraph2 = "1011010000" else '0'; 
		reg_q401 <= '1' when reg_fullgraph2 = "1011010001" else '0'; 
		reg_q2666 <= '1' when reg_fullgraph2 = "1011010010" else '0'; 
		reg_q286 <= '1' when reg_fullgraph2 = "1011010011" else '0'; 
		reg_q2658 <= '1' when reg_fullgraph2 = "1011010100" else '0'; 
		reg_q754 <= '1' when reg_fullgraph2 = "1011010101" else '0'; 
		reg_q345 <= '1' when reg_fullgraph2 = "1011010110" else '0'; 
		reg_q1021 <= '1' when reg_fullgraph2 = "1011010111" else '0'; 
		reg_q2539 <= '1' when reg_fullgraph2 = "1011011000" else '0'; 
		reg_q1163 <= '1' when reg_fullgraph2 = "1011011001" else '0'; 
		reg_q1165 <= '1' when reg_fullgraph2 = "1011011010" else '0'; 
		reg_q411 <= '1' when reg_fullgraph2 = "1011011011" else '0'; 
		reg_q720 <= '1' when reg_fullgraph2 = "1011011100" else '0'; 
		reg_q1292 <= '1' when reg_fullgraph2 = "1011011101" else '0'; 
		reg_q1294 <= '1' when reg_fullgraph2 = "1011011110" else '0'; 
		reg_q2553 <= '1' when reg_fullgraph2 = "1011011111" else '0'; 
		reg_q1449 <= '1' when reg_fullgraph2 = "1011100000" else '0'; 
		reg_q1100 <= '1' when reg_fullgraph2 = "1011100001" else '0'; 
		reg_q424 <= '1' when reg_fullgraph2 = "1011100010" else '0'; 
		reg_q1177 <= '1' when reg_fullgraph2 = "1011100011" else '0'; 
		reg_q2355 <= '1' when reg_fullgraph2 = "1011100100" else '0'; 
		reg_q732 <= '1' when reg_fullgraph2 = "1011100101" else '0'; 
		reg_q434 <= '1' when reg_fullgraph2 = "1011100110" else '0'; 
		reg_q2551 <= '1' when reg_fullgraph2 = "1011100111" else '0'; 
		reg_q2044 <= '1' when reg_fullgraph2 = "1011101000" else '0'; 
		reg_q2046 <= '1' when reg_fullgraph2 = "1011101001" else '0'; 
		reg_q2541 <= '1' when reg_fullgraph2 = "1011101010" else '0'; 
		reg_q1588 <= '1' when reg_fullgraph2 = "1011101011" else '0'; 
		reg_q2693 <= '1' when reg_fullgraph2 = "1011101100" else '0'; 
		reg_q2543 <= '1' when reg_fullgraph2 = "1011101101" else '0'; 
		reg_q2545 <= '1' when reg_fullgraph2 = "1011101110" else '0'; 
		reg_q2347 <= '1' when reg_fullgraph2 = "1011101111" else '0'; 
		reg_q1740 <= '1' when reg_fullgraph2 = "1011110000" else '0'; 
		reg_q1329 <= '1' when reg_fullgraph2 = "1011110001" else '0'; 
		reg_q2632 <= '1' when reg_fullgraph2 = "1011110010" else '0'; 
		reg_q1303 <= '1' when reg_fullgraph2 = "1011110011" else '0'; 
		reg_q309 <= '1' when reg_fullgraph2 = "1011110100" else '0'; 
		reg_q216 <= '1' when reg_fullgraph2 = "1011110101" else '0'; 
		reg_q2134 <= '1' when reg_fullgraph2 = "1011110110" else '0'; 
		reg_q770 <= '1' when reg_fullgraph2 = "1011110111" else '0'; 
		reg_q155 <= '1' when reg_fullgraph2 = "1011111000" else '0'; 
		reg_q2140 <= '1' when reg_fullgraph2 = "1011111001" else '0'; 
		reg_q383 <= '1' when reg_fullgraph2 = "1011111010" else '0'; 
		reg_q1633 <= '1' when reg_fullgraph2 = "1011111011" else '0'; 
		reg_q772 <= '1' when reg_fullgraph2 = "1011111100" else '0'; 
		reg_q1155 <= '1' when reg_fullgraph2 = "1011111101" else '0'; 
		reg_q927 <= '1' when reg_fullgraph2 = "1011111110" else '0'; 
		reg_q929 <= '1' when reg_fullgraph2 = "1011111111" else '0'; 
		reg_q1969 <= '1' when reg_fullgraph2 = "1100000000" else '0'; 
		reg_q1415 <= '1' when reg_fullgraph2 = "1100000001" else '0'; 
		reg_q1417 <= '1' when reg_fullgraph2 = "1100000010" else '0'; 
		reg_q153 <= '1' when reg_fullgraph2 = "1100000011" else '0'; 
		reg_q1288 <= '1' when reg_fullgraph2 = "1100000100" else '0'; 
		reg_q1276 <= '1' when reg_fullgraph2 = "1100000101" else '0'; 
		reg_q2048 <= '1' when reg_fullgraph2 = "1100000110" else '0'; 
		reg_q218 <= '1' when reg_fullgraph2 = "1100000111" else '0'; 
		reg_q1149 <= '1' when reg_fullgraph2 = "1100001000" else '0'; 
		reg_q259 <= '1' when reg_fullgraph2 = "1100001001" else '0'; 
		reg_q2327 <= '1' when reg_fullgraph2 = "1100001010" else '0'; 
		reg_q266 <= '1' when reg_fullgraph2 = "1100001011" else '0'; 
		reg_q746 <= '1' when reg_fullgraph2 = "1100001100" else '0'; 
		reg_q774 <= '1' when reg_fullgraph2 = "1100001101" else '0'; 
		reg_q776 <= '1' when reg_fullgraph2 = "1100001110" else '0'; 
		reg_q389 <= '1' when reg_fullgraph2 = "1100001111" else '0'; 
		reg_q1598 <= '1' when reg_fullgraph2 = "1100010000" else '0'; 
		reg_q1004 <= '1' when reg_fullgraph2 = "1100010001" else '0'; 
		reg_q1419 <= '1' when reg_fullgraph2 = "1100010010" else '0'; 
		reg_q1278 <= '1' when reg_fullgraph2 = "1100010011" else '0'; 
		reg_q1654 <= '1' when reg_fullgraph2 = "1100010100" else '0'; 
		reg_q1458 <= '1' when reg_fullgraph2 = "1100010101" else '0'; 
		reg_q1641 <= '1' when reg_fullgraph2 = "1100010110" else '0'; 
		reg_q1600 <= '1' when reg_fullgraph2 = "1100010111" else '0'; 
		reg_q2097 <= '1' when reg_fullgraph2 = "1100011000" else '0'; 
		reg_q1290 <= '1' when reg_fullgraph2 = "1100011001" else '0'; 
		reg_q740 <= '1' when reg_fullgraph2 = "1100011010" else '0'; 
		reg_q677 <= '1' when reg_fullgraph2 = "1100011011" else '0'; 
		reg_q2050 <= '1' when reg_fullgraph2 = "1100011100" else '0'; 
--end decoder 

reg_q178_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q178 AND symb_decoder(16#72#)) OR
 					(reg_q178 AND symb_decoder(16#6f#)) OR
 					(reg_q178 AND symb_decoder(16#38#)) OR
 					(reg_q178 AND symb_decoder(16#5a#)) OR
 					(reg_q178 AND symb_decoder(16#40#)) OR
 					(reg_q178 AND symb_decoder(16#d6#)) OR
 					(reg_q178 AND symb_decoder(16#19#)) OR
 					(reg_q178 AND symb_decoder(16#d3#)) OR
 					(reg_q178 AND symb_decoder(16#65#)) OR
 					(reg_q178 AND symb_decoder(16#59#)) OR
 					(reg_q178 AND symb_decoder(16#25#)) OR
 					(reg_q178 AND symb_decoder(16#fb#)) OR
 					(reg_q178 AND symb_decoder(16#fa#)) OR
 					(reg_q178 AND symb_decoder(16#a0#)) OR
 					(reg_q178 AND symb_decoder(16#bf#)) OR
 					(reg_q178 AND symb_decoder(16#4f#)) OR
 					(reg_q178 AND symb_decoder(16#f2#)) OR
 					(reg_q178 AND symb_decoder(16#ec#)) OR
 					(reg_q178 AND symb_decoder(16#36#)) OR
 					(reg_q178 AND symb_decoder(16#57#)) OR
 					(reg_q178 AND symb_decoder(16#ea#)) OR
 					(reg_q178 AND symb_decoder(16#94#)) OR
 					(reg_q178 AND symb_decoder(16#ba#)) OR
 					(reg_q178 AND symb_decoder(16#17#)) OR
 					(reg_q178 AND symb_decoder(16#56#)) OR
 					(reg_q178 AND symb_decoder(16#32#)) OR
 					(reg_q178 AND symb_decoder(16#e4#)) OR
 					(reg_q178 AND symb_decoder(16#a5#)) OR
 					(reg_q178 AND symb_decoder(16#70#)) OR
 					(reg_q178 AND symb_decoder(16#07#)) OR
 					(reg_q178 AND symb_decoder(16#ca#)) OR
 					(reg_q178 AND symb_decoder(16#9d#)) OR
 					(reg_q178 AND symb_decoder(16#12#)) OR
 					(reg_q178 AND symb_decoder(16#f9#)) OR
 					(reg_q178 AND symb_decoder(16#87#)) OR
 					(reg_q178 AND symb_decoder(16#58#)) OR
 					(reg_q178 AND symb_decoder(16#c1#)) OR
 					(reg_q178 AND symb_decoder(16#54#)) OR
 					(reg_q178 AND symb_decoder(16#cd#)) OR
 					(reg_q178 AND symb_decoder(16#5f#)) OR
 					(reg_q178 AND symb_decoder(16#f8#)) OR
 					(reg_q178 AND symb_decoder(16#cc#)) OR
 					(reg_q178 AND symb_decoder(16#e1#)) OR
 					(reg_q178 AND symb_decoder(16#8d#)) OR
 					(reg_q178 AND symb_decoder(16#92#)) OR
 					(reg_q178 AND symb_decoder(16#c2#)) OR
 					(reg_q178 AND symb_decoder(16#d9#)) OR
 					(reg_q178 AND symb_decoder(16#f7#)) OR
 					(reg_q178 AND symb_decoder(16#3d#)) OR
 					(reg_q178 AND symb_decoder(16#85#)) OR
 					(reg_q178 AND symb_decoder(16#24#)) OR
 					(reg_q178 AND symb_decoder(16#bc#)) OR
 					(reg_q178 AND symb_decoder(16#02#)) OR
 					(reg_q178 AND symb_decoder(16#95#)) OR
 					(reg_q178 AND symb_decoder(16#1b#)) OR
 					(reg_q178 AND symb_decoder(16#ed#)) OR
 					(reg_q178 AND symb_decoder(16#2e#)) OR
 					(reg_q178 AND symb_decoder(16#44#)) OR
 					(reg_q178 AND symb_decoder(16#bb#)) OR
 					(reg_q178 AND symb_decoder(16#b4#)) OR
 					(reg_q178 AND symb_decoder(16#9b#)) OR
 					(reg_q178 AND symb_decoder(16#a6#)) OR
 					(reg_q178 AND symb_decoder(16#5b#)) OR
 					(reg_q178 AND symb_decoder(16#0b#)) OR
 					(reg_q178 AND symb_decoder(16#ad#)) OR
 					(reg_q178 AND symb_decoder(16#93#)) OR
 					(reg_q178 AND symb_decoder(16#81#)) OR
 					(reg_q178 AND symb_decoder(16#1d#)) OR
 					(reg_q178 AND symb_decoder(16#d1#)) OR
 					(reg_q178 AND symb_decoder(16#f3#)) OR
 					(reg_q178 AND symb_decoder(16#e5#)) OR
 					(reg_q178 AND symb_decoder(16#89#)) OR
 					(reg_q178 AND symb_decoder(16#97#)) OR
 					(reg_q178 AND symb_decoder(16#ff#)) OR
 					(reg_q178 AND symb_decoder(16#49#)) OR
 					(reg_q178 AND symb_decoder(16#29#)) OR
 					(reg_q178 AND symb_decoder(16#5d#)) OR
 					(reg_q178 AND symb_decoder(16#dd#)) OR
 					(reg_q178 AND symb_decoder(16#2f#)) OR
 					(reg_q178 AND symb_decoder(16#67#)) OR
 					(reg_q178 AND symb_decoder(16#eb#)) OR
 					(reg_q178 AND symb_decoder(16#c7#)) OR
 					(reg_q178 AND symb_decoder(16#c4#)) OR
 					(reg_q178 AND symb_decoder(16#a8#)) OR
 					(reg_q178 AND symb_decoder(16#35#)) OR
 					(reg_q178 AND symb_decoder(16#a4#)) OR
 					(reg_q178 AND symb_decoder(16#01#)) OR
 					(reg_q178 AND symb_decoder(16#ee#)) OR
 					(reg_q178 AND symb_decoder(16#2d#)) OR
 					(reg_q178 AND symb_decoder(16#11#)) OR
 					(reg_q178 AND symb_decoder(16#b6#)) OR
 					(reg_q178 AND symb_decoder(16#fe#)) OR
 					(reg_q178 AND symb_decoder(16#d7#)) OR
 					(reg_q178 AND symb_decoder(16#be#)) OR
 					(reg_q178 AND symb_decoder(16#4e#)) OR
 					(reg_q178 AND symb_decoder(16#8a#)) OR
 					(reg_q178 AND symb_decoder(16#d0#)) OR
 					(reg_q178 AND symb_decoder(16#30#)) OR
 					(reg_q178 AND symb_decoder(16#7d#)) OR
 					(reg_q178 AND symb_decoder(16#af#)) OR
 					(reg_q178 AND symb_decoder(16#84#)) OR
 					(reg_q178 AND symb_decoder(16#8f#)) OR
 					(reg_q178 AND symb_decoder(16#a2#)) OR
 					(reg_q178 AND symb_decoder(16#48#)) OR
 					(reg_q178 AND symb_decoder(16#5c#)) OR
 					(reg_q178 AND symb_decoder(16#63#)) OR
 					(reg_q178 AND symb_decoder(16#9f#)) OR
 					(reg_q178 AND symb_decoder(16#53#)) OR
 					(reg_q178 AND symb_decoder(16#c8#)) OR
 					(reg_q178 AND symb_decoder(16#31#)) OR
 					(reg_q178 AND symb_decoder(16#a7#)) OR
 					(reg_q178 AND symb_decoder(16#dc#)) OR
 					(reg_q178 AND symb_decoder(16#64#)) OR
 					(reg_q178 AND symb_decoder(16#00#)) OR
 					(reg_q178 AND symb_decoder(16#b1#)) OR
 					(reg_q178 AND symb_decoder(16#55#)) OR
 					(reg_q178 AND symb_decoder(16#7c#)) OR
 					(reg_q178 AND symb_decoder(16#2c#)) OR
 					(reg_q178 AND symb_decoder(16#ce#)) OR
 					(reg_q178 AND symb_decoder(16#fd#)) OR
 					(reg_q178 AND symb_decoder(16#18#)) OR
 					(reg_q178 AND symb_decoder(16#09#)) OR
 					(reg_q178 AND symb_decoder(16#e2#)) OR
 					(reg_q178 AND symb_decoder(16#a9#)) OR
 					(reg_q178 AND symb_decoder(16#b0#)) OR
 					(reg_q178 AND symb_decoder(16#0e#)) OR
 					(reg_q178 AND symb_decoder(16#6b#)) OR
 					(reg_q178 AND symb_decoder(16#42#)) OR
 					(reg_q178 AND symb_decoder(16#39#)) OR
 					(reg_q178 AND symb_decoder(16#4a#)) OR
 					(reg_q178 AND symb_decoder(16#03#)) OR
 					(reg_q178 AND symb_decoder(16#37#)) OR
 					(reg_q178 AND symb_decoder(16#f1#)) OR
 					(reg_q178 AND symb_decoder(16#91#)) OR
 					(reg_q178 AND symb_decoder(16#1c#)) OR
 					(reg_q178 AND symb_decoder(16#0c#)) OR
 					(reg_q178 AND symb_decoder(16#50#)) OR
 					(reg_q178 AND symb_decoder(16#db#)) OR
 					(reg_q178 AND symb_decoder(16#9c#)) OR
 					(reg_q178 AND symb_decoder(16#b2#)) OR
 					(reg_q178 AND symb_decoder(16#9a#)) OR
 					(reg_q178 AND symb_decoder(16#0a#)) OR
 					(reg_q178 AND symb_decoder(16#bd#)) OR
 					(reg_q178 AND symb_decoder(16#7e#)) OR
 					(reg_q178 AND symb_decoder(16#88#)) OR
 					(reg_q178 AND symb_decoder(16#c0#)) OR
 					(reg_q178 AND symb_decoder(16#ef#)) OR
 					(reg_q178 AND symb_decoder(16#23#)) OR
 					(reg_q178 AND symb_decoder(16#15#)) OR
 					(reg_q178 AND symb_decoder(16#79#)) OR
 					(reg_q178 AND symb_decoder(16#90#)) OR
 					(reg_q178 AND symb_decoder(16#ae#)) OR
 					(reg_q178 AND symb_decoder(16#3a#)) OR
 					(reg_q178 AND symb_decoder(16#fc#)) OR
 					(reg_q178 AND symb_decoder(16#8b#)) OR
 					(reg_q178 AND symb_decoder(16#26#)) OR
 					(reg_q178 AND symb_decoder(16#1f#)) OR
 					(reg_q178 AND symb_decoder(16#86#)) OR
 					(reg_q178 AND symb_decoder(16#68#)) OR
 					(reg_q178 AND symb_decoder(16#83#)) OR
 					(reg_q178 AND symb_decoder(16#6c#)) OR
 					(reg_q178 AND symb_decoder(16#a3#)) OR
 					(reg_q178 AND symb_decoder(16#4d#)) OR
 					(reg_q178 AND symb_decoder(16#de#)) OR
 					(reg_q178 AND symb_decoder(16#6a#)) OR
 					(reg_q178 AND symb_decoder(16#06#)) OR
 					(reg_q178 AND symb_decoder(16#c9#)) OR
 					(reg_q178 AND symb_decoder(16#99#)) OR
 					(reg_q178 AND symb_decoder(16#0f#)) OR
 					(reg_q178 AND symb_decoder(16#75#)) OR
 					(reg_q178 AND symb_decoder(16#f6#)) OR
 					(reg_q178 AND symb_decoder(16#98#)) OR
 					(reg_q178 AND symb_decoder(16#33#)) OR
 					(reg_q178 AND symb_decoder(16#a1#)) OR
 					(reg_q178 AND symb_decoder(16#9e#)) OR
 					(reg_q178 AND symb_decoder(16#51#)) OR
 					(reg_q178 AND symb_decoder(16#0d#)) OR
 					(reg_q178 AND symb_decoder(16#d5#)) OR
 					(reg_q178 AND symb_decoder(16#3c#)) OR
 					(reg_q178 AND symb_decoder(16#80#)) OR
 					(reg_q178 AND symb_decoder(16#62#)) OR
 					(reg_q178 AND symb_decoder(16#73#)) OR
 					(reg_q178 AND symb_decoder(16#f4#)) OR
 					(reg_q178 AND symb_decoder(16#3e#)) OR
 					(reg_q178 AND symb_decoder(16#28#)) OR
 					(reg_q178 AND symb_decoder(16#e8#)) OR
 					(reg_q178 AND symb_decoder(16#77#)) OR
 					(reg_q178 AND symb_decoder(16#e0#)) OR
 					(reg_q178 AND symb_decoder(16#e3#)) OR
 					(reg_q178 AND symb_decoder(16#6e#)) OR
 					(reg_q178 AND symb_decoder(16#f0#)) OR
 					(reg_q178 AND symb_decoder(16#e6#)) OR
 					(reg_q178 AND symb_decoder(16#27#)) OR
 					(reg_q178 AND symb_decoder(16#43#)) OR
 					(reg_q178 AND symb_decoder(16#6d#)) OR
 					(reg_q178 AND symb_decoder(16#7a#)) OR
 					(reg_q178 AND symb_decoder(16#10#)) OR
 					(reg_q178 AND symb_decoder(16#1e#)) OR
 					(reg_q178 AND symb_decoder(16#22#)) OR
 					(reg_q178 AND symb_decoder(16#05#)) OR
 					(reg_q178 AND symb_decoder(16#b9#)) OR
 					(reg_q178 AND symb_decoder(16#82#)) OR
 					(reg_q178 AND symb_decoder(16#b5#)) OR
 					(reg_q178 AND symb_decoder(16#34#)) OR
 					(reg_q178 AND symb_decoder(16#d8#)) OR
 					(reg_q178 AND symb_decoder(16#ab#)) OR
 					(reg_q178 AND symb_decoder(16#08#)) OR
 					(reg_q178 AND symb_decoder(16#2b#)) OR
 					(reg_q178 AND symb_decoder(16#74#)) OR
 					(reg_q178 AND symb_decoder(16#cb#)) OR
 					(reg_q178 AND symb_decoder(16#b7#)) OR
 					(reg_q178 AND symb_decoder(16#78#)) OR
 					(reg_q178 AND symb_decoder(16#7b#)) OR
 					(reg_q178 AND symb_decoder(16#8e#)) OR
 					(reg_q178 AND symb_decoder(16#b3#)) OR
 					(reg_q178 AND symb_decoder(16#e7#)) OR
 					(reg_q178 AND symb_decoder(16#7f#)) OR
 					(reg_q178 AND symb_decoder(16#61#)) OR
 					(reg_q178 AND symb_decoder(16#1a#)) OR
 					(reg_q178 AND symb_decoder(16#b8#)) OR
 					(reg_q178 AND symb_decoder(16#e9#)) OR
 					(reg_q178 AND symb_decoder(16#47#)) OR
 					(reg_q178 AND symb_decoder(16#71#)) OR
 					(reg_q178 AND symb_decoder(16#8c#)) OR
 					(reg_q178 AND symb_decoder(16#60#)) OR
 					(reg_q178 AND symb_decoder(16#3f#)) OR
 					(reg_q178 AND symb_decoder(16#df#)) OR
 					(reg_q178 AND symb_decoder(16#c5#)) OR
 					(reg_q178 AND symb_decoder(16#13#)) OR
 					(reg_q178 AND symb_decoder(16#16#)) OR
 					(reg_q178 AND symb_decoder(16#aa#)) OR
 					(reg_q178 AND symb_decoder(16#4b#)) OR
 					(reg_q178 AND symb_decoder(16#14#)) OR
 					(reg_q178 AND symb_decoder(16#cf#)) OR
 					(reg_q178 AND symb_decoder(16#da#)) OR
 					(reg_q178 AND symb_decoder(16#76#)) OR
 					(reg_q178 AND symb_decoder(16#66#)) OR
 					(reg_q178 AND symb_decoder(16#96#)) OR
 					(reg_q178 AND symb_decoder(16#d4#)) OR
 					(reg_q178 AND symb_decoder(16#45#)) OR
 					(reg_q178 AND symb_decoder(16#21#)) OR
 					(reg_q178 AND symb_decoder(16#3b#)) OR
 					(reg_q178 AND symb_decoder(16#04#)) OR
 					(reg_q178 AND symb_decoder(16#20#)) OR
 					(reg_q178 AND symb_decoder(16#46#)) OR
 					(reg_q178 AND symb_decoder(16#c6#)) OR
 					(reg_q178 AND symb_decoder(16#2a#)) OR
 					(reg_q178 AND symb_decoder(16#41#)) OR
 					(reg_q178 AND symb_decoder(16#52#)) OR
 					(reg_q178 AND symb_decoder(16#d2#)) OR
 					(reg_q178 AND symb_decoder(16#5e#)) OR
 					(reg_q178 AND symb_decoder(16#69#)) OR
 					(reg_q178 AND symb_decoder(16#f5#)) OR
 					(reg_q178 AND symb_decoder(16#c3#)) OR
 					(reg_q178 AND symb_decoder(16#4c#)) OR
 					(reg_q178 AND symb_decoder(16#ac#));
reg_q178_init <= '0' ;
	p_reg_q178: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q178 <= reg_q178_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q178 <= reg_q178_init;
        else
          reg_q178 <= reg_q178_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q899_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q899 AND symb_decoder(16#1d#)) OR
 					(reg_q899 AND symb_decoder(16#1e#)) OR
 					(reg_q899 AND symb_decoder(16#71#)) OR
 					(reg_q899 AND symb_decoder(16#9f#)) OR
 					(reg_q899 AND symb_decoder(16#ea#)) OR
 					(reg_q899 AND symb_decoder(16#28#)) OR
 					(reg_q899 AND symb_decoder(16#af#)) OR
 					(reg_q899 AND symb_decoder(16#b7#)) OR
 					(reg_q899 AND symb_decoder(16#14#)) OR
 					(reg_q899 AND symb_decoder(16#23#)) OR
 					(reg_q899 AND symb_decoder(16#b9#)) OR
 					(reg_q899 AND symb_decoder(16#0d#)) OR
 					(reg_q899 AND symb_decoder(16#25#)) OR
 					(reg_q899 AND symb_decoder(16#cd#)) OR
 					(reg_q899 AND symb_decoder(16#54#)) OR
 					(reg_q899 AND symb_decoder(16#98#)) OR
 					(reg_q899 AND symb_decoder(16#77#)) OR
 					(reg_q899 AND symb_decoder(16#29#)) OR
 					(reg_q899 AND symb_decoder(16#82#)) OR
 					(reg_q899 AND symb_decoder(16#9c#)) OR
 					(reg_q899 AND symb_decoder(16#9d#)) OR
 					(reg_q899 AND symb_decoder(16#df#)) OR
 					(reg_q899 AND symb_decoder(16#6c#)) OR
 					(reg_q899 AND symb_decoder(16#a8#)) OR
 					(reg_q899 AND symb_decoder(16#4c#)) OR
 					(reg_q899 AND symb_decoder(16#dd#)) OR
 					(reg_q899 AND symb_decoder(16#21#)) OR
 					(reg_q899 AND symb_decoder(16#2c#)) OR
 					(reg_q899 AND symb_decoder(16#39#)) OR
 					(reg_q899 AND symb_decoder(16#eb#)) OR
 					(reg_q899 AND symb_decoder(16#8f#)) OR
 					(reg_q899 AND symb_decoder(16#e9#)) OR
 					(reg_q899 AND symb_decoder(16#5b#)) OR
 					(reg_q899 AND symb_decoder(16#a3#)) OR
 					(reg_q899 AND symb_decoder(16#81#)) OR
 					(reg_q899 AND symb_decoder(16#0a#)) OR
 					(reg_q899 AND symb_decoder(16#e1#)) OR
 					(reg_q899 AND symb_decoder(16#e6#)) OR
 					(reg_q899 AND symb_decoder(16#68#)) OR
 					(reg_q899 AND symb_decoder(16#c1#)) OR
 					(reg_q899 AND symb_decoder(16#89#)) OR
 					(reg_q899 AND symb_decoder(16#bf#)) OR
 					(reg_q899 AND symb_decoder(16#95#)) OR
 					(reg_q899 AND symb_decoder(16#63#)) OR
 					(reg_q899 AND symb_decoder(16#87#)) OR
 					(reg_q899 AND symb_decoder(16#02#)) OR
 					(reg_q899 AND symb_decoder(16#d6#)) OR
 					(reg_q899 AND symb_decoder(16#de#)) OR
 					(reg_q899 AND symb_decoder(16#e4#)) OR
 					(reg_q899 AND symb_decoder(16#61#)) OR
 					(reg_q899 AND symb_decoder(16#a4#)) OR
 					(reg_q899 AND symb_decoder(16#52#)) OR
 					(reg_q899 AND symb_decoder(16#be#)) OR
 					(reg_q899 AND symb_decoder(16#e3#)) OR
 					(reg_q899 AND symb_decoder(16#96#)) OR
 					(reg_q899 AND symb_decoder(16#5a#)) OR
 					(reg_q899 AND symb_decoder(16#6e#)) OR
 					(reg_q899 AND symb_decoder(16#37#)) OR
 					(reg_q899 AND symb_decoder(16#2d#)) OR
 					(reg_q899 AND symb_decoder(16#f8#)) OR
 					(reg_q899 AND symb_decoder(16#d4#)) OR
 					(reg_q899 AND symb_decoder(16#27#)) OR
 					(reg_q899 AND symb_decoder(16#72#)) OR
 					(reg_q899 AND symb_decoder(16#6a#)) OR
 					(reg_q899 AND symb_decoder(16#c0#)) OR
 					(reg_q899 AND symb_decoder(16#5d#)) OR
 					(reg_q899 AND symb_decoder(16#31#)) OR
 					(reg_q899 AND symb_decoder(16#b5#)) OR
 					(reg_q899 AND symb_decoder(16#5c#)) OR
 					(reg_q899 AND symb_decoder(16#10#)) OR
 					(reg_q899 AND symb_decoder(16#8a#)) OR
 					(reg_q899 AND symb_decoder(16#97#)) OR
 					(reg_q899 AND symb_decoder(16#01#)) OR
 					(reg_q899 AND symb_decoder(16#db#)) OR
 					(reg_q899 AND symb_decoder(16#67#)) OR
 					(reg_q899 AND symb_decoder(16#c7#)) OR
 					(reg_q899 AND symb_decoder(16#d2#)) OR
 					(reg_q899 AND symb_decoder(16#7a#)) OR
 					(reg_q899 AND symb_decoder(16#19#)) OR
 					(reg_q899 AND symb_decoder(16#57#)) OR
 					(reg_q899 AND symb_decoder(16#2a#)) OR
 					(reg_q899 AND symb_decoder(16#36#)) OR
 					(reg_q899 AND symb_decoder(16#56#)) OR
 					(reg_q899 AND symb_decoder(16#1b#)) OR
 					(reg_q899 AND symb_decoder(16#9e#)) OR
 					(reg_q899 AND symb_decoder(16#4f#)) OR
 					(reg_q899 AND symb_decoder(16#41#)) OR
 					(reg_q899 AND symb_decoder(16#e7#)) OR
 					(reg_q899 AND symb_decoder(16#60#)) OR
 					(reg_q899 AND symb_decoder(16#17#)) OR
 					(reg_q899 AND symb_decoder(16#f2#)) OR
 					(reg_q899 AND symb_decoder(16#1f#)) OR
 					(reg_q899 AND symb_decoder(16#78#)) OR
 					(reg_q899 AND symb_decoder(16#33#)) OR
 					(reg_q899 AND symb_decoder(16#b6#)) OR
 					(reg_q899 AND symb_decoder(16#8d#)) OR
 					(reg_q899 AND symb_decoder(16#f9#)) OR
 					(reg_q899 AND symb_decoder(16#51#)) OR
 					(reg_q899 AND symb_decoder(16#ff#)) OR
 					(reg_q899 AND symb_decoder(16#00#)) OR
 					(reg_q899 AND symb_decoder(16#24#)) OR
 					(reg_q899 AND symb_decoder(16#59#)) OR
 					(reg_q899 AND symb_decoder(16#5e#)) OR
 					(reg_q899 AND symb_decoder(16#1c#)) OR
 					(reg_q899 AND symb_decoder(16#b3#)) OR
 					(reg_q899 AND symb_decoder(16#58#)) OR
 					(reg_q899 AND symb_decoder(16#0b#)) OR
 					(reg_q899 AND symb_decoder(16#3f#)) OR
 					(reg_q899 AND symb_decoder(16#da#)) OR
 					(reg_q899 AND symb_decoder(16#f7#)) OR
 					(reg_q899 AND symb_decoder(16#1a#)) OR
 					(reg_q899 AND symb_decoder(16#3d#)) OR
 					(reg_q899 AND symb_decoder(16#e8#)) OR
 					(reg_q899 AND symb_decoder(16#40#)) OR
 					(reg_q899 AND symb_decoder(16#f6#)) OR
 					(reg_q899 AND symb_decoder(16#e0#)) OR
 					(reg_q899 AND symb_decoder(16#c6#)) OR
 					(reg_q899 AND symb_decoder(16#07#)) OR
 					(reg_q899 AND symb_decoder(16#04#)) OR
 					(reg_q899 AND symb_decoder(16#a7#)) OR
 					(reg_q899 AND symb_decoder(16#c8#)) OR
 					(reg_q899 AND symb_decoder(16#88#)) OR
 					(reg_q899 AND symb_decoder(16#bb#)) OR
 					(reg_q899 AND symb_decoder(16#d9#)) OR
 					(reg_q899 AND symb_decoder(16#ad#)) OR
 					(reg_q899 AND symb_decoder(16#f4#)) OR
 					(reg_q899 AND symb_decoder(16#cf#)) OR
 					(reg_q899 AND symb_decoder(16#20#)) OR
 					(reg_q899 AND symb_decoder(16#e5#)) OR
 					(reg_q899 AND symb_decoder(16#b2#)) OR
 					(reg_q899 AND symb_decoder(16#a2#)) OR
 					(reg_q899 AND symb_decoder(16#fa#)) OR
 					(reg_q899 AND symb_decoder(16#22#)) OR
 					(reg_q899 AND symb_decoder(16#03#)) OR
 					(reg_q899 AND symb_decoder(16#49#)) OR
 					(reg_q899 AND symb_decoder(16#b0#)) OR
 					(reg_q899 AND symb_decoder(16#46#)) OR
 					(reg_q899 AND symb_decoder(16#65#)) OR
 					(reg_q899 AND symb_decoder(16#11#)) OR
 					(reg_q899 AND symb_decoder(16#80#)) OR
 					(reg_q899 AND symb_decoder(16#70#)) OR
 					(reg_q899 AND symb_decoder(16#42#)) OR
 					(reg_q899 AND symb_decoder(16#0c#)) OR
 					(reg_q899 AND symb_decoder(16#ae#)) OR
 					(reg_q899 AND symb_decoder(16#b8#)) OR
 					(reg_q899 AND symb_decoder(16#bd#)) OR
 					(reg_q899 AND symb_decoder(16#fd#)) OR
 					(reg_q899 AND symb_decoder(16#93#)) OR
 					(reg_q899 AND symb_decoder(16#ac#)) OR
 					(reg_q899 AND symb_decoder(16#91#)) OR
 					(reg_q899 AND symb_decoder(16#f3#)) OR
 					(reg_q899 AND symb_decoder(16#3c#)) OR
 					(reg_q899 AND symb_decoder(16#5f#)) OR
 					(reg_q899 AND symb_decoder(16#9b#)) OR
 					(reg_q899 AND symb_decoder(16#d1#)) OR
 					(reg_q899 AND symb_decoder(16#08#)) OR
 					(reg_q899 AND symb_decoder(16#c5#)) OR
 					(reg_q899 AND symb_decoder(16#ab#)) OR
 					(reg_q899 AND symb_decoder(16#cb#)) OR
 					(reg_q899 AND symb_decoder(16#12#)) OR
 					(reg_q899 AND symb_decoder(16#85#)) OR
 					(reg_q899 AND symb_decoder(16#6b#)) OR
 					(reg_q899 AND symb_decoder(16#18#)) OR
 					(reg_q899 AND symb_decoder(16#d0#)) OR
 					(reg_q899 AND symb_decoder(16#90#)) OR
 					(reg_q899 AND symb_decoder(16#0e#)) OR
 					(reg_q899 AND symb_decoder(16#ee#)) OR
 					(reg_q899 AND symb_decoder(16#4a#)) OR
 					(reg_q899 AND symb_decoder(16#16#)) OR
 					(reg_q899 AND symb_decoder(16#15#)) OR
 					(reg_q899 AND symb_decoder(16#7f#)) OR
 					(reg_q899 AND symb_decoder(16#6f#)) OR
 					(reg_q899 AND symb_decoder(16#e2#)) OR
 					(reg_q899 AND symb_decoder(16#ce#)) OR
 					(reg_q899 AND symb_decoder(16#c2#)) OR
 					(reg_q899 AND symb_decoder(16#d7#)) OR
 					(reg_q899 AND symb_decoder(16#7b#)) OR
 					(reg_q899 AND symb_decoder(16#f1#)) OR
 					(reg_q899 AND symb_decoder(16#76#)) OR
 					(reg_q899 AND symb_decoder(16#84#)) OR
 					(reg_q899 AND symb_decoder(16#f0#)) OR
 					(reg_q899 AND symb_decoder(16#8b#)) OR
 					(reg_q899 AND symb_decoder(16#4b#)) OR
 					(reg_q899 AND symb_decoder(16#a5#)) OR
 					(reg_q899 AND symb_decoder(16#fb#)) OR
 					(reg_q899 AND symb_decoder(16#7d#)) OR
 					(reg_q899 AND symb_decoder(16#50#)) OR
 					(reg_q899 AND symb_decoder(16#30#)) OR
 					(reg_q899 AND symb_decoder(16#79#)) OR
 					(reg_q899 AND symb_decoder(16#34#)) OR
 					(reg_q899 AND symb_decoder(16#4e#)) OR
 					(reg_q899 AND symb_decoder(16#13#)) OR
 					(reg_q899 AND symb_decoder(16#b4#)) OR
 					(reg_q899 AND symb_decoder(16#bc#)) OR
 					(reg_q899 AND symb_decoder(16#fe#)) OR
 					(reg_q899 AND symb_decoder(16#7e#)) OR
 					(reg_q899 AND symb_decoder(16#d3#)) OR
 					(reg_q899 AND symb_decoder(16#92#)) OR
 					(reg_q899 AND symb_decoder(16#75#)) OR
 					(reg_q899 AND symb_decoder(16#c3#)) OR
 					(reg_q899 AND symb_decoder(16#53#)) OR
 					(reg_q899 AND symb_decoder(16#69#)) OR
 					(reg_q899 AND symb_decoder(16#2f#)) OR
 					(reg_q899 AND symb_decoder(16#44#)) OR
 					(reg_q899 AND symb_decoder(16#3e#)) OR
 					(reg_q899 AND symb_decoder(16#7c#)) OR
 					(reg_q899 AND symb_decoder(16#fc#)) OR
 					(reg_q899 AND symb_decoder(16#3b#)) OR
 					(reg_q899 AND symb_decoder(16#45#)) OR
 					(reg_q899 AND symb_decoder(16#62#)) OR
 					(reg_q899 AND symb_decoder(16#2b#)) OR
 					(reg_q899 AND symb_decoder(16#ec#)) OR
 					(reg_q899 AND symb_decoder(16#05#)) OR
 					(reg_q899 AND symb_decoder(16#64#)) OR
 					(reg_q899 AND symb_decoder(16#a9#)) OR
 					(reg_q899 AND symb_decoder(16#35#)) OR
 					(reg_q899 AND symb_decoder(16#3a#)) OR
 					(reg_q899 AND symb_decoder(16#ba#)) OR
 					(reg_q899 AND symb_decoder(16#74#)) OR
 					(reg_q899 AND symb_decoder(16#ca#)) OR
 					(reg_q899 AND symb_decoder(16#94#)) OR
 					(reg_q899 AND symb_decoder(16#6d#)) OR
 					(reg_q899 AND symb_decoder(16#0f#)) OR
 					(reg_q899 AND symb_decoder(16#26#)) OR
 					(reg_q899 AND symb_decoder(16#43#)) OR
 					(reg_q899 AND symb_decoder(16#8e#)) OR
 					(reg_q899 AND symb_decoder(16#9a#)) OR
 					(reg_q899 AND symb_decoder(16#09#)) OR
 					(reg_q899 AND symb_decoder(16#c9#)) OR
 					(reg_q899 AND symb_decoder(16#32#)) OR
 					(reg_q899 AND symb_decoder(16#66#)) OR
 					(reg_q899 AND symb_decoder(16#c4#)) OR
 					(reg_q899 AND symb_decoder(16#a0#)) OR
 					(reg_q899 AND symb_decoder(16#a1#)) OR
 					(reg_q899 AND symb_decoder(16#86#)) OR
 					(reg_q899 AND symb_decoder(16#73#)) OR
 					(reg_q899 AND symb_decoder(16#cc#)) OR
 					(reg_q899 AND symb_decoder(16#48#)) OR
 					(reg_q899 AND symb_decoder(16#aa#)) OR
 					(reg_q899 AND symb_decoder(16#d8#)) OR
 					(reg_q899 AND symb_decoder(16#4d#)) OR
 					(reg_q899 AND symb_decoder(16#ef#)) OR
 					(reg_q899 AND symb_decoder(16#2e#)) OR
 					(reg_q899 AND symb_decoder(16#47#)) OR
 					(reg_q899 AND symb_decoder(16#38#)) OR
 					(reg_q899 AND symb_decoder(16#99#)) OR
 					(reg_q899 AND symb_decoder(16#83#)) OR
 					(reg_q899 AND symb_decoder(16#dc#)) OR
 					(reg_q899 AND symb_decoder(16#d5#)) OR
 					(reg_q899 AND symb_decoder(16#ed#)) OR
 					(reg_q899 AND symb_decoder(16#55#)) OR
 					(reg_q899 AND symb_decoder(16#b1#)) OR
 					(reg_q899 AND symb_decoder(16#8c#)) OR
 					(reg_q899 AND symb_decoder(16#f5#)) OR
 					(reg_q899 AND symb_decoder(16#06#)) OR
 					(reg_q899 AND symb_decoder(16#a6#));
reg_q899_init <= '0' ;
	p_reg_q899: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q899 <= reg_q899_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q899 <= reg_q899_init;
        else
          reg_q899 <= reg_q899_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q225_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q225 AND symb_decoder(16#46#)) OR
 					(reg_q225 AND symb_decoder(16#d3#)) OR
 					(reg_q225 AND symb_decoder(16#20#)) OR
 					(reg_q225 AND symb_decoder(16#84#)) OR
 					(reg_q225 AND symb_decoder(16#ee#)) OR
 					(reg_q225 AND symb_decoder(16#71#)) OR
 					(reg_q225 AND symb_decoder(16#ed#)) OR
 					(reg_q225 AND symb_decoder(16#b4#)) OR
 					(reg_q225 AND symb_decoder(16#dc#)) OR
 					(reg_q225 AND symb_decoder(16#e5#)) OR
 					(reg_q225 AND symb_decoder(16#3b#)) OR
 					(reg_q225 AND symb_decoder(16#92#)) OR
 					(reg_q225 AND symb_decoder(16#a8#)) OR
 					(reg_q225 AND symb_decoder(16#c0#)) OR
 					(reg_q225 AND symb_decoder(16#01#)) OR
 					(reg_q225 AND symb_decoder(16#99#)) OR
 					(reg_q225 AND symb_decoder(16#dd#)) OR
 					(reg_q225 AND symb_decoder(16#56#)) OR
 					(reg_q225 AND symb_decoder(16#c5#)) OR
 					(reg_q225 AND symb_decoder(16#14#)) OR
 					(reg_q225 AND symb_decoder(16#95#)) OR
 					(reg_q225 AND symb_decoder(16#0e#)) OR
 					(reg_q225 AND symb_decoder(16#d8#)) OR
 					(reg_q225 AND symb_decoder(16#94#)) OR
 					(reg_q225 AND symb_decoder(16#53#)) OR
 					(reg_q225 AND symb_decoder(16#fd#)) OR
 					(reg_q225 AND symb_decoder(16#db#)) OR
 					(reg_q225 AND symb_decoder(16#36#)) OR
 					(reg_q225 AND symb_decoder(16#e2#)) OR
 					(reg_q225 AND symb_decoder(16#48#)) OR
 					(reg_q225 AND symb_decoder(16#72#)) OR
 					(reg_q225 AND symb_decoder(16#b0#)) OR
 					(reg_q225 AND symb_decoder(16#f2#)) OR
 					(reg_q225 AND symb_decoder(16#64#)) OR
 					(reg_q225 AND symb_decoder(16#05#)) OR
 					(reg_q225 AND symb_decoder(16#55#)) OR
 					(reg_q225 AND symb_decoder(16#4b#)) OR
 					(reg_q225 AND symb_decoder(16#8b#)) OR
 					(reg_q225 AND symb_decoder(16#bb#)) OR
 					(reg_q225 AND symb_decoder(16#34#)) OR
 					(reg_q225 AND symb_decoder(16#0f#)) OR
 					(reg_q225 AND symb_decoder(16#0a#)) OR
 					(reg_q225 AND symb_decoder(16#51#)) OR
 					(reg_q225 AND symb_decoder(16#30#)) OR
 					(reg_q225 AND symb_decoder(16#cd#)) OR
 					(reg_q225 AND symb_decoder(16#54#)) OR
 					(reg_q225 AND symb_decoder(16#aa#)) OR
 					(reg_q225 AND symb_decoder(16#7a#)) OR
 					(reg_q225 AND symb_decoder(16#9c#)) OR
 					(reg_q225 AND symb_decoder(16#6b#)) OR
 					(reg_q225 AND symb_decoder(16#ad#)) OR
 					(reg_q225 AND symb_decoder(16#f0#)) OR
 					(reg_q225 AND symb_decoder(16#0d#)) OR
 					(reg_q225 AND symb_decoder(16#86#)) OR
 					(reg_q225 AND symb_decoder(16#85#)) OR
 					(reg_q225 AND symb_decoder(16#1f#)) OR
 					(reg_q225 AND symb_decoder(16#1a#)) OR
 					(reg_q225 AND symb_decoder(16#3a#)) OR
 					(reg_q225 AND symb_decoder(16#6c#)) OR
 					(reg_q225 AND symb_decoder(16#a7#)) OR
 					(reg_q225 AND symb_decoder(16#3c#)) OR
 					(reg_q225 AND symb_decoder(16#d5#)) OR
 					(reg_q225 AND symb_decoder(16#2d#)) OR
 					(reg_q225 AND symb_decoder(16#4a#)) OR
 					(reg_q225 AND symb_decoder(16#49#)) OR
 					(reg_q225 AND symb_decoder(16#f4#)) OR
 					(reg_q225 AND symb_decoder(16#b3#)) OR
 					(reg_q225 AND symb_decoder(16#d9#)) OR
 					(reg_q225 AND symb_decoder(16#04#)) OR
 					(reg_q225 AND symb_decoder(16#f7#)) OR
 					(reg_q225 AND symb_decoder(16#96#)) OR
 					(reg_q225 AND symb_decoder(16#32#)) OR
 					(reg_q225 AND symb_decoder(16#8c#)) OR
 					(reg_q225 AND symb_decoder(16#65#)) OR
 					(reg_q225 AND symb_decoder(16#c6#)) OR
 					(reg_q225 AND symb_decoder(16#9a#)) OR
 					(reg_q225 AND symb_decoder(16#e4#)) OR
 					(reg_q225 AND symb_decoder(16#d2#)) OR
 					(reg_q225 AND symb_decoder(16#e0#)) OR
 					(reg_q225 AND symb_decoder(16#eb#)) OR
 					(reg_q225 AND symb_decoder(16#d1#)) OR
 					(reg_q225 AND symb_decoder(16#38#)) OR
 					(reg_q225 AND symb_decoder(16#fc#)) OR
 					(reg_q225 AND symb_decoder(16#63#)) OR
 					(reg_q225 AND symb_decoder(16#28#)) OR
 					(reg_q225 AND symb_decoder(16#93#)) OR
 					(reg_q225 AND symb_decoder(16#13#)) OR
 					(reg_q225 AND symb_decoder(16#23#)) OR
 					(reg_q225 AND symb_decoder(16#45#)) OR
 					(reg_q225 AND symb_decoder(16#4c#)) OR
 					(reg_q225 AND symb_decoder(16#00#)) OR
 					(reg_q225 AND symb_decoder(16#d0#)) OR
 					(reg_q225 AND symb_decoder(16#df#)) OR
 					(reg_q225 AND symb_decoder(16#e8#)) OR
 					(reg_q225 AND symb_decoder(16#a6#)) OR
 					(reg_q225 AND symb_decoder(16#06#)) OR
 					(reg_q225 AND symb_decoder(16#f5#)) OR
 					(reg_q225 AND symb_decoder(16#08#)) OR
 					(reg_q225 AND symb_decoder(16#09#)) OR
 					(reg_q225 AND symb_decoder(16#6e#)) OR
 					(reg_q225 AND symb_decoder(16#78#)) OR
 					(reg_q225 AND symb_decoder(16#83#)) OR
 					(reg_q225 AND symb_decoder(16#88#)) OR
 					(reg_q225 AND symb_decoder(16#29#)) OR
 					(reg_q225 AND symb_decoder(16#cb#)) OR
 					(reg_q225 AND symb_decoder(16#5b#)) OR
 					(reg_q225 AND symb_decoder(16#f3#)) OR
 					(reg_q225 AND symb_decoder(16#fb#)) OR
 					(reg_q225 AND symb_decoder(16#ec#)) OR
 					(reg_q225 AND symb_decoder(16#26#)) OR
 					(reg_q225 AND symb_decoder(16#5a#)) OR
 					(reg_q225 AND symb_decoder(16#15#)) OR
 					(reg_q225 AND symb_decoder(16#8d#)) OR
 					(reg_q225 AND symb_decoder(16#2b#)) OR
 					(reg_q225 AND symb_decoder(16#e9#)) OR
 					(reg_q225 AND symb_decoder(16#02#)) OR
 					(reg_q225 AND symb_decoder(16#1e#)) OR
 					(reg_q225 AND symb_decoder(16#ba#)) OR
 					(reg_q225 AND symb_decoder(16#31#)) OR
 					(reg_q225 AND symb_decoder(16#c2#)) OR
 					(reg_q225 AND symb_decoder(16#79#)) OR
 					(reg_q225 AND symb_decoder(16#a5#)) OR
 					(reg_q225 AND symb_decoder(16#f8#)) OR
 					(reg_q225 AND symb_decoder(16#43#)) OR
 					(reg_q225 AND symb_decoder(16#67#)) OR
 					(reg_q225 AND symb_decoder(16#ae#)) OR
 					(reg_q225 AND symb_decoder(16#e1#)) OR
 					(reg_q225 AND symb_decoder(16#ce#)) OR
 					(reg_q225 AND symb_decoder(16#57#)) OR
 					(reg_q225 AND symb_decoder(16#8f#)) OR
 					(reg_q225 AND symb_decoder(16#19#)) OR
 					(reg_q225 AND symb_decoder(16#c7#)) OR
 					(reg_q225 AND symb_decoder(16#c9#)) OR
 					(reg_q225 AND symb_decoder(16#9d#)) OR
 					(reg_q225 AND symb_decoder(16#7d#)) OR
 					(reg_q225 AND symb_decoder(16#da#)) OR
 					(reg_q225 AND symb_decoder(16#c4#)) OR
 					(reg_q225 AND symb_decoder(16#6a#)) OR
 					(reg_q225 AND symb_decoder(16#ff#)) OR
 					(reg_q225 AND symb_decoder(16#76#)) OR
 					(reg_q225 AND symb_decoder(16#cf#)) OR
 					(reg_q225 AND symb_decoder(16#9e#)) OR
 					(reg_q225 AND symb_decoder(16#6d#)) OR
 					(reg_q225 AND symb_decoder(16#24#)) OR
 					(reg_q225 AND symb_decoder(16#3f#)) OR
 					(reg_q225 AND symb_decoder(16#62#)) OR
 					(reg_q225 AND symb_decoder(16#27#)) OR
 					(reg_q225 AND symb_decoder(16#a9#)) OR
 					(reg_q225 AND symb_decoder(16#ca#)) OR
 					(reg_q225 AND symb_decoder(16#f6#)) OR
 					(reg_q225 AND symb_decoder(16#c1#)) OR
 					(reg_q225 AND symb_decoder(16#3e#)) OR
 					(reg_q225 AND symb_decoder(16#af#)) OR
 					(reg_q225 AND symb_decoder(16#1c#)) OR
 					(reg_q225 AND symb_decoder(16#bd#)) OR
 					(reg_q225 AND symb_decoder(16#7e#)) OR
 					(reg_q225 AND symb_decoder(16#f1#)) OR
 					(reg_q225 AND symb_decoder(16#97#)) OR
 					(reg_q225 AND symb_decoder(16#6f#)) OR
 					(reg_q225 AND symb_decoder(16#bc#)) OR
 					(reg_q225 AND symb_decoder(16#44#)) OR
 					(reg_q225 AND symb_decoder(16#37#)) OR
 					(reg_q225 AND symb_decoder(16#82#)) OR
 					(reg_q225 AND symb_decoder(16#5d#)) OR
 					(reg_q225 AND symb_decoder(16#47#)) OR
 					(reg_q225 AND symb_decoder(16#81#)) OR
 					(reg_q225 AND symb_decoder(16#9b#)) OR
 					(reg_q225 AND symb_decoder(16#2c#)) OR
 					(reg_q225 AND symb_decoder(16#5c#)) OR
 					(reg_q225 AND symb_decoder(16#74#)) OR
 					(reg_q225 AND symb_decoder(16#4e#)) OR
 					(reg_q225 AND symb_decoder(16#03#)) OR
 					(reg_q225 AND symb_decoder(16#7c#)) OR
 					(reg_q225 AND symb_decoder(16#0c#)) OR
 					(reg_q225 AND symb_decoder(16#c8#)) OR
 					(reg_q225 AND symb_decoder(16#11#)) OR
 					(reg_q225 AND symb_decoder(16#a2#)) OR
 					(reg_q225 AND symb_decoder(16#b2#)) OR
 					(reg_q225 AND symb_decoder(16#35#)) OR
 					(reg_q225 AND symb_decoder(16#98#)) OR
 					(reg_q225 AND symb_decoder(16#66#)) OR
 					(reg_q225 AND symb_decoder(16#39#)) OR
 					(reg_q225 AND symb_decoder(16#8a#)) OR
 					(reg_q225 AND symb_decoder(16#2a#)) OR
 					(reg_q225 AND symb_decoder(16#69#)) OR
 					(reg_q225 AND symb_decoder(16#b5#)) OR
 					(reg_q225 AND symb_decoder(16#16#)) OR
 					(reg_q225 AND symb_decoder(16#58#)) OR
 					(reg_q225 AND symb_decoder(16#a4#)) OR
 					(reg_q225 AND symb_decoder(16#be#)) OR
 					(reg_q225 AND symb_decoder(16#cc#)) OR
 					(reg_q225 AND symb_decoder(16#b7#)) OR
 					(reg_q225 AND symb_decoder(16#e3#)) OR
 					(reg_q225 AND symb_decoder(16#33#)) OR
 					(reg_q225 AND symb_decoder(16#25#)) OR
 					(reg_q225 AND symb_decoder(16#41#)) OR
 					(reg_q225 AND symb_decoder(16#80#)) OR
 					(reg_q225 AND symb_decoder(16#a1#)) OR
 					(reg_q225 AND symb_decoder(16#77#)) OR
 					(reg_q225 AND symb_decoder(16#9f#)) OR
 					(reg_q225 AND symb_decoder(16#ef#)) OR
 					(reg_q225 AND symb_decoder(16#7f#)) OR
 					(reg_q225 AND symb_decoder(16#ac#)) OR
 					(reg_q225 AND symb_decoder(16#2e#)) OR
 					(reg_q225 AND symb_decoder(16#b1#)) OR
 					(reg_q225 AND symb_decoder(16#1b#)) OR
 					(reg_q225 AND symb_decoder(16#12#)) OR
 					(reg_q225 AND symb_decoder(16#87#)) OR
 					(reg_q225 AND symb_decoder(16#3d#)) OR
 					(reg_q225 AND symb_decoder(16#40#)) OR
 					(reg_q225 AND symb_decoder(16#60#)) OR
 					(reg_q225 AND symb_decoder(16#e6#)) OR
 					(reg_q225 AND symb_decoder(16#5f#)) OR
 					(reg_q225 AND symb_decoder(16#a3#)) OR
 					(reg_q225 AND symb_decoder(16#52#)) OR
 					(reg_q225 AND symb_decoder(16#2f#)) OR
 					(reg_q225 AND symb_decoder(16#5e#)) OR
 					(reg_q225 AND symb_decoder(16#d6#)) OR
 					(reg_q225 AND symb_decoder(16#70#)) OR
 					(reg_q225 AND symb_decoder(16#bf#)) OR
 					(reg_q225 AND symb_decoder(16#21#)) OR
 					(reg_q225 AND symb_decoder(16#18#)) OR
 					(reg_q225 AND symb_decoder(16#d4#)) OR
 					(reg_q225 AND symb_decoder(16#fa#)) OR
 					(reg_q225 AND symb_decoder(16#22#)) OR
 					(reg_q225 AND symb_decoder(16#e7#)) OR
 					(reg_q225 AND symb_decoder(16#fe#)) OR
 					(reg_q225 AND symb_decoder(16#42#)) OR
 					(reg_q225 AND symb_decoder(16#89#)) OR
 					(reg_q225 AND symb_decoder(16#d7#)) OR
 					(reg_q225 AND symb_decoder(16#07#)) OR
 					(reg_q225 AND symb_decoder(16#de#)) OR
 					(reg_q225 AND symb_decoder(16#59#)) OR
 					(reg_q225 AND symb_decoder(16#ab#)) OR
 					(reg_q225 AND symb_decoder(16#1d#)) OR
 					(reg_q225 AND symb_decoder(16#50#)) OR
 					(reg_q225 AND symb_decoder(16#0b#)) OR
 					(reg_q225 AND symb_decoder(16#91#)) OR
 					(reg_q225 AND symb_decoder(16#10#)) OR
 					(reg_q225 AND symb_decoder(16#17#)) OR
 					(reg_q225 AND symb_decoder(16#c3#)) OR
 					(reg_q225 AND symb_decoder(16#73#)) OR
 					(reg_q225 AND symb_decoder(16#4d#)) OR
 					(reg_q225 AND symb_decoder(16#90#)) OR
 					(reg_q225 AND symb_decoder(16#b8#)) OR
 					(reg_q225 AND symb_decoder(16#7b#)) OR
 					(reg_q225 AND symb_decoder(16#4f#)) OR
 					(reg_q225 AND symb_decoder(16#ea#)) OR
 					(reg_q225 AND symb_decoder(16#f9#)) OR
 					(reg_q225 AND symb_decoder(16#8e#)) OR
 					(reg_q225 AND symb_decoder(16#68#)) OR
 					(reg_q225 AND symb_decoder(16#b9#)) OR
 					(reg_q225 AND symb_decoder(16#a0#)) OR
 					(reg_q225 AND symb_decoder(16#75#)) OR
 					(reg_q225 AND symb_decoder(16#b6#)) OR
 					(reg_q225 AND symb_decoder(16#61#));
reg_q225_init <= '0' ;
	p_reg_q225: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q225 <= reg_q225_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q225 <= reg_q225_init;
        else
          reg_q225 <= reg_q225_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1297_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1297 AND symb_decoder(16#24#)) OR
 					(reg_q1297 AND symb_decoder(16#64#)) OR
 					(reg_q1297 AND symb_decoder(16#eb#)) OR
 					(reg_q1297 AND symb_decoder(16#3a#)) OR
 					(reg_q1297 AND symb_decoder(16#45#)) OR
 					(reg_q1297 AND symb_decoder(16#01#)) OR
 					(reg_q1297 AND symb_decoder(16#d8#)) OR
 					(reg_q1297 AND symb_decoder(16#b2#)) OR
 					(reg_q1297 AND symb_decoder(16#6b#)) OR
 					(reg_q1297 AND symb_decoder(16#65#)) OR
 					(reg_q1297 AND symb_decoder(16#86#)) OR
 					(reg_q1297 AND symb_decoder(16#92#)) OR
 					(reg_q1297 AND symb_decoder(16#87#)) OR
 					(reg_q1297 AND symb_decoder(16#22#)) OR
 					(reg_q1297 AND symb_decoder(16#2a#)) OR
 					(reg_q1297 AND symb_decoder(16#55#)) OR
 					(reg_q1297 AND symb_decoder(16#13#)) OR
 					(reg_q1297 AND symb_decoder(16#e5#)) OR
 					(reg_q1297 AND symb_decoder(16#a3#)) OR
 					(reg_q1297 AND symb_decoder(16#12#)) OR
 					(reg_q1297 AND symb_decoder(16#8a#)) OR
 					(reg_q1297 AND symb_decoder(16#fd#)) OR
 					(reg_q1297 AND symb_decoder(16#41#)) OR
 					(reg_q1297 AND symb_decoder(16#08#)) OR
 					(reg_q1297 AND symb_decoder(16#71#)) OR
 					(reg_q1297 AND symb_decoder(16#4a#)) OR
 					(reg_q1297 AND symb_decoder(16#9d#)) OR
 					(reg_q1297 AND symb_decoder(16#3c#)) OR
 					(reg_q1297 AND symb_decoder(16#70#)) OR
 					(reg_q1297 AND symb_decoder(16#7e#)) OR
 					(reg_q1297 AND symb_decoder(16#69#)) OR
 					(reg_q1297 AND symb_decoder(16#80#)) OR
 					(reg_q1297 AND symb_decoder(16#78#)) OR
 					(reg_q1297 AND symb_decoder(16#06#)) OR
 					(reg_q1297 AND symb_decoder(16#19#)) OR
 					(reg_q1297 AND symb_decoder(16#2f#)) OR
 					(reg_q1297 AND symb_decoder(16#59#)) OR
 					(reg_q1297 AND symb_decoder(16#fe#)) OR
 					(reg_q1297 AND symb_decoder(16#e4#)) OR
 					(reg_q1297 AND symb_decoder(16#91#)) OR
 					(reg_q1297 AND symb_decoder(16#6c#)) OR
 					(reg_q1297 AND symb_decoder(16#2e#)) OR
 					(reg_q1297 AND symb_decoder(16#99#)) OR
 					(reg_q1297 AND symb_decoder(16#a2#)) OR
 					(reg_q1297 AND symb_decoder(16#94#)) OR
 					(reg_q1297 AND symb_decoder(16#21#)) OR
 					(reg_q1297 AND symb_decoder(16#8b#)) OR
 					(reg_q1297 AND symb_decoder(16#74#)) OR
 					(reg_q1297 AND symb_decoder(16#e7#)) OR
 					(reg_q1297 AND symb_decoder(16#6f#)) OR
 					(reg_q1297 AND symb_decoder(16#fa#)) OR
 					(reg_q1297 AND symb_decoder(16#a8#)) OR
 					(reg_q1297 AND symb_decoder(16#57#)) OR
 					(reg_q1297 AND symb_decoder(16#f6#)) OR
 					(reg_q1297 AND symb_decoder(16#f2#)) OR
 					(reg_q1297 AND symb_decoder(16#d5#)) OR
 					(reg_q1297 AND symb_decoder(16#35#)) OR
 					(reg_q1297 AND symb_decoder(16#43#)) OR
 					(reg_q1297 AND symb_decoder(16#51#)) OR
 					(reg_q1297 AND symb_decoder(16#27#)) OR
 					(reg_q1297 AND symb_decoder(16#18#)) OR
 					(reg_q1297 AND symb_decoder(16#a4#)) OR
 					(reg_q1297 AND symb_decoder(16#0d#)) OR
 					(reg_q1297 AND symb_decoder(16#b1#)) OR
 					(reg_q1297 AND symb_decoder(16#85#)) OR
 					(reg_q1297 AND symb_decoder(16#33#)) OR
 					(reg_q1297 AND symb_decoder(16#b3#)) OR
 					(reg_q1297 AND symb_decoder(16#11#)) OR
 					(reg_q1297 AND symb_decoder(16#98#)) OR
 					(reg_q1297 AND symb_decoder(16#e2#)) OR
 					(reg_q1297 AND symb_decoder(16#cc#)) OR
 					(reg_q1297 AND symb_decoder(16#32#)) OR
 					(reg_q1297 AND symb_decoder(16#ef#)) OR
 					(reg_q1297 AND symb_decoder(16#14#)) OR
 					(reg_q1297 AND symb_decoder(16#c0#)) OR
 					(reg_q1297 AND symb_decoder(16#d6#)) OR
 					(reg_q1297 AND symb_decoder(16#77#)) OR
 					(reg_q1297 AND symb_decoder(16#44#)) OR
 					(reg_q1297 AND symb_decoder(16#7c#)) OR
 					(reg_q1297 AND symb_decoder(16#e8#)) OR
 					(reg_q1297 AND symb_decoder(16#e1#)) OR
 					(reg_q1297 AND symb_decoder(16#31#)) OR
 					(reg_q1297 AND symb_decoder(16#b0#)) OR
 					(reg_q1297 AND symb_decoder(16#96#)) OR
 					(reg_q1297 AND symb_decoder(16#1b#)) OR
 					(reg_q1297 AND symb_decoder(16#4c#)) OR
 					(reg_q1297 AND symb_decoder(16#34#)) OR
 					(reg_q1297 AND symb_decoder(16#bc#)) OR
 					(reg_q1297 AND symb_decoder(16#a1#)) OR
 					(reg_q1297 AND symb_decoder(16#2b#)) OR
 					(reg_q1297 AND symb_decoder(16#ee#)) OR
 					(reg_q1297 AND symb_decoder(16#f1#)) OR
 					(reg_q1297 AND symb_decoder(16#56#)) OR
 					(reg_q1297 AND symb_decoder(16#50#)) OR
 					(reg_q1297 AND symb_decoder(16#5a#)) OR
 					(reg_q1297 AND symb_decoder(16#81#)) OR
 					(reg_q1297 AND symb_decoder(16#10#)) OR
 					(reg_q1297 AND symb_decoder(16#a7#)) OR
 					(reg_q1297 AND symb_decoder(16#ca#)) OR
 					(reg_q1297 AND symb_decoder(16#ed#)) OR
 					(reg_q1297 AND symb_decoder(16#8c#)) OR
 					(reg_q1297 AND symb_decoder(16#c5#)) OR
 					(reg_q1297 AND symb_decoder(16#b9#)) OR
 					(reg_q1297 AND symb_decoder(16#d3#)) OR
 					(reg_q1297 AND symb_decoder(16#6d#)) OR
 					(reg_q1297 AND symb_decoder(16#a6#)) OR
 					(reg_q1297 AND symb_decoder(16#4f#)) OR
 					(reg_q1297 AND symb_decoder(16#09#)) OR
 					(reg_q1297 AND symb_decoder(16#bb#)) OR
 					(reg_q1297 AND symb_decoder(16#26#)) OR
 					(reg_q1297 AND symb_decoder(16#da#)) OR
 					(reg_q1297 AND symb_decoder(16#9e#)) OR
 					(reg_q1297 AND symb_decoder(16#3b#)) OR
 					(reg_q1297 AND symb_decoder(16#fc#)) OR
 					(reg_q1297 AND symb_decoder(16#47#)) OR
 					(reg_q1297 AND symb_decoder(16#63#)) OR
 					(reg_q1297 AND symb_decoder(16#e6#)) OR
 					(reg_q1297 AND symb_decoder(16#4d#)) OR
 					(reg_q1297 AND symb_decoder(16#16#)) OR
 					(reg_q1297 AND symb_decoder(16#c9#)) OR
 					(reg_q1297 AND symb_decoder(16#be#)) OR
 					(reg_q1297 AND symb_decoder(16#ba#)) OR
 					(reg_q1297 AND symb_decoder(16#e0#)) OR
 					(reg_q1297 AND symb_decoder(16#76#)) OR
 					(reg_q1297 AND symb_decoder(16#9f#)) OR
 					(reg_q1297 AND symb_decoder(16#39#)) OR
 					(reg_q1297 AND symb_decoder(16#0a#)) OR
 					(reg_q1297 AND symb_decoder(16#c3#)) OR
 					(reg_q1297 AND symb_decoder(16#2d#)) OR
 					(reg_q1297 AND symb_decoder(16#c7#)) OR
 					(reg_q1297 AND symb_decoder(16#1f#)) OR
 					(reg_q1297 AND symb_decoder(16#1c#)) OR
 					(reg_q1297 AND symb_decoder(16#2c#)) OR
 					(reg_q1297 AND symb_decoder(16#88#)) OR
 					(reg_q1297 AND symb_decoder(16#6e#)) OR
 					(reg_q1297 AND symb_decoder(16#c1#)) OR
 					(reg_q1297 AND symb_decoder(16#db#)) OR
 					(reg_q1297 AND symb_decoder(16#ff#)) OR
 					(reg_q1297 AND symb_decoder(16#c6#)) OR
 					(reg_q1297 AND symb_decoder(16#a5#)) OR
 					(reg_q1297 AND symb_decoder(16#f3#)) OR
 					(reg_q1297 AND symb_decoder(16#f4#)) OR
 					(reg_q1297 AND symb_decoder(16#f5#)) OR
 					(reg_q1297 AND symb_decoder(16#f7#)) OR
 					(reg_q1297 AND symb_decoder(16#1e#)) OR
 					(reg_q1297 AND symb_decoder(16#00#)) OR
 					(reg_q1297 AND symb_decoder(16#b5#)) OR
 					(reg_q1297 AND symb_decoder(16#17#)) OR
 					(reg_q1297 AND symb_decoder(16#ec#)) OR
 					(reg_q1297 AND symb_decoder(16#1d#)) OR
 					(reg_q1297 AND symb_decoder(16#82#)) OR
 					(reg_q1297 AND symb_decoder(16#9c#)) OR
 					(reg_q1297 AND symb_decoder(16#bd#)) OR
 					(reg_q1297 AND symb_decoder(16#b8#)) OR
 					(reg_q1297 AND symb_decoder(16#c8#)) OR
 					(reg_q1297 AND symb_decoder(16#67#)) OR
 					(reg_q1297 AND symb_decoder(16#4b#)) OR
 					(reg_q1297 AND symb_decoder(16#30#)) OR
 					(reg_q1297 AND symb_decoder(16#20#)) OR
 					(reg_q1297 AND symb_decoder(16#fb#)) OR
 					(reg_q1297 AND symb_decoder(16#f0#)) OR
 					(reg_q1297 AND symb_decoder(16#1a#)) OR
 					(reg_q1297 AND symb_decoder(16#4e#)) OR
 					(reg_q1297 AND symb_decoder(16#b7#)) OR
 					(reg_q1297 AND symb_decoder(16#9a#)) OR
 					(reg_q1297 AND symb_decoder(16#ac#)) OR
 					(reg_q1297 AND symb_decoder(16#83#)) OR
 					(reg_q1297 AND symb_decoder(16#48#)) OR
 					(reg_q1297 AND symb_decoder(16#8d#)) OR
 					(reg_q1297 AND symb_decoder(16#29#)) OR
 					(reg_q1297 AND symb_decoder(16#97#)) OR
 					(reg_q1297 AND symb_decoder(16#23#)) OR
 					(reg_q1297 AND symb_decoder(16#d2#)) OR
 					(reg_q1297 AND symb_decoder(16#5e#)) OR
 					(reg_q1297 AND symb_decoder(16#0b#)) OR
 					(reg_q1297 AND symb_decoder(16#b4#)) OR
 					(reg_q1297 AND symb_decoder(16#8f#)) OR
 					(reg_q1297 AND symb_decoder(16#15#)) OR
 					(reg_q1297 AND symb_decoder(16#dd#)) OR
 					(reg_q1297 AND symb_decoder(16#03#)) OR
 					(reg_q1297 AND symb_decoder(16#62#)) OR
 					(reg_q1297 AND symb_decoder(16#42#)) OR
 					(reg_q1297 AND symb_decoder(16#58#)) OR
 					(reg_q1297 AND symb_decoder(16#3d#)) OR
 					(reg_q1297 AND symb_decoder(16#6a#)) OR
 					(reg_q1297 AND symb_decoder(16#61#)) OR
 					(reg_q1297 AND symb_decoder(16#cf#)) OR
 					(reg_q1297 AND symb_decoder(16#f9#)) OR
 					(reg_q1297 AND symb_decoder(16#d1#)) OR
 					(reg_q1297 AND symb_decoder(16#a9#)) OR
 					(reg_q1297 AND symb_decoder(16#f8#)) OR
 					(reg_q1297 AND symb_decoder(16#c4#)) OR
 					(reg_q1297 AND symb_decoder(16#ad#)) OR
 					(reg_q1297 AND symb_decoder(16#b6#)) OR
 					(reg_q1297 AND symb_decoder(16#72#)) OR
 					(reg_q1297 AND symb_decoder(16#40#)) OR
 					(reg_q1297 AND symb_decoder(16#84#)) OR
 					(reg_q1297 AND symb_decoder(16#02#)) OR
 					(reg_q1297 AND symb_decoder(16#ea#)) OR
 					(reg_q1297 AND symb_decoder(16#c2#)) OR
 					(reg_q1297 AND symb_decoder(16#53#)) OR
 					(reg_q1297 AND symb_decoder(16#5b#)) OR
 					(reg_q1297 AND symb_decoder(16#75#)) OR
 					(reg_q1297 AND symb_decoder(16#df#)) OR
 					(reg_q1297 AND symb_decoder(16#0f#)) OR
 					(reg_q1297 AND symb_decoder(16#bf#)) OR
 					(reg_q1297 AND symb_decoder(16#28#)) OR
 					(reg_q1297 AND symb_decoder(16#0c#)) OR
 					(reg_q1297 AND symb_decoder(16#49#)) OR
 					(reg_q1297 AND symb_decoder(16#68#)) OR
 					(reg_q1297 AND symb_decoder(16#ce#)) OR
 					(reg_q1297 AND symb_decoder(16#3f#)) OR
 					(reg_q1297 AND symb_decoder(16#25#)) OR
 					(reg_q1297 AND symb_decoder(16#04#)) OR
 					(reg_q1297 AND symb_decoder(16#93#)) OR
 					(reg_q1297 AND symb_decoder(16#52#)) OR
 					(reg_q1297 AND symb_decoder(16#d0#)) OR
 					(reg_q1297 AND symb_decoder(16#37#)) OR
 					(reg_q1297 AND symb_decoder(16#89#)) OR
 					(reg_q1297 AND symb_decoder(16#7f#)) OR
 					(reg_q1297 AND symb_decoder(16#de#)) OR
 					(reg_q1297 AND symb_decoder(16#0e#)) OR
 					(reg_q1297 AND symb_decoder(16#36#)) OR
 					(reg_q1297 AND symb_decoder(16#54#)) OR
 					(reg_q1297 AND symb_decoder(16#cd#)) OR
 					(reg_q1297 AND symb_decoder(16#46#)) OR
 					(reg_q1297 AND symb_decoder(16#79#)) OR
 					(reg_q1297 AND symb_decoder(16#9b#)) OR
 					(reg_q1297 AND symb_decoder(16#dc#)) OR
 					(reg_q1297 AND symb_decoder(16#d9#)) OR
 					(reg_q1297 AND symb_decoder(16#3e#)) OR
 					(reg_q1297 AND symb_decoder(16#aa#)) OR
 					(reg_q1297 AND symb_decoder(16#7b#)) OR
 					(reg_q1297 AND symb_decoder(16#5c#)) OR
 					(reg_q1297 AND symb_decoder(16#60#)) OR
 					(reg_q1297 AND symb_decoder(16#e3#)) OR
 					(reg_q1297 AND symb_decoder(16#38#)) OR
 					(reg_q1297 AND symb_decoder(16#95#)) OR
 					(reg_q1297 AND symb_decoder(16#05#)) OR
 					(reg_q1297 AND symb_decoder(16#a0#)) OR
 					(reg_q1297 AND symb_decoder(16#8e#)) OR
 					(reg_q1297 AND symb_decoder(16#7d#)) OR
 					(reg_q1297 AND symb_decoder(16#73#)) OR
 					(reg_q1297 AND symb_decoder(16#7a#)) OR
 					(reg_q1297 AND symb_decoder(16#5d#)) OR
 					(reg_q1297 AND symb_decoder(16#5f#)) OR
 					(reg_q1297 AND symb_decoder(16#ab#)) OR
 					(reg_q1297 AND symb_decoder(16#66#)) OR
 					(reg_q1297 AND symb_decoder(16#d7#)) OR
 					(reg_q1297 AND symb_decoder(16#d4#)) OR
 					(reg_q1297 AND symb_decoder(16#90#)) OR
 					(reg_q1297 AND symb_decoder(16#af#)) OR
 					(reg_q1297 AND symb_decoder(16#e9#)) OR
 					(reg_q1297 AND symb_decoder(16#ae#)) OR
 					(reg_q1297 AND symb_decoder(16#07#)) OR
 					(reg_q1297 AND symb_decoder(16#cb#));
reg_q1297_init <= '0' ;
	p_reg_q1297: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1297 <= reg_q1297_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1297 <= reg_q1297_init;
        else
          reg_q1297 <= reg_q1297_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph7

reg_q1876_in <= (reg_q1874 AND symb_decoder(16#54#)) OR
 					(reg_q1874 AND symb_decoder(16#74#));
reg_q1878_in <= (reg_q1876 AND symb_decoder(16#61#)) OR
 					(reg_q1876 AND symb_decoder(16#41#));
reg_q1792_in <= (reg_q1790 AND symb_decoder(16#69#)) OR
 					(reg_q1790 AND symb_decoder(16#49#));
reg_q1794_in <= (reg_q1792 AND symb_decoder(16#4d#)) OR
 					(reg_q1792 AND symb_decoder(16#6d#));
reg_q1852_in <= (reg_q1850 AND symb_decoder(16#65#)) OR
 					(reg_q1850 AND symb_decoder(16#45#));
reg_q1854_in <= (reg_q1852 AND symb_decoder(16#72#)) OR
 					(reg_q1852 AND symb_decoder(16#52#));
reg_q889_in <= (reg_q887 AND symb_decoder(16#5b#));
reg_q532_in <= (reg_q530 AND symb_decoder(16#2e#));
reg_q534_in <= (reg_q532 AND symb_decoder(16#39#)) OR
 					(reg_q532 AND symb_decoder(16#35#)) OR
 					(reg_q532 AND symb_decoder(16#30#)) OR
 					(reg_q532 AND symb_decoder(16#33#)) OR
 					(reg_q532 AND symb_decoder(16#38#)) OR
 					(reg_q532 AND symb_decoder(16#36#)) OR
 					(reg_q532 AND symb_decoder(16#37#)) OR
 					(reg_q532 AND symb_decoder(16#34#)) OR
 					(reg_q532 AND symb_decoder(16#31#)) OR
 					(reg_q532 AND symb_decoder(16#32#)) OR
 					(reg_q534 AND symb_decoder(16#32#)) OR
 					(reg_q534 AND symb_decoder(16#34#)) OR
 					(reg_q534 AND symb_decoder(16#36#)) OR
 					(reg_q534 AND symb_decoder(16#38#)) OR
 					(reg_q534 AND symb_decoder(16#33#)) OR
 					(reg_q534 AND symb_decoder(16#35#)) OR
 					(reg_q534 AND symb_decoder(16#37#)) OR
 					(reg_q534 AND symb_decoder(16#31#)) OR
 					(reg_q534 AND symb_decoder(16#30#)) OR
 					(reg_q534 AND symb_decoder(16#39#));
reg_q2419_in <= (reg_q2417 AND symb_decoder(16#45#)) OR
 					(reg_q2417 AND symb_decoder(16#65#));
reg_q2421_in <= (reg_q2419 AND symb_decoder(16#73#)) OR
 					(reg_q2419 AND symb_decoder(16#53#));
reg_q1770_in <= (reg_q1768 AND symb_decoder(16#0a#)) OR
 					(reg_q1768 AND symb_decoder(16#20#)) OR
 					(reg_q1768 AND symb_decoder(16#0c#)) OR
 					(reg_q1768 AND symb_decoder(16#09#)) OR
 					(reg_q1768 AND symb_decoder(16#0d#));
reg_q616_in <= (reg_q616 AND symb_decoder(16#31#)) OR
 					(reg_q616 AND symb_decoder(16#35#)) OR
 					(reg_q616 AND symb_decoder(16#30#)) OR
 					(reg_q616 AND symb_decoder(16#32#)) OR
 					(reg_q616 AND symb_decoder(16#38#)) OR
 					(reg_q616 AND symb_decoder(16#33#)) OR
 					(reg_q616 AND symb_decoder(16#37#)) OR
 					(reg_q616 AND symb_decoder(16#39#)) OR
 					(reg_q616 AND symb_decoder(16#34#)) OR
 					(reg_q616 AND symb_decoder(16#36#)) OR
 					(reg_q614 AND symb_decoder(16#30#)) OR
 					(reg_q614 AND symb_decoder(16#31#)) OR
 					(reg_q614 AND symb_decoder(16#36#)) OR
 					(reg_q614 AND symb_decoder(16#35#)) OR
 					(reg_q614 AND symb_decoder(16#33#)) OR
 					(reg_q614 AND symb_decoder(16#38#)) OR
 					(reg_q614 AND symb_decoder(16#34#)) OR
 					(reg_q614 AND symb_decoder(16#32#)) OR
 					(reg_q614 AND symb_decoder(16#39#)) OR
 					(reg_q614 AND symb_decoder(16#37#));
reg_q526_in <= (reg_q526 AND symb_decoder(16#37#)) OR
 					(reg_q526 AND symb_decoder(16#39#)) OR
 					(reg_q526 AND symb_decoder(16#36#)) OR
 					(reg_q526 AND symb_decoder(16#31#)) OR
 					(reg_q526 AND symb_decoder(16#35#)) OR
 					(reg_q526 AND symb_decoder(16#30#)) OR
 					(reg_q526 AND symb_decoder(16#33#)) OR
 					(reg_q526 AND symb_decoder(16#32#)) OR
 					(reg_q526 AND symb_decoder(16#34#)) OR
 					(reg_q526 AND symb_decoder(16#38#)) OR
 					(reg_q524 AND symb_decoder(16#30#)) OR
 					(reg_q524 AND symb_decoder(16#39#)) OR
 					(reg_q524 AND symb_decoder(16#31#)) OR
 					(reg_q524 AND symb_decoder(16#36#)) OR
 					(reg_q524 AND symb_decoder(16#32#)) OR
 					(reg_q524 AND symb_decoder(16#34#)) OR
 					(reg_q524 AND symb_decoder(16#37#)) OR
 					(reg_q524 AND symb_decoder(16#38#)) OR
 					(reg_q524 AND symb_decoder(16#33#)) OR
 					(reg_q524 AND symb_decoder(16#35#));
reg_q945_in <= (reg_q943 AND symb_decoder(16#2e#));
reg_q947_in <= (reg_q945 AND symb_decoder(16#33#)) OR
 					(reg_q945 AND symb_decoder(16#36#)) OR
 					(reg_q945 AND symb_decoder(16#37#)) OR
 					(reg_q945 AND symb_decoder(16#30#)) OR
 					(reg_q945 AND symb_decoder(16#31#)) OR
 					(reg_q945 AND symb_decoder(16#34#)) OR
 					(reg_q945 AND symb_decoder(16#38#)) OR
 					(reg_q945 AND symb_decoder(16#32#)) OR
 					(reg_q945 AND symb_decoder(16#35#)) OR
 					(reg_q945 AND symb_decoder(16#39#)) OR
 					(reg_q947 AND symb_decoder(16#31#)) OR
 					(reg_q947 AND symb_decoder(16#34#)) OR
 					(reg_q947 AND symb_decoder(16#36#)) OR
 					(reg_q947 AND symb_decoder(16#38#)) OR
 					(reg_q947 AND symb_decoder(16#30#)) OR
 					(reg_q947 AND symb_decoder(16#33#)) OR
 					(reg_q947 AND symb_decoder(16#39#)) OR
 					(reg_q947 AND symb_decoder(16#37#)) OR
 					(reg_q947 AND symb_decoder(16#32#)) OR
 					(reg_q947 AND symb_decoder(16#35#));
reg_q791_in <= (reg_q789 AND symb_decoder(16#5e#));
reg_q856_in <= (reg_q854 AND symb_decoder(16#72#)) OR
 					(reg_q854 AND symb_decoder(16#52#));
reg_q858_in <= (reg_q856 AND symb_decoder(16#49#)) OR
 					(reg_q856 AND symb_decoder(16#69#));
reg_q1215_in <= (reg_q1213 AND symb_decoder(16#4d#)) OR
 					(reg_q1213 AND symb_decoder(16#6d#));
reg_q1217_in <= (reg_q1215 AND symb_decoder(16#45#)) OR
 					(reg_q1215 AND symb_decoder(16#65#));
reg_q937_in <= (reg_q955 AND symb_decoder(16#00#)) OR
 					(reg_q933 AND symb_decoder(16#00#));
reg_q939_in <= (reg_q937 AND symb_decoder(16#33#)) OR
 					(reg_q937 AND symb_decoder(16#31#)) OR
 					(reg_q937 AND symb_decoder(16#39#)) OR
 					(reg_q937 AND symb_decoder(16#32#)) OR
 					(reg_q937 AND symb_decoder(16#37#)) OR
 					(reg_q937 AND symb_decoder(16#30#)) OR
 					(reg_q937 AND symb_decoder(16#34#)) OR
 					(reg_q937 AND symb_decoder(16#36#)) OR
 					(reg_q937 AND symb_decoder(16#35#)) OR
 					(reg_q937 AND symb_decoder(16#38#)) OR
 					(reg_q939 AND symb_decoder(16#39#)) OR
 					(reg_q939 AND symb_decoder(16#35#)) OR
 					(reg_q939 AND symb_decoder(16#32#)) OR
 					(reg_q939 AND symb_decoder(16#34#)) OR
 					(reg_q939 AND symb_decoder(16#36#)) OR
 					(reg_q939 AND symb_decoder(16#31#)) OR
 					(reg_q939 AND symb_decoder(16#33#)) OR
 					(reg_q939 AND symb_decoder(16#38#)) OR
 					(reg_q939 AND symb_decoder(16#37#)) OR
 					(reg_q939 AND symb_decoder(16#30#));
reg_q1866_in <= (reg_q1864 AND symb_decoder(16#2e#));
reg_q2002_in <= (reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2001 AND symb_decoder(16#54#)) OR
 					(reg_q2001 AND symb_decoder(16#74#));
reg_q520_in <= (reg_q518 AND symb_decoder(16#5f#));
reg_q522_in <= (reg_q520 AND symb_decoder(16#39#)) OR
 					(reg_q520 AND symb_decoder(16#30#)) OR
 					(reg_q520 AND symb_decoder(16#37#)) OR
 					(reg_q520 AND symb_decoder(16#32#)) OR
 					(reg_q520 AND symb_decoder(16#31#)) OR
 					(reg_q520 AND symb_decoder(16#33#)) OR
 					(reg_q520 AND symb_decoder(16#34#)) OR
 					(reg_q520 AND symb_decoder(16#35#)) OR
 					(reg_q520 AND symb_decoder(16#36#)) OR
 					(reg_q520 AND symb_decoder(16#38#)) OR
 					(reg_q522 AND symb_decoder(16#32#)) OR
 					(reg_q522 AND symb_decoder(16#31#)) OR
 					(reg_q522 AND symb_decoder(16#35#)) OR
 					(reg_q522 AND symb_decoder(16#34#)) OR
 					(reg_q522 AND symb_decoder(16#37#)) OR
 					(reg_q522 AND symb_decoder(16#39#)) OR
 					(reg_q522 AND symb_decoder(16#36#)) OR
 					(reg_q522 AND symb_decoder(16#38#)) OR
 					(reg_q522 AND symb_decoder(16#30#)) OR
 					(reg_q522 AND symb_decoder(16#33#));
reg_q2528_in <= (reg_q2526 AND symb_decoder(16#3b#));
reg_q2530_in <= (reg_q2528 AND symb_decoder(16#31#)) OR
 					(reg_q2528 AND symb_decoder(16#32#)) OR
 					(reg_q2528 AND symb_decoder(16#34#)) OR
 					(reg_q2528 AND symb_decoder(16#33#)) OR
 					(reg_q2528 AND symb_decoder(16#36#)) OR
 					(reg_q2528 AND symb_decoder(16#38#)) OR
 					(reg_q2528 AND symb_decoder(16#30#)) OR
 					(reg_q2528 AND symb_decoder(16#35#)) OR
 					(reg_q2528 AND symb_decoder(16#39#)) OR
 					(reg_q2528 AND symb_decoder(16#37#)) OR
 					(reg_q2530 AND symb_decoder(16#32#)) OR
 					(reg_q2530 AND symb_decoder(16#35#)) OR
 					(reg_q2530 AND symb_decoder(16#39#)) OR
 					(reg_q2530 AND symb_decoder(16#37#)) OR
 					(reg_q2530 AND symb_decoder(16#36#)) OR
 					(reg_q2530 AND symb_decoder(16#34#)) OR
 					(reg_q2530 AND symb_decoder(16#31#)) OR
 					(reg_q2530 AND symb_decoder(16#33#)) OR
 					(reg_q2530 AND symb_decoder(16#38#)) OR
 					(reg_q2530 AND symb_decoder(16#30#));
reg_q2445_in <= (reg_q2443 AND symb_decoder(16#6f#)) OR
 					(reg_q2443 AND symb_decoder(16#4f#));
reg_q2447_in <= (reg_q2445 AND symb_decoder(16#61#)) OR
 					(reg_q2445 AND symb_decoder(16#41#));
reg_q1874_in <= (reg_q1872 AND symb_decoder(16#52#)) OR
 					(reg_q1872 AND symb_decoder(16#72#));
reg_q2078_in <= (reg_q2076 AND symb_decoder(16#65#));
reg_q2080_in <= (reg_q2078 AND symb_decoder(16#72#));
reg_q2178_in <= (reg_q2176 AND symb_decoder(16#69#)) OR
 					(reg_q2176 AND symb_decoder(16#49#));
reg_q2180_in <= (reg_q2178 AND symb_decoder(16#43#)) OR
 					(reg_q2178 AND symb_decoder(16#63#));
reg_q590_in <= (reg_q588 AND symb_decoder(16#54#)) OR
 					(reg_q588 AND symb_decoder(16#74#));
reg_q592_in <= (reg_q590 AND symb_decoder(16#69#)) OR
 					(reg_q590 AND symb_decoder(16#49#));
reg_q1387_in <= (reg_q1385 AND symb_decoder(16#41#)) OR
 					(reg_q1385 AND symb_decoder(16#61#));
reg_q1389_in <= (reg_q1387 AND symb_decoder(16#4d#)) OR
 					(reg_q1387 AND symb_decoder(16#6d#));
reg_q2405_in <= (reg_q2403 AND symb_decoder(16#62#)) OR
 					(reg_q2403 AND symb_decoder(16#42#));
reg_q2407_in <= (reg_q2405 AND symb_decoder(16#61#)) OR
 					(reg_q2405 AND symb_decoder(16#41#));
reg_q1920_in <= (reg_q1918 AND symb_decoder(16#57#)) OR
 					(reg_q1918 AND symb_decoder(16#77#));
reg_q1409_in <= (reg_q1407 AND symb_decoder(16#41#)) OR
 					(reg_q1407 AND symb_decoder(16#61#));
reg_q1411_in <= (reg_q1409 AND symb_decoder(16#6b#)) OR
 					(reg_q1409 AND symb_decoder(16#4b#));
reg_q2064_in <= (reg_q2062 AND symb_decoder(16#32#));
reg_q960_in <= (reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q960 AND symb_decoder(16#35#)) OR
 					(reg_q960 AND symb_decoder(16#37#)) OR
 					(reg_q960 AND symb_decoder(16#38#)) OR
 					(reg_q960 AND symb_decoder(16#30#)) OR
 					(reg_q960 AND symb_decoder(16#36#)) OR
 					(reg_q960 AND symb_decoder(16#39#)) OR
 					(reg_q960 AND symb_decoder(16#32#)) OR
 					(reg_q960 AND symb_decoder(16#33#)) OR
 					(reg_q960 AND symb_decoder(16#34#)) OR
 					(reg_q960 AND symb_decoder(16#31#)) OR
 					(reg_q959 AND symb_decoder(16#37#)) OR
 					(reg_q959 AND symb_decoder(16#31#)) OR
 					(reg_q959 AND symb_decoder(16#33#)) OR
 					(reg_q959 AND symb_decoder(16#32#)) OR
 					(reg_q959 AND symb_decoder(16#30#)) OR
 					(reg_q959 AND symb_decoder(16#35#)) OR
 					(reg_q959 AND symb_decoder(16#38#)) OR
 					(reg_q959 AND symb_decoder(16#34#)) OR
 					(reg_q959 AND symb_decoder(16#39#)) OR
 					(reg_q959 AND symb_decoder(16#36#));
reg_q874_in <= (reg_q872 AND symb_decoder(16#5c#));
reg_q876_in <= (reg_q874 AND symb_decoder(16#5d#));
reg_q949_in <= (reg_q947 AND symb_decoder(16#2e#));
reg_q951_in <= (reg_q949 AND symb_decoder(16#35#)) OR
 					(reg_q949 AND symb_decoder(16#31#)) OR
 					(reg_q949 AND symb_decoder(16#34#)) OR
 					(reg_q949 AND symb_decoder(16#36#)) OR
 					(reg_q949 AND symb_decoder(16#33#)) OR
 					(reg_q949 AND symb_decoder(16#38#)) OR
 					(reg_q949 AND symb_decoder(16#32#)) OR
 					(reg_q949 AND symb_decoder(16#39#)) OR
 					(reg_q949 AND symb_decoder(16#30#)) OR
 					(reg_q949 AND symb_decoder(16#37#)) OR
 					(reg_q951 AND symb_decoder(16#39#)) OR
 					(reg_q951 AND symb_decoder(16#33#)) OR
 					(reg_q951 AND symb_decoder(16#32#)) OR
 					(reg_q951 AND symb_decoder(16#34#)) OR
 					(reg_q951 AND symb_decoder(16#37#)) OR
 					(reg_q951 AND symb_decoder(16#35#)) OR
 					(reg_q951 AND symb_decoder(16#38#)) OR
 					(reg_q951 AND symb_decoder(16#36#)) OR
 					(reg_q951 AND symb_decoder(16#31#)) OR
 					(reg_q951 AND symb_decoder(16#30#));
reg_q12_in <= (reg_q10 AND symb_decoder(16#6c#)) OR
 					(reg_q10 AND symb_decoder(16#4c#));
reg_q2409_in <= (reg_q2407 AND symb_decoder(16#72#)) OR
 					(reg_q2407 AND symb_decoder(16#52#));
reg_q882_in <= (reg_q880 AND symb_decoder(16#4d#)) OR
 					(reg_q880 AND symb_decoder(16#6b#)) OR
 					(reg_q880 AND symb_decoder(16#54#)) OR
 					(reg_q880 AND symb_decoder(16#62#)) OR
 					(reg_q880 AND symb_decoder(16#46#)) OR
 					(reg_q880 AND symb_decoder(16#4e#)) OR
 					(reg_q880 AND symb_decoder(16#51#)) OR
 					(reg_q880 AND symb_decoder(16#71#)) OR
 					(reg_q880 AND symb_decoder(16#67#)) OR
 					(reg_q880 AND symb_decoder(16#55#)) OR
 					(reg_q880 AND symb_decoder(16#50#)) OR
 					(reg_q880 AND symb_decoder(16#7a#)) OR
 					(reg_q880 AND symb_decoder(16#56#)) OR
 					(reg_q880 AND symb_decoder(16#70#)) OR
 					(reg_q880 AND symb_decoder(16#4f#)) OR
 					(reg_q880 AND symb_decoder(16#69#)) OR
 					(reg_q880 AND symb_decoder(16#58#)) OR
 					(reg_q880 AND symb_decoder(16#5a#)) OR
 					(reg_q880 AND symb_decoder(16#6a#)) OR
 					(reg_q880 AND symb_decoder(16#73#)) OR
 					(reg_q880 AND symb_decoder(16#41#)) OR
 					(reg_q880 AND symb_decoder(16#76#)) OR
 					(reg_q880 AND symb_decoder(16#77#)) OR
 					(reg_q880 AND symb_decoder(16#6c#)) OR
 					(reg_q880 AND symb_decoder(16#59#)) OR
 					(reg_q880 AND symb_decoder(16#6f#)) OR
 					(reg_q880 AND symb_decoder(16#45#)) OR
 					(reg_q880 AND symb_decoder(16#68#)) OR
 					(reg_q880 AND symb_decoder(16#6d#)) OR
 					(reg_q880 AND symb_decoder(16#49#)) OR
 					(reg_q880 AND symb_decoder(16#42#)) OR
 					(reg_q880 AND symb_decoder(16#53#)) OR
 					(reg_q880 AND symb_decoder(16#79#)) OR
 					(reg_q880 AND symb_decoder(16#6e#)) OR
 					(reg_q880 AND symb_decoder(16#4c#)) OR
 					(reg_q880 AND symb_decoder(16#74#)) OR
 					(reg_q880 AND symb_decoder(16#4a#)) OR
 					(reg_q880 AND symb_decoder(16#4b#)) OR
 					(reg_q880 AND symb_decoder(16#43#)) OR
 					(reg_q880 AND symb_decoder(16#52#)) OR
 					(reg_q880 AND symb_decoder(16#61#)) OR
 					(reg_q880 AND symb_decoder(16#57#)) OR
 					(reg_q880 AND symb_decoder(16#65#)) OR
 					(reg_q880 AND symb_decoder(16#75#)) OR
 					(reg_q880 AND symb_decoder(16#44#)) OR
 					(reg_q880 AND symb_decoder(16#47#)) OR
 					(reg_q880 AND symb_decoder(16#78#)) OR
 					(reg_q880 AND symb_decoder(16#64#)) OR
 					(reg_q880 AND symb_decoder(16#66#)) OR
 					(reg_q880 AND symb_decoder(16#63#)) OR
 					(reg_q880 AND symb_decoder(16#72#)) OR
 					(reg_q880 AND symb_decoder(16#48#));
reg_q2429_in <= (reg_q2427 AND symb_decoder(16#63#)) OR
 					(reg_q2427 AND symb_decoder(16#43#));
reg_q2526_in <= (reg_q2526 AND symb_decoder(16#35#)) OR
 					(reg_q2526 AND symb_decoder(16#32#)) OR
 					(reg_q2526 AND symb_decoder(16#39#)) OR
 					(reg_q2526 AND symb_decoder(16#36#)) OR
 					(reg_q2526 AND symb_decoder(16#38#)) OR
 					(reg_q2526 AND symb_decoder(16#33#)) OR
 					(reg_q2526 AND symb_decoder(16#37#)) OR
 					(reg_q2526 AND symb_decoder(16#34#)) OR
 					(reg_q2526 AND symb_decoder(16#31#)) OR
 					(reg_q2526 AND symb_decoder(16#30#)) OR
 					(reg_q2524 AND symb_decoder(16#37#)) OR
 					(reg_q2524 AND symb_decoder(16#35#)) OR
 					(reg_q2524 AND symb_decoder(16#30#)) OR
 					(reg_q2524 AND symb_decoder(16#36#)) OR
 					(reg_q2524 AND symb_decoder(16#31#)) OR
 					(reg_q2524 AND symb_decoder(16#39#)) OR
 					(reg_q2524 AND symb_decoder(16#38#)) OR
 					(reg_q2524 AND symb_decoder(16#33#)) OR
 					(reg_q2524 AND symb_decoder(16#32#)) OR
 					(reg_q2524 AND symb_decoder(16#34#));
reg_q2423_in <= (reg_q2421 AND symb_decoder(16#74#)) OR
 					(reg_q2421 AND symb_decoder(16#54#));
reg_q2425_in <= (reg_q2423 AND symb_decoder(16#61#)) OR
 					(reg_q2423 AND symb_decoder(16#41#));
reg_q2196_in <= (reg_q2194 AND symb_decoder(16#44#)) OR
 					(reg_q2194 AND symb_decoder(16#64#));
reg_q2198_in <= (reg_q2196 AND symb_decoder(16#41#)) OR
 					(reg_q2196 AND symb_decoder(16#61#));
reg_q854_in <= (reg_q852 AND symb_decoder(16#44#)) OR
 					(reg_q852 AND symb_decoder(16#64#));
reg_q612_in <= (reg_q610 AND symb_decoder(16#32#));
reg_q614_in <= (reg_q612 AND symb_decoder(16#65#)) OR
 					(reg_q612 AND symb_decoder(16#45#));
reg_q34_in <= (reg_q32 AND symb_decoder(16#54#)) OR
 					(reg_q32 AND symb_decoder(16#74#));
reg_q36_in <= (reg_q34 AND symb_decoder(16#45#)) OR
 					(reg_q34 AND symb_decoder(16#65#));
reg_q2072_in <= (reg_q2070 AND symb_decoder(16#50#));
reg_q884_in <= (reg_q882 AND symb_decoder(16#3a#));
reg_q1207_in <= (reg_q1207 AND symb_decoder(16#38#)) OR
 					(reg_q1207 AND symb_decoder(16#32#)) OR
 					(reg_q1207 AND symb_decoder(16#34#)) OR
 					(reg_q1207 AND symb_decoder(16#30#)) OR
 					(reg_q1207 AND symb_decoder(16#33#)) OR
 					(reg_q1207 AND symb_decoder(16#35#)) OR
 					(reg_q1207 AND symb_decoder(16#36#)) OR
 					(reg_q1207 AND symb_decoder(16#39#)) OR
 					(reg_q1207 AND symb_decoder(16#37#)) OR
 					(reg_q1207 AND symb_decoder(16#31#)) OR
 					(reg_q1205 AND symb_decoder(16#38#)) OR
 					(reg_q1205 AND symb_decoder(16#35#)) OR
 					(reg_q1205 AND symb_decoder(16#39#)) OR
 					(reg_q1205 AND symb_decoder(16#37#)) OR
 					(reg_q1205 AND symb_decoder(16#31#)) OR
 					(reg_q1205 AND symb_decoder(16#36#)) OR
 					(reg_q1205 AND symb_decoder(16#34#)) OR
 					(reg_q1205 AND symb_decoder(16#30#)) OR
 					(reg_q1205 AND symb_decoder(16#32#)) OR
 					(reg_q1205 AND symb_decoder(16#33#));
reg_q1985_in <= (reg_q1985 AND symb_decoder(16#30#)) OR
 					(reg_q1985 AND symb_decoder(16#35#)) OR
 					(reg_q1985 AND symb_decoder(16#31#)) OR
 					(reg_q1985 AND symb_decoder(16#36#)) OR
 					(reg_q1985 AND symb_decoder(16#34#)) OR
 					(reg_q1985 AND symb_decoder(16#39#)) OR
 					(reg_q1985 AND symb_decoder(16#32#)) OR
 					(reg_q1985 AND symb_decoder(16#33#)) OR
 					(reg_q1985 AND symb_decoder(16#37#)) OR
 					(reg_q1985 AND symb_decoder(16#38#)) OR
 					(reg_q1983 AND symb_decoder(16#33#)) OR
 					(reg_q1983 AND symb_decoder(16#31#)) OR
 					(reg_q1983 AND symb_decoder(16#34#)) OR
 					(reg_q1983 AND symb_decoder(16#30#)) OR
 					(reg_q1983 AND symb_decoder(16#32#)) OR
 					(reg_q1983 AND symb_decoder(16#39#)) OR
 					(reg_q1983 AND symb_decoder(16#36#)) OR
 					(reg_q1983 AND symb_decoder(16#37#)) OR
 					(reg_q1983 AND symb_decoder(16#38#)) OR
 					(reg_q1983 AND symb_decoder(16#35#));
reg_q1401_in <= (reg_q1399 AND symb_decoder(16#42#)) OR
 					(reg_q1399 AND symb_decoder(16#62#));
reg_q1403_in <= (reg_q1401 AND symb_decoder(16#45#)) OR
 					(reg_q1401 AND symb_decoder(16#65#));
reg_q38_in <= (reg_q36 AND symb_decoder(16#44#)) OR
 					(reg_q36 AND symb_decoder(16#64#));
reg_q1916_in <= (reg_q1914 AND symb_decoder(16#65#)) OR
 					(reg_q1914 AND symb_decoder(16#45#));
reg_q1800_in <= (reg_q1798 AND symb_decoder(16#53#)) OR
 					(reg_q1798 AND symb_decoder(16#73#));
reg_q1226_in <= (reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1225 AND symb_decoder(16#47#)) OR
 					(reg_q1225 AND symb_decoder(16#67#));
reg_q2093_in <= (reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2092 AND symb_decoder(16#75#)) OR
 					(reg_q2092 AND symb_decoder(16#55#));
reg_q758_in <= (reg_q756 AND symb_decoder(16#44#)) OR
 					(reg_q756 AND symb_decoder(16#64#));
reg_q2182_in <= (reg_q2180 AND symb_decoder(16#54#)) OR
 					(reg_q2180 AND symb_decoder(16#74#));
reg_q2184_in <= (reg_q2182 AND symb_decoder(16#69#)) OR
 					(reg_q2182 AND symb_decoder(16#49#));
reg_q598_in <= (reg_q596 AND symb_decoder(16#50#)) OR
 					(reg_q596 AND symb_decoder(16#70#));
reg_q600_in <= (reg_q598 AND symb_decoder(16#52#)) OR
 					(reg_q598 AND symb_decoder(16#72#));
reg_q1981_in <= (reg_q1981 AND symb_decoder(16#37#)) OR
 					(reg_q1981 AND symb_decoder(16#32#)) OR
 					(reg_q1981 AND symb_decoder(16#34#)) OR
 					(reg_q1981 AND symb_decoder(16#33#)) OR
 					(reg_q1981 AND symb_decoder(16#38#)) OR
 					(reg_q1981 AND symb_decoder(16#31#)) OR
 					(reg_q1981 AND symb_decoder(16#36#)) OR
 					(reg_q1981 AND symb_decoder(16#30#)) OR
 					(reg_q1981 AND symb_decoder(16#35#)) OR
 					(reg_q1981 AND symb_decoder(16#39#)) OR
 					(reg_q1979 AND symb_decoder(16#31#)) OR
 					(reg_q1979 AND symb_decoder(16#36#)) OR
 					(reg_q1979 AND symb_decoder(16#34#)) OR
 					(reg_q1979 AND symb_decoder(16#39#)) OR
 					(reg_q1979 AND symb_decoder(16#38#)) OR
 					(reg_q1979 AND symb_decoder(16#37#)) OR
 					(reg_q1979 AND symb_decoder(16#30#)) OR
 					(reg_q1979 AND symb_decoder(16#32#)) OR
 					(reg_q1979 AND symb_decoder(16#35#)) OR
 					(reg_q1979 AND symb_decoder(16#33#));
reg_q2062_in <= (reg_q2060 AND symb_decoder(16#66#));
reg_q1393_in <= (reg_q1391 AND symb_decoder(16#3a#));
reg_q474_in <= (reg_q472 AND symb_decoder(16#32#));
reg_q476_in <= (reg_q474 AND symb_decoder(16#30#));
reg_q2395_in <= (reg_q2393 AND symb_decoder(16#4f#)) OR
 					(reg_q2393 AND symb_decoder(16#6f#));
reg_q2397_in <= (reg_q2395 AND symb_decoder(16#6d#)) OR
 					(reg_q2395 AND symb_decoder(16#4d#));
reg_q1205_in <= (reg_q1203 AND symb_decoder(16#4e#)) OR
 					(reg_q1203 AND symb_decoder(16#6e#));
reg_q1924_in <= (reg_q1922 AND symb_decoder(16#42#)) OR
 					(reg_q1922 AND symb_decoder(16#62#));
reg_q2439_in <= (reg_q2437 AND symb_decoder(16#54#)) OR
 					(reg_q2437 AND symb_decoder(16#74#));
reg_q2441_in <= (reg_q2439 AND symb_decoder(16#61#)) OR
 					(reg_q2439 AND symb_decoder(16#41#));
reg_q630_in <= (reg_q628 AND symb_decoder(16#52#)) OR
 					(reg_q628 AND symb_decoder(16#72#));
reg_q1850_in <= (reg_q1848 AND symb_decoder(16#53#)) OR
 					(reg_q1848 AND symb_decoder(16#73#));
reg_q1888_in <= (reg_q1886 AND symb_decoder(16#48#)) OR
 					(reg_q1886 AND symb_decoder(16#68#));
reg_q1890_in <= (reg_q1888 AND symb_decoder(16#61#)) OR
 					(reg_q1888 AND symb_decoder(16#41#));
reg_q528_in <= (reg_q526 AND symb_decoder(16#2e#));
reg_q530_in <= (reg_q528 AND symb_decoder(16#35#)) OR
 					(reg_q528 AND symb_decoder(16#39#)) OR
 					(reg_q528 AND symb_decoder(16#31#)) OR
 					(reg_q528 AND symb_decoder(16#38#)) OR
 					(reg_q528 AND symb_decoder(16#34#)) OR
 					(reg_q528 AND symb_decoder(16#32#)) OR
 					(reg_q528 AND symb_decoder(16#33#)) OR
 					(reg_q528 AND symb_decoder(16#36#)) OR
 					(reg_q528 AND symb_decoder(16#37#)) OR
 					(reg_q528 AND symb_decoder(16#30#)) OR
 					(reg_q530 AND symb_decoder(16#31#)) OR
 					(reg_q530 AND symb_decoder(16#35#)) OR
 					(reg_q530 AND symb_decoder(16#36#)) OR
 					(reg_q530 AND symb_decoder(16#39#)) OR
 					(reg_q530 AND symb_decoder(16#30#)) OR
 					(reg_q530 AND symb_decoder(16#34#)) OR
 					(reg_q530 AND symb_decoder(16#37#)) OR
 					(reg_q530 AND symb_decoder(16#32#)) OR
 					(reg_q530 AND symb_decoder(16#38#)) OR
 					(reg_q530 AND symb_decoder(16#33#));
reg_q606_in <= (reg_q604 AND symb_decoder(16#56#)) OR
 					(reg_q604 AND symb_decoder(16#76#));
reg_q608_in <= (reg_q606 AND symb_decoder(16#30#)) OR
 					(reg_q606 AND symb_decoder(16#32#)) OR
 					(reg_q606 AND symb_decoder(16#31#)) OR
 					(reg_q606 AND symb_decoder(16#37#)) OR
 					(reg_q606 AND symb_decoder(16#39#)) OR
 					(reg_q606 AND symb_decoder(16#35#)) OR
 					(reg_q606 AND symb_decoder(16#34#)) OR
 					(reg_q606 AND symb_decoder(16#36#)) OR
 					(reg_q606 AND symb_decoder(16#33#)) OR
 					(reg_q606 AND symb_decoder(16#38#)) OR
 					(reg_q608 AND symb_decoder(16#39#)) OR
 					(reg_q608 AND symb_decoder(16#33#)) OR
 					(reg_q608 AND symb_decoder(16#37#)) OR
 					(reg_q608 AND symb_decoder(16#38#)) OR
 					(reg_q608 AND symb_decoder(16#31#)) OR
 					(reg_q608 AND symb_decoder(16#34#)) OR
 					(reg_q608 AND symb_decoder(16#32#)) OR
 					(reg_q608 AND symb_decoder(16#35#)) OR
 					(reg_q608 AND symb_decoder(16#30#)) OR
 					(reg_q608 AND symb_decoder(16#36#));
reg_q2431_in <= (reg_q2429 AND symb_decoder(16#4f#)) OR
 					(reg_q2429 AND symb_decoder(16#6f#));
reg_q2433_in <= (reg_q2431 AND symb_decoder(16#4e#)) OR
 					(reg_q2431 AND symb_decoder(16#6e#));
reg_q1987_in <= (reg_q1985 AND symb_decoder(16#2e#));
reg_q1989_in <= (reg_q1987 AND symb_decoder(16#30#)) OR
 					(reg_q1987 AND symb_decoder(16#34#)) OR
 					(reg_q1987 AND symb_decoder(16#32#)) OR
 					(reg_q1987 AND symb_decoder(16#39#)) OR
 					(reg_q1987 AND symb_decoder(16#38#)) OR
 					(reg_q1987 AND symb_decoder(16#33#)) OR
 					(reg_q1987 AND symb_decoder(16#37#)) OR
 					(reg_q1987 AND symb_decoder(16#31#)) OR
 					(reg_q1987 AND symb_decoder(16#35#)) OR
 					(reg_q1987 AND symb_decoder(16#36#)) OR
 					(reg_q1989 AND symb_decoder(16#33#)) OR
 					(reg_q1989 AND symb_decoder(16#39#)) OR
 					(reg_q1989 AND symb_decoder(16#35#)) OR
 					(reg_q1989 AND symb_decoder(16#32#)) OR
 					(reg_q1989 AND symb_decoder(16#36#)) OR
 					(reg_q1989 AND symb_decoder(16#34#)) OR
 					(reg_q1989 AND symb_decoder(16#38#)) OR
 					(reg_q1989 AND symb_decoder(16#30#)) OR
 					(reg_q1989 AND symb_decoder(16#31#)) OR
 					(reg_q1989 AND symb_decoder(16#37#));
reg_q1832_in <= (reg_q1830 AND symb_decoder(16#68#)) OR
 					(reg_q1830 AND symb_decoder(16#48#));
reg_q1834_in <= (reg_q1832 AND symb_decoder(16#77#)) OR
 					(reg_q1832 AND symb_decoder(16#57#));
reg_q799_in <= (reg_q797 AND symb_decoder(16#2e#));
reg_q801_in <= (reg_q799 AND symb_decoder(16#33#)) OR
 					(reg_q799 AND symb_decoder(16#30#)) OR
 					(reg_q799 AND symb_decoder(16#34#)) OR
 					(reg_q799 AND symb_decoder(16#39#)) OR
 					(reg_q799 AND symb_decoder(16#38#)) OR
 					(reg_q799 AND symb_decoder(16#37#)) OR
 					(reg_q799 AND symb_decoder(16#36#)) OR
 					(reg_q799 AND symb_decoder(16#35#)) OR
 					(reg_q799 AND symb_decoder(16#31#)) OR
 					(reg_q799 AND symb_decoder(16#32#)) OR
 					(reg_q801 AND symb_decoder(16#37#)) OR
 					(reg_q801 AND symb_decoder(16#35#)) OR
 					(reg_q801 AND symb_decoder(16#30#)) OR
 					(reg_q801 AND symb_decoder(16#32#)) OR
 					(reg_q801 AND symb_decoder(16#38#)) OR
 					(reg_q801 AND symb_decoder(16#39#)) OR
 					(reg_q801 AND symb_decoder(16#31#)) OR
 					(reg_q801 AND symb_decoder(16#36#)) OR
 					(reg_q801 AND symb_decoder(16#34#)) OR
 					(reg_q801 AND symb_decoder(16#33#));
reg_q2415_in <= (reg_q2413 AND symb_decoder(16#49#)) OR
 					(reg_q2413 AND symb_decoder(16#69#));
reg_q1910_in <= (reg_q1908 AND symb_decoder(16#4d#)) OR
 					(reg_q1908 AND symb_decoder(16#6d#));
reg_q1912_in <= (reg_q1910 AND symb_decoder(16#4f#)) OR
 					(reg_q1910 AND symb_decoder(16#6f#));
reg_q578_in <= (reg_q576 AND symb_decoder(16#31#));
reg_q580_in <= (reg_q578 AND symb_decoder(16#25#));
reg_q1818_in <= (reg_q1816 AND symb_decoder(16#76#)) OR
 					(reg_q1816 AND symb_decoder(16#56#));
reg_q1820_in <= (reg_q1818 AND symb_decoder(16#37#)) OR
 					(reg_q1818 AND symb_decoder(16#36#)) OR
 					(reg_q1818 AND symb_decoder(16#30#)) OR
 					(reg_q1818 AND symb_decoder(16#38#)) OR
 					(reg_q1818 AND symb_decoder(16#39#)) OR
 					(reg_q1818 AND symb_decoder(16#32#)) OR
 					(reg_q1818 AND symb_decoder(16#31#)) OR
 					(reg_q1818 AND symb_decoder(16#33#)) OR
 					(reg_q1818 AND symb_decoder(16#34#)) OR
 					(reg_q1818 AND symb_decoder(16#35#)) OR
 					(reg_q1820 AND symb_decoder(16#30#)) OR
 					(reg_q1820 AND symb_decoder(16#33#)) OR
 					(reg_q1820 AND symb_decoder(16#36#)) OR
 					(reg_q1820 AND symb_decoder(16#39#)) OR
 					(reg_q1820 AND symb_decoder(16#37#)) OR
 					(reg_q1820 AND symb_decoder(16#35#)) OR
 					(reg_q1820 AND symb_decoder(16#32#)) OR
 					(reg_q1820 AND symb_decoder(16#31#)) OR
 					(reg_q1820 AND symb_decoder(16#34#)) OR
 					(reg_q1820 AND symb_decoder(16#38#));
reg_q1842_in <= (reg_q1840 AND symb_decoder(16#4c#)) OR
 					(reg_q1840 AND symb_decoder(16#6c#));
reg_q1844_in <= (reg_q1842 AND symb_decoder(16#45#)) OR
 					(reg_q1842 AND symb_decoder(16#65#));
reg_q18_in <= (reg_q16 AND symb_decoder(16#69#)) OR
 					(reg_q16 AND symb_decoder(16#49#));
reg_q1646_in <= (reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q1645 AND symb_decoder(16#72#)) OR
 					(reg_q1645 AND symb_decoder(16#52#));
reg_q506_in <= (reg_q504 AND symb_decoder(16#3a#));
reg_q508_in <= (reg_q506 AND symb_decoder(16#25#));
reg_q628_in <= (reg_q626 AND symb_decoder(16#45#)) OR
 					(reg_q626 AND symb_decoder(16#65#));
reg_q131_in <= (reg_q129 AND symb_decoder(16#63#)) OR
 					(reg_q129 AND symb_decoder(16#43#));
reg_q1381_in <= (reg_q1379 AND symb_decoder(16#45#)) OR
 					(reg_q1379 AND symb_decoder(16#65#));
reg_q1948_in <= (reg_q1946 AND symb_decoder(16#41#)) OR
 					(reg_q1946 AND symb_decoder(16#61#));
reg_q1950_in <= (reg_q1948 AND symb_decoder(16#72#)) OR
 					(reg_q1948 AND symb_decoder(16#52#));
reg_q1605_in <= (reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q1604 AND symb_decoder(16#6e#)) OR
 					(reg_q1604 AND symb_decoder(16#4e#));
reg_q14_in <= (reg_q12 AND symb_decoder(16#45#)) OR
 					(reg_q12 AND symb_decoder(16#65#));
reg_q1979_in <= (reg_q1997 AND symb_decoder(16#23#)) OR
 					(reg_q1975 AND symb_decoder(16#23#));
reg_q795_in <= (reg_q813 AND symb_decoder(16#5e#)) OR
 					(reg_q791 AND symb_decoder(16#5e#));
reg_q797_in <= (reg_q795 AND symb_decoder(16#33#)) OR
 					(reg_q795 AND symb_decoder(16#30#)) OR
 					(reg_q795 AND symb_decoder(16#34#)) OR
 					(reg_q795 AND symb_decoder(16#36#)) OR
 					(reg_q795 AND symb_decoder(16#38#)) OR
 					(reg_q795 AND symb_decoder(16#35#)) OR
 					(reg_q795 AND symb_decoder(16#39#)) OR
 					(reg_q795 AND symb_decoder(16#37#)) OR
 					(reg_q795 AND symb_decoder(16#32#)) OR
 					(reg_q795 AND symb_decoder(16#31#)) OR
 					(reg_q797 AND symb_decoder(16#33#)) OR
 					(reg_q797 AND symb_decoder(16#37#)) OR
 					(reg_q797 AND symb_decoder(16#31#)) OR
 					(reg_q797 AND symb_decoder(16#32#)) OR
 					(reg_q797 AND symb_decoder(16#34#)) OR
 					(reg_q797 AND symb_decoder(16#36#)) OR
 					(reg_q797 AND symb_decoder(16#35#)) OR
 					(reg_q797 AND symb_decoder(16#38#)) OR
 					(reg_q797 AND symb_decoder(16#39#)) OR
 					(reg_q797 AND symb_decoder(16#30#));
reg_q510_in <= (reg_q508 AND symb_decoder(16#32#));
reg_q1814_in <= (reg_q1812 AND symb_decoder(16#52#)) OR
 					(reg_q1812 AND symb_decoder(16#72#));
reg_q562_in <= (reg_q560 AND symb_decoder(16#64#)) OR
 					(reg_q560 AND symb_decoder(16#44#));
reg_q564_in <= (reg_q562 AND symb_decoder(16#59#)) OR
 					(reg_q562 AND symb_decoder(16#79#));
reg_q943_in <= (reg_q943 AND symb_decoder(16#36#)) OR
 					(reg_q943 AND symb_decoder(16#37#)) OR
 					(reg_q943 AND symb_decoder(16#34#)) OR
 					(reg_q943 AND symb_decoder(16#32#)) OR
 					(reg_q943 AND symb_decoder(16#31#)) OR
 					(reg_q943 AND symb_decoder(16#38#)) OR
 					(reg_q943 AND symb_decoder(16#35#)) OR
 					(reg_q943 AND symb_decoder(16#30#)) OR
 					(reg_q943 AND symb_decoder(16#33#)) OR
 					(reg_q943 AND symb_decoder(16#39#)) OR
 					(reg_q941 AND symb_decoder(16#38#)) OR
 					(reg_q941 AND symb_decoder(16#30#)) OR
 					(reg_q941 AND symb_decoder(16#37#)) OR
 					(reg_q941 AND symb_decoder(16#34#)) OR
 					(reg_q941 AND symb_decoder(16#39#)) OR
 					(reg_q941 AND symb_decoder(16#32#)) OR
 					(reg_q941 AND symb_decoder(16#36#)) OR
 					(reg_q941 AND symb_decoder(16#31#)) OR
 					(reg_q941 AND symb_decoder(16#35#)) OR
 					(reg_q941 AND symb_decoder(16#33#));
reg_q1942_in <= (reg_q1940 AND symb_decoder(16#50#)) OR
 					(reg_q1940 AND symb_decoder(16#70#));
reg_q1944_in <= (reg_q1942 AND symb_decoder(16#59#)) OR
 					(reg_q1942 AND symb_decoder(16#79#));
reg_q634_in <= (reg_q632 AND symb_decoder(16#6f#)) OR
 					(reg_q632 AND symb_decoder(16#4f#));
reg_q1213_in <= (reg_q1211 AND symb_decoder(16#49#)) OR
 					(reg_q1211 AND symb_decoder(16#69#));
reg_q1858_in <= (reg_q1856 AND symb_decoder(16#49#)) OR
 					(reg_q1856 AND symb_decoder(16#69#));
reg_q1860_in <= (reg_q1858 AND symb_decoder(16#64#)) OR
 					(reg_q1858 AND symb_decoder(16#44#));
reg_q1836_in <= (reg_q1834 AND symb_decoder(16#49#)) OR
 					(reg_q1834 AND symb_decoder(16#69#));
reg_q1525_in <= (reg_q1523 AND symb_decoder(16#45#)) OR
 					(reg_q1523 AND symb_decoder(16#65#));
reg_q878_in <= (reg_q876 AND symb_decoder(16#37#)) OR
 					(reg_q876 AND symb_decoder(16#33#)) OR
 					(reg_q876 AND symb_decoder(16#32#)) OR
 					(reg_q876 AND symb_decoder(16#36#)) OR
 					(reg_q876 AND symb_decoder(16#34#)) OR
 					(reg_q876 AND symb_decoder(16#30#)) OR
 					(reg_q876 AND symb_decoder(16#31#)) OR
 					(reg_q876 AND symb_decoder(16#35#)) OR
 					(reg_q876 AND symb_decoder(16#39#)) OR
 					(reg_q876 AND symb_decoder(16#38#));
reg_q1464_in <= (reg_q1462 AND symb_decoder(16#41#)) OR
 					(reg_q1462 AND symb_decoder(16#61#));
reg_q787_in <= (reg_q785 AND symb_decoder(16#4e#)) OR
 					(reg_q785 AND symb_decoder(16#6e#));
reg_q1862_in <= (reg_q1860 AND symb_decoder(16#6f#)) OR
 					(reg_q1860 AND symb_decoder(16#4f#));
reg_q1922_in <= (reg_q1920 AND symb_decoder(16#45#)) OR
 					(reg_q1920 AND symb_decoder(16#65#));
reg_q1550_in <= (reg_q1548 AND symb_decoder(16#74#)) OR
 					(reg_q1548 AND symb_decoder(16#54#));
reg_q1870_in <= (reg_q1868 AND symb_decoder(16#50#)) OR
 					(reg_q1868 AND symb_decoder(16#70#));
reg_q1991_in <= (reg_q1989 AND symb_decoder(16#2e#));
reg_q1993_in <= (reg_q1991 AND symb_decoder(16#39#)) OR
 					(reg_q1991 AND symb_decoder(16#34#)) OR
 					(reg_q1991 AND symb_decoder(16#37#)) OR
 					(reg_q1991 AND symb_decoder(16#31#)) OR
 					(reg_q1991 AND symb_decoder(16#38#)) OR
 					(reg_q1991 AND symb_decoder(16#35#)) OR
 					(reg_q1991 AND symb_decoder(16#30#)) OR
 					(reg_q1991 AND symb_decoder(16#32#)) OR
 					(reg_q1991 AND symb_decoder(16#33#)) OR
 					(reg_q1991 AND symb_decoder(16#36#)) OR
 					(reg_q1993 AND symb_decoder(16#34#)) OR
 					(reg_q1993 AND symb_decoder(16#39#)) OR
 					(reg_q1993 AND symb_decoder(16#33#)) OR
 					(reg_q1993 AND symb_decoder(16#38#)) OR
 					(reg_q1993 AND symb_decoder(16#36#)) OR
 					(reg_q1993 AND symb_decoder(16#32#)) OR
 					(reg_q1993 AND symb_decoder(16#30#)) OR
 					(reg_q1993 AND symb_decoder(16#37#)) OR
 					(reg_q1993 AND symb_decoder(16#31#)) OR
 					(reg_q1993 AND symb_decoder(16#35#));
reg_q803_in <= (reg_q801 AND symb_decoder(16#2e#));
reg_q807_in <= (reg_q805 AND symb_decoder(16#2e#));
reg_q809_in <= (reg_q807 AND symb_decoder(16#34#)) OR
 					(reg_q807 AND symb_decoder(16#38#)) OR
 					(reg_q807 AND symb_decoder(16#35#)) OR
 					(reg_q807 AND symb_decoder(16#31#)) OR
 					(reg_q807 AND symb_decoder(16#39#)) OR
 					(reg_q807 AND symb_decoder(16#37#)) OR
 					(reg_q807 AND symb_decoder(16#32#)) OR
 					(reg_q807 AND symb_decoder(16#36#)) OR
 					(reg_q807 AND symb_decoder(16#33#)) OR
 					(reg_q807 AND symb_decoder(16#30#)) OR
 					(reg_q809 AND symb_decoder(16#32#)) OR
 					(reg_q809 AND symb_decoder(16#35#)) OR
 					(reg_q809 AND symb_decoder(16#39#)) OR
 					(reg_q809 AND symb_decoder(16#38#)) OR
 					(reg_q809 AND symb_decoder(16#33#)) OR
 					(reg_q809 AND symb_decoder(16#31#)) OR
 					(reg_q809 AND symb_decoder(16#30#)) OR
 					(reg_q809 AND symb_decoder(16#37#)) OR
 					(reg_q809 AND symb_decoder(16#36#)) OR
 					(reg_q809 AND symb_decoder(16#34#));
reg_q478_in <= (reg_q476 AND symb_decoder(16#30#));
reg_q524_in <= (reg_q522 AND symb_decoder(16#2e#));
reg_q805_in <= (reg_q803 AND symb_decoder(16#37#)) OR
 					(reg_q803 AND symb_decoder(16#30#)) OR
 					(reg_q803 AND symb_decoder(16#38#)) OR
 					(reg_q803 AND symb_decoder(16#33#)) OR
 					(reg_q803 AND symb_decoder(16#39#)) OR
 					(reg_q803 AND symb_decoder(16#35#)) OR
 					(reg_q803 AND symb_decoder(16#36#)) OR
 					(reg_q803 AND symb_decoder(16#34#)) OR
 					(reg_q803 AND symb_decoder(16#32#)) OR
 					(reg_q803 AND symb_decoder(16#31#)) OR
 					(reg_q805 AND symb_decoder(16#36#)) OR
 					(reg_q805 AND symb_decoder(16#30#)) OR
 					(reg_q805 AND symb_decoder(16#33#)) OR
 					(reg_q805 AND symb_decoder(16#39#)) OR
 					(reg_q805 AND symb_decoder(16#38#)) OR
 					(reg_q805 AND symb_decoder(16#34#)) OR
 					(reg_q805 AND symb_decoder(16#32#)) OR
 					(reg_q805 AND symb_decoder(16#37#)) OR
 					(reg_q805 AND symb_decoder(16#31#)) OR
 					(reg_q805 AND symb_decoder(16#35#));
reg_q1219_in <= (reg_q1217 AND symb_decoder(16#38#)) OR
 					(reg_q1217 AND symb_decoder(16#30#)) OR
 					(reg_q1217 AND symb_decoder(16#35#)) OR
 					(reg_q1217 AND symb_decoder(16#33#)) OR
 					(reg_q1217 AND symb_decoder(16#31#)) OR
 					(reg_q1217 AND symb_decoder(16#37#)) OR
 					(reg_q1217 AND symb_decoder(16#32#)) OR
 					(reg_q1217 AND symb_decoder(16#34#)) OR
 					(reg_q1217 AND symb_decoder(16#36#)) OR
 					(reg_q1217 AND symb_decoder(16#39#)) OR
 					(reg_q1219 AND symb_decoder(16#37#)) OR
 					(reg_q1219 AND symb_decoder(16#31#)) OR
 					(reg_q1219 AND symb_decoder(16#35#)) OR
 					(reg_q1219 AND symb_decoder(16#34#)) OR
 					(reg_q1219 AND symb_decoder(16#39#)) OR
 					(reg_q1219 AND symb_decoder(16#32#)) OR
 					(reg_q1219 AND symb_decoder(16#38#)) OR
 					(reg_q1219 AND symb_decoder(16#36#)) OR
 					(reg_q1219 AND symb_decoder(16#33#)) OR
 					(reg_q1219 AND symb_decoder(16#30#));
reg_q1796_in <= (reg_q1794 AND symb_decoder(16#42#)) OR
 					(reg_q1794 AND symb_decoder(16#62#));
reg_q648_in <= (reg_q646 AND symb_decoder(16#32#));
reg_q650_in <= (reg_q648 AND symb_decoder(16#31#));
reg_q1822_in <= (reg_q1820 AND symb_decoder(16#2e#));
reg_q1824_in <= (reg_q1822 AND symb_decoder(16#39#)) OR
 					(reg_q1822 AND symb_decoder(16#33#)) OR
 					(reg_q1822 AND symb_decoder(16#36#)) OR
 					(reg_q1822 AND symb_decoder(16#35#)) OR
 					(reg_q1822 AND symb_decoder(16#30#)) OR
 					(reg_q1822 AND symb_decoder(16#34#)) OR
 					(reg_q1822 AND symb_decoder(16#38#)) OR
 					(reg_q1822 AND symb_decoder(16#37#)) OR
 					(reg_q1822 AND symb_decoder(16#31#)) OR
 					(reg_q1822 AND symb_decoder(16#32#)) OR
 					(reg_q1824 AND symb_decoder(16#37#)) OR
 					(reg_q1824 AND symb_decoder(16#34#)) OR
 					(reg_q1824 AND symb_decoder(16#38#)) OR
 					(reg_q1824 AND symb_decoder(16#30#)) OR
 					(reg_q1824 AND symb_decoder(16#35#)) OR
 					(reg_q1824 AND symb_decoder(16#39#)) OR
 					(reg_q1824 AND symb_decoder(16#36#)) OR
 					(reg_q1824 AND symb_decoder(16#31#)) OR
 					(reg_q1824 AND symb_decoder(16#33#)) OR
 					(reg_q1824 AND symb_decoder(16#32#));
reg_q2192_in <= (reg_q2190 AND symb_decoder(16#6c#)) OR
 					(reg_q2190 AND symb_decoder(16#4c#));
reg_q1397_in <= (reg_q1395 AND symb_decoder(16#43#)) OR
 					(reg_q1395 AND symb_decoder(16#63#));
reg_q789_in <= (reg_q787 AND symb_decoder(16#46#)) OR
 					(reg_q787 AND symb_decoder(16#66#));
reg_q1830_in <= (reg_q1828 AND symb_decoder(16#63#)) OR
 					(reg_q1828 AND symb_decoder(16#43#));
reg_q1113_in <= (reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q1112 AND symb_decoder(16#66#)) OR
 					(reg_q1112 AND symb_decoder(16#46#));
reg_q1983_in <= (reg_q1981 AND symb_decoder(16#2e#));
reg_q1872_in <= (reg_q1870 AND symb_decoder(16#4f#)) OR
 					(reg_q1870 AND symb_decoder(16#6f#));
reg_q2186_in <= (reg_q2184 AND symb_decoder(16#6f#)) OR
 					(reg_q2184 AND symb_decoder(16#4f#));
reg_q2188_in <= (reg_q2186 AND symb_decoder(16#6e#)) OR
 					(reg_q2186 AND symb_decoder(16#4e#));
reg_q2162_in <= (reg_q2160 AND symb_decoder(16#64#)) OR
 					(reg_q2160 AND symb_decoder(16#44#));
reg_q1846_in <= (reg_q1844 AND symb_decoder(16#52#)) OR
 					(reg_q1844 AND symb_decoder(16#72#));
reg_q540_in <= (reg_q538 AND symb_decoder(16#32#));
reg_q542_in <= (reg_q540 AND symb_decoder(16#30#));
reg_q1798_in <= (reg_q1796 AND symb_decoder(16#75#)) OR
 					(reg_q1796 AND symb_decoder(16#55#));
reg_q1936_in <= (reg_q1934 AND symb_decoder(16#64#)) OR
 					(reg_q1934 AND symb_decoder(16#44#));
reg_q2200_in <= (reg_q2198 AND symb_decoder(16#65#)) OR
 					(reg_q2198 AND symb_decoder(16#45#));
reg_q941_in <= (reg_q939 AND symb_decoder(16#2e#));
reg_q572_in <= (reg_q570 AND symb_decoder(16#31#));
reg_q574_in <= (reg_q572 AND symb_decoder(16#25#));
reg_q862_in <= (reg_q860 AND symb_decoder(16#45#)) OR
 					(reg_q860 AND symb_decoder(16#65#));
reg_q1161_in <= (reg_q1159 AND symb_decoder(16#43#)) OR
 					(reg_q1159 AND symb_decoder(16#63#));
reg_q2524_in <= (reg_q2522 AND symb_decoder(16#72#)) OR
 					(reg_q2522 AND symb_decoder(16#52#));
reg_q638_in <= (reg_q636 AND symb_decoder(16#6c#)) OR
 					(reg_q636 AND symb_decoder(16#4c#));
reg_q640_in <= (reg_q638 AND symb_decoder(16#49#)) OR
 					(reg_q638 AND symb_decoder(16#69#));
reg_q594_in <= (reg_q592 AND symb_decoder(16#58#)) OR
 					(reg_q592 AND symb_decoder(16#78#));
reg_q32_in <= (reg_q30 AND symb_decoder(16#55#)) OR
 					(reg_q30 AND symb_decoder(16#75#));
reg_q872_in <= (reg_q870 AND symb_decoder(16#54#)) OR
 					(reg_q870 AND symb_decoder(16#74#));
reg_q2468_in <= (reg_q2695 AND symb_decoder(16#2a#));
reg_q866_in <= (reg_q864 AND symb_decoder(16#6c#)) OR
 					(reg_q864 AND symb_decoder(16#4c#));
reg_q868_in <= (reg_q866 AND symb_decoder(16#49#)) OR
 					(reg_q866 AND symb_decoder(16#69#));
reg_q870_in <= (reg_q868 AND symb_decoder(16#73#)) OR
 					(reg_q868 AND symb_decoder(16#53#));
reg_q1399_in <= (reg_q1397 AND symb_decoder(16#59#)) OR
 					(reg_q1397 AND symb_decoder(16#79#));
reg_q1928_in <= (reg_q1926 AND symb_decoder(16#42#)) OR
 					(reg_q1926 AND symb_decoder(16#62#));
reg_q642_in <= (reg_q640 AND symb_decoder(16#6e#)) OR
 					(reg_q640 AND symb_decoder(16#4e#));
reg_q644_in <= (reg_q642 AND symb_decoder(16#65#)) OR
 					(reg_q642 AND symb_decoder(16#45#));
reg_q2487_in <= (reg_q2485 AND symb_decoder(16#50#));
reg_q2489_in <= (reg_q2487 AND symb_decoder(16#4f#));
reg_q636_in <= (reg_q634 AND symb_decoder(16#6e#)) OR
 					(reg_q634 AND symb_decoder(16#4e#));
reg_q552_in <= (reg_q550 AND symb_decoder(16#54#)) OR
 					(reg_q550 AND symb_decoder(16#74#));
reg_q554_in <= (reg_q552 AND symb_decoder(16#5f#));
reg_q1365_in <= (reg_q1363 AND symb_decoder(16#32#));
reg_q1367_in <= (reg_q1365 AND symb_decoder(16#45#)) OR
 					(reg_q1365 AND symb_decoder(16#65#));
reg_q1812_in <= (reg_q1810 AND symb_decoder(16#45#)) OR
 					(reg_q1810 AND symb_decoder(16#65#));
reg_q1371_in <= (reg_q1369 AND symb_decoder(16#45#)) OR
 					(reg_q1369 AND symb_decoder(16#65#));
reg_q2399_in <= (reg_q2397 AND symb_decoder(16#50#)) OR
 					(reg_q2397 AND symb_decoder(16#70#));
reg_q2401_in <= (reg_q2399 AND symb_decoder(16#72#)) OR
 					(reg_q2399 AND symb_decoder(16#52#));
reg_q1908_in <= (reg_q1906 AND symb_decoder(16#65#)) OR
 					(reg_q1906 AND symb_decoder(16#45#));
reg_q584_in <= (reg_q582 AND symb_decoder(16#31#));
reg_q586_in <= (reg_q584 AND symb_decoder(16#6f#)) OR
 					(reg_q584 AND symb_decoder(16#4f#));
reg_q576_in <= (reg_q574 AND symb_decoder(16#32#));
reg_q20_in <= (reg_q18 AND symb_decoder(16#73#)) OR
 					(reg_q18 AND symb_decoder(16#53#));
reg_q2435_in <= (reg_q2433 AND symb_decoder(16#65#)) OR
 					(reg_q2433 AND symb_decoder(16#45#));
reg_q2437_in <= (reg_q2435 AND symb_decoder(16#63#)) OR
 					(reg_q2435 AND symb_decoder(16#43#));
reg_q2413_in <= (reg_q2411 AND symb_decoder(16#73#)) OR
 					(reg_q2411 AND symb_decoder(16#53#));
reg_q560_in <= (reg_q558 AND symb_decoder(16#4f#)) OR
 					(reg_q558 AND symb_decoder(16#6f#));
reg_q1804_in <= (reg_q1802 AND symb_decoder(16#53#)) OR
 					(reg_q1802 AND symb_decoder(16#73#));
reg_q1806_in <= (reg_q1804 AND symb_decoder(16#65#)) OR
 					(reg_q1804 AND symb_decoder(16#45#));
reg_q472_in <= (reg_q470 AND symb_decoder(16#25#));
reg_q546_in <= (reg_q544 AND symb_decoder(16#50#)) OR
 					(reg_q544 AND symb_decoder(16#70#));
reg_q548_in <= (reg_q546 AND symb_decoder(16#6f#)) OR
 					(reg_q546 AND symb_decoder(16#4f#));
reg_q2493_in <= (reg_q2491 AND symb_decoder(16#54#));
reg_q582_in <= (reg_q580 AND symb_decoder(16#32#));
reg_q492_in <= (reg_q490 AND symb_decoder(16#30#));
reg_q494_in <= (reg_q492 AND symb_decoder(16#6f#)) OR
 					(reg_q492 AND symb_decoder(16#4f#));
reg_q602_in <= (reg_q600 AND symb_decoder(16#6f#)) OR
 					(reg_q600 AND symb_decoder(16#4f#));
reg_q2082_in <= (reg_q2080 AND symb_decoder(16#76#));
reg_q2084_in <= (reg_q2082 AND symb_decoder(16#65#));
reg_q2190_in <= (reg_q2188 AND symb_decoder(16#41#)) OR
 					(reg_q2188 AND symb_decoder(16#61#));
reg_q1838_in <= (reg_q1836 AND symb_decoder(16#6e#)) OR
 					(reg_q1836 AND symb_decoder(16#4e#));
reg_q1898_in <= (reg_q1896 AND symb_decoder(16#6e#)) OR
 					(reg_q1896 AND symb_decoder(16#4e#));
reg_q1900_in <= (reg_q1898 AND symb_decoder(16#65#)) OR
 					(reg_q1898 AND symb_decoder(16#45#));
reg_q8_in <= (reg_q6 AND symb_decoder(16#66#)) OR
 					(reg_q6 AND symb_decoder(16#46#));
reg_q496_in <= (reg_q494 AND symb_decoder(16#6e#)) OR
 					(reg_q494 AND symb_decoder(16#4e#));
reg_q498_in <= (reg_q496 AND symb_decoder(16#6c#)) OR
 					(reg_q496 AND symb_decoder(16#4c#));
reg_q462_in <= (reg_q460 AND symb_decoder(16#3d#));
reg_q464_in <= (reg_q462 AND symb_decoder(16#46#)) OR
 					(reg_q462 AND symb_decoder(16#66#));
reg_q568_in <= (reg_q566 AND symb_decoder(16#25#));
reg_q1930_in <= (reg_q1928 AND symb_decoder(16#61#)) OR
 					(reg_q1928 AND symb_decoder(16#41#));
reg_q1932_in <= (reg_q1930 AND symb_decoder(16#73#)) OR
 					(reg_q1930 AND symb_decoder(16#53#));
reg_q512_in <= (reg_q510 AND symb_decoder(16#30#));
reg_q1914_in <= (reg_q1912 AND symb_decoder(16#54#)) OR
 					(reg_q1912 AND symb_decoder(16#74#));
reg_q1379_in <= (reg_q1377 AND symb_decoder(16#6c#)) OR
 					(reg_q1377 AND symb_decoder(16#4c#));
reg_q1199_in <= (reg_q1197 AND symb_decoder(16#74#)) OR
 					(reg_q1197 AND symb_decoder(16#54#));
reg_q544_in <= (reg_q542 AND symb_decoder(16#5b#));
reg_q470_in <= (reg_q468 AND symb_decoder(16#72#)) OR
 					(reg_q468 AND symb_decoder(16#52#));
reg_q2508_in <= (reg_q2506 AND symb_decoder(16#52#));
reg_q480_in <= (reg_q478 AND symb_decoder(16#2e#));
reg_q482_in <= (reg_q480 AND symb_decoder(16#32#));
reg_q500_in <= (reg_q498 AND symb_decoder(16#49#)) OR
 					(reg_q498 AND symb_decoder(16#69#));
reg_q1894_in <= (reg_q1892 AND symb_decoder(16#4f#)) OR
 					(reg_q1892 AND symb_decoder(16#6f#));
reg_q1896_in <= (reg_q1894 AND symb_decoder(16#77#)) OR
 					(reg_q1894 AND symb_decoder(16#57#));
reg_q820_in <= (reg_q818 AND symb_decoder(16#6d#)) OR
 					(reg_q818 AND symb_decoder(16#4d#));
reg_q905_in <= (reg_q903 AND symb_decoder(16#61#)) OR
 					(reg_q903 AND symb_decoder(16#41#));
reg_q24_in <= (reg_q22 AND symb_decoder(16#45#)) OR
 					(reg_q22 AND symb_decoder(16#65#));
reg_q1856_in <= (reg_q1854 AND symb_decoder(16#56#)) OR
 					(reg_q1854 AND symb_decoder(16#76#));
reg_q1203_in <= (reg_q1201 AND symb_decoder(16#4f#)) OR
 					(reg_q1201 AND symb_decoder(16#6f#));
reg_q1934_in <= (reg_q1932 AND symb_decoder(16#45#)) OR
 					(reg_q1932 AND symb_decoder(16#65#));
reg_q736_in <= (reg_q734 AND symb_decoder(16#63#)) OR
 					(reg_q734 AND symb_decoder(16#43#));
reg_q484_in <= (reg_q482 AND symb_decoder(16#2e#));
reg_q486_in <= (reg_q484 AND symb_decoder(16#30#));
reg_q550_in <= (reg_q548 AND symb_decoder(16#52#)) OR
 					(reg_q548 AND symb_decoder(16#72#));
reg_q2086_in <= (reg_q2084 AND symb_decoder(16#72#));
reg_q2088_in <= (reg_q2086 AND symb_decoder(16#3a#));
reg_q514_in <= (reg_q512 AND symb_decoder(16#5b#));
reg_q468_in <= (reg_q466 AND symb_decoder(16#41#)) OR
 					(reg_q466 AND symb_decoder(16#61#));
reg_q1902_in <= (reg_q1900 AND symb_decoder(16#54#)) OR
 					(reg_q1900 AND symb_decoder(16#74#));
reg_q28_in <= (reg_q26 AND symb_decoder(16#45#)) OR
 					(reg_q26 AND symb_decoder(16#65#));
reg_q30_in <= (reg_q28 AND symb_decoder(16#43#)) OR
 					(reg_q28 AND symb_decoder(16#63#));
reg_q917_in <= (reg_q915 AND symb_decoder(16#61#)) OR
 					(reg_q915 AND symb_decoder(16#41#));
reg_q2443_in <= (reg_q2441 AND symb_decoder(16#44#)) OR
 					(reg_q2441 AND symb_decoder(16#64#));
reg_q1808_in <= (reg_q1806 AND symb_decoder(16#52#)) OR
 					(reg_q1806 AND symb_decoder(16#72#));
reg_q1810_in <= (reg_q1808 AND symb_decoder(16#56#)) OR
 					(reg_q1808 AND symb_decoder(16#76#));
reg_q1369_in <= (reg_q1367 AND symb_decoder(16#78#)) OR
 					(reg_q1367 AND symb_decoder(16#58#));
reg_q588_in <= (reg_q586 AND symb_decoder(16#50#)) OR
 					(reg_q586 AND symb_decoder(16#70#));
reg_q1892_in <= (reg_q1890 AND symb_decoder(16#64#)) OR
 					(reg_q1890 AND symb_decoder(16#44#));
reg_q538_in <= (reg_q536 AND symb_decoder(16#25#));
reg_q1391_in <= (reg_q1389 AND symb_decoder(16#45#)) OR
 					(reg_q1389 AND symb_decoder(16#65#));
reg_q502_in <= (reg_q500 AND symb_decoder(16#4e#)) OR
 					(reg_q500 AND symb_decoder(16#6e#));
reg_q504_in <= (reg_q502 AND symb_decoder(16#45#)) OR
 					(reg_q502 AND symb_decoder(16#65#));
reg_q466_in <= (reg_q464 AND symb_decoder(16#45#)) OR
 					(reg_q464 AND symb_decoder(16#65#));
reg_q2463_in <= (reg_q2461 AND symb_decoder(16#46#)) OR
 					(reg_q2461 AND symb_decoder(16#66#));
reg_q2391_in <= (reg_q2389 AND symb_decoder(16#61#)) OR
 					(reg_q2389 AND symb_decoder(16#41#));
reg_q2325_in <= (reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2324 AND symb_decoder(16#22#));
reg_q26_in <= (reg_q24 AND symb_decoder(16#78#)) OR
 					(reg_q24 AND symb_decoder(16#58#));
reg_q903_in <= (reg_q901 AND symb_decoder(16#0d#));
reg_q518_in <= (reg_q516 AND symb_decoder(16#50#)) OR
 					(reg_q516 AND symb_decoder(16#70#));
reg_q1840_in <= (reg_q1838 AND symb_decoder(16#64#)) OR
 					(reg_q1838 AND symb_decoder(16#44#));
reg_q624_in <= (reg_q622 AND symb_decoder(16#52#)) OR
 					(reg_q622 AND symb_decoder(16#72#));
reg_q626_in <= (reg_q624 AND symb_decoder(16#56#)) OR
 					(reg_q624 AND symb_decoder(16#76#));
reg_q516_in <= (reg_q514 AND symb_decoder(16#49#)) OR
 					(reg_q514 AND symb_decoder(16#69#));
reg_q1946_in <= (reg_q1944 AND symb_decoder(16#77#)) OR
 					(reg_q1944 AND symb_decoder(16#57#));
reg_q1864_in <= (reg_q1862 AND symb_decoder(16#52#)) OR
 					(reg_q1862 AND symb_decoder(16#72#));
reg_q1940_in <= (reg_q1938 AND symb_decoder(16#73#)) OR
 					(reg_q1938 AND symb_decoder(16#53#));
reg_q42_in <= (reg_q40 AND symb_decoder(16#2e#));
reg_q44_in <= (reg_q42 AND symb_decoder(16#2e#));
reg_q2202_in <= (reg_q2200 AND symb_decoder(16#6d#)) OR
 					(reg_q2200 AND symb_decoder(16#4d#));
reg_q2520_in <= (reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2518 AND symb_decoder(16#2f#));
reg_q860_in <= (reg_q858 AND symb_decoder(16#56#)) OR
 					(reg_q858 AND symb_decoder(16#76#));
reg_q1031_in <= (reg_q1029 AND symb_decoder(16#69#)) OR
 					(reg_q1029 AND symb_decoder(16#49#));
reg_q2393_in <= (reg_q2391 AND symb_decoder(16#43#)) OR
 					(reg_q2391 AND symb_decoder(16#63#));
reg_q2204_in <= (reg_q2202 AND symb_decoder(16#4f#)) OR
 					(reg_q2202 AND symb_decoder(16#6f#));
reg_q2206_in <= (reg_q2204 AND symb_decoder(16#4e#)) OR
 					(reg_q2204 AND symb_decoder(16#6e#));
reg_q646_in <= (reg_q644 AND symb_decoder(16#25#));
reg_q2403_in <= (reg_q2401 AND symb_decoder(16#4f#)) OR
 					(reg_q2401 AND symb_decoder(16#6f#));
reg_q1952_in <= (reg_q1950 AND symb_decoder(16#45#)) OR
 					(reg_q1950 AND symb_decoder(16#65#));
reg_q1405_in <= (reg_q1403 AND symb_decoder(16#52#)) OR
 					(reg_q1403 AND symb_decoder(16#72#));
reg_q1407_in <= (reg_q1405 AND symb_decoder(16#70#)) OR
 					(reg_q1405 AND symb_decoder(16#50#));
reg_q622_in <= (reg_q620 AND symb_decoder(16#65#)) OR
 					(reg_q620 AND symb_decoder(16#45#));
reg_q488_in <= (reg_q486 AND symb_decoder(16#25#));
reg_q490_in <= (reg_q488 AND symb_decoder(16#32#));
reg_q40_in <= (reg_q38 AND symb_decoder(16#2e#));
reg_q654_in <= (reg_q652 AND symb_decoder(16#32#));
reg_q656_in <= (reg_q654 AND symb_decoder(16#31#));
reg_q570_in <= (reg_q568 AND symb_decoder(16#32#));
reg_q822_in <= (reg_q820 AND symb_decoder(16#69#)) OR
 					(reg_q820 AND symb_decoder(16#49#));
reg_q1363_in <= (reg_q1361 AND symb_decoder(16#30#));
reg_q2522_in <= (reg_q2520 AND symb_decoder(16#67#)) OR
 					(reg_q2520 AND symb_decoder(16#47#));
reg_q652_in <= (reg_q650 AND symb_decoder(16#25#));
reg_q1413_in <= (reg_q1411 AND symb_decoder(16#79#)) OR
 					(reg_q1411 AND symb_decoder(16#59#));
reg_q610_in <= (reg_q608 AND symb_decoder(16#25#));
reg_q536_in <= (reg_q534 AND symb_decoder(16#5d#));
reg_q2056_in <= (reg_q2054 AND symb_decoder(16#68#));
reg_q2058_in <= (reg_q2056 AND symb_decoder(16#65#));
reg_q660_in <= (reg_q658 AND symb_decoder(16#32#));
reg_q662_in <= (reg_q660 AND symb_decoder(16#31#));
reg_q2060_in <= (reg_q2058 AND symb_decoder(16#65#));
reg_q658_in <= (reg_q656 AND symb_decoder(16#25#));
reg_q2076_in <= (reg_q2074 AND symb_decoder(16#53#));
reg_fullgraph7_init <= "000000000";

reg_fullgraph7_sel <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & reg_q2076_in & reg_q658_in & reg_q2060_in & reg_q662_in & reg_q660_in & reg_q2058_in & reg_q2056_in & reg_q536_in & reg_q610_in & reg_q1413_in & reg_q652_in & reg_q2522_in & reg_q1363_in & reg_q822_in & reg_q570_in & reg_q656_in & reg_q654_in & reg_q40_in & reg_q490_in & reg_q488_in & reg_q622_in & reg_q1407_in & reg_q1405_in & reg_q1952_in & reg_q2403_in & reg_q646_in & reg_q2206_in & reg_q2204_in & reg_q2393_in & reg_q1031_in & reg_q860_in & reg_q2520_in & reg_q2202_in & reg_q44_in & reg_q42_in & reg_q1940_in & reg_q1864_in & reg_q1946_in & reg_q516_in & reg_q626_in & reg_q624_in & reg_q1840_in & reg_q518_in & reg_q903_in & reg_q26_in & reg_q2325_in & reg_q2391_in & reg_q2463_in & reg_q466_in & reg_q504_in & reg_q502_in & reg_q1391_in & reg_q538_in & reg_q1892_in & reg_q588_in & reg_q1369_in & reg_q1810_in & reg_q1808_in & reg_q2443_in & reg_q917_in & reg_q30_in & reg_q28_in & reg_q1902_in & reg_q468_in & reg_q514_in & reg_q2088_in & reg_q2086_in & reg_q550_in & reg_q486_in & reg_q484_in & reg_q736_in & reg_q1934_in & reg_q1203_in & reg_q1856_in & reg_q24_in & reg_q905_in & reg_q820_in & reg_q1896_in & reg_q1894_in & reg_q500_in & reg_q482_in & reg_q480_in & reg_q2508_in & reg_q470_in & reg_q544_in & reg_q1199_in & reg_q1379_in & reg_q1914_in & reg_q512_in & reg_q1932_in & reg_q1930_in & reg_q568_in & reg_q464_in & reg_q462_in & reg_q498_in & reg_q496_in & reg_q8_in & reg_q1900_in & reg_q1898_in & reg_q1838_in & reg_q2190_in & reg_q2084_in & reg_q2082_in & reg_q602_in & reg_q494_in & reg_q492_in & reg_q582_in & reg_q2493_in & reg_q548_in & reg_q546_in & reg_q472_in & reg_q1806_in & reg_q1804_in & reg_q560_in & reg_q2413_in & reg_q2437_in & reg_q2435_in & reg_q20_in & reg_q576_in & reg_q586_in & reg_q584_in & reg_q1908_in & reg_q2401_in & reg_q2399_in & reg_q1371_in & reg_q1812_in & reg_q1367_in & reg_q1365_in & reg_q554_in & reg_q552_in & reg_q636_in & reg_q2489_in & reg_q2487_in & reg_q644_in & reg_q642_in & reg_q1928_in & reg_q1399_in & reg_q870_in & reg_q868_in & reg_q866_in & reg_q2468_in & reg_q872_in & reg_q32_in & reg_q594_in & reg_q640_in & reg_q638_in & reg_q2524_in & reg_q1161_in & reg_q862_in & reg_q574_in & reg_q572_in & reg_q941_in & reg_q2200_in & reg_q1936_in & reg_q1798_in & reg_q542_in & reg_q540_in & reg_q1846_in & reg_q2162_in & reg_q2188_in & reg_q2186_in & reg_q1872_in & reg_q1983_in & reg_q1113_in & reg_q1830_in & reg_q789_in & reg_q1397_in & reg_q2192_in & reg_q1824_in & reg_q1822_in & reg_q650_in & reg_q648_in & reg_q1796_in & reg_q1219_in & reg_q805_in & reg_q524_in & reg_q478_in & reg_q809_in & reg_q807_in & reg_q803_in & reg_q1993_in & reg_q1991_in & reg_q1870_in & reg_q1550_in & reg_q1922_in & reg_q1862_in & reg_q787_in & reg_q1464_in & reg_q878_in & reg_q1525_in & reg_q1836_in & reg_q1860_in & reg_q1858_in & reg_q1213_in & reg_q634_in & reg_q1944_in & reg_q1942_in & reg_q943_in & reg_q564_in & reg_q562_in & reg_q1814_in & reg_q510_in & reg_q797_in & reg_q795_in & reg_q1979_in & reg_q14_in & reg_q1605_in & reg_q1950_in & reg_q1948_in & reg_q1381_in & reg_q131_in & reg_q628_in & reg_q508_in & reg_q506_in & reg_q1646_in & reg_q18_in & reg_q1844_in & reg_q1842_in & reg_q1820_in & reg_q1818_in & reg_q580_in & reg_q578_in & reg_q1912_in & reg_q1910_in & reg_q2415_in & reg_q801_in & reg_q799_in & reg_q1834_in & reg_q1832_in & reg_q1989_in & reg_q1987_in & reg_q2433_in & reg_q2431_in & reg_q608_in & reg_q606_in & reg_q530_in & reg_q528_in & reg_q1890_in & reg_q1888_in & reg_q1850_in & reg_q630_in & reg_q2441_in & reg_q2439_in & reg_q1924_in & reg_q1205_in & reg_q2397_in & reg_q2395_in & reg_q476_in & reg_q474_in & reg_q1393_in & reg_q2062_in & reg_q1981_in & reg_q600_in & reg_q598_in & reg_q2184_in & reg_q2182_in & reg_q758_in & reg_q2093_in & reg_q1226_in & reg_q1800_in & reg_q1916_in & reg_q38_in & reg_q1403_in & reg_q1401_in & reg_q1985_in & reg_q1207_in & reg_q884_in & reg_q2072_in & reg_q36_in & reg_q34_in & reg_q614_in & reg_q612_in & reg_q854_in & reg_q2198_in & reg_q2196_in & reg_q2425_in & reg_q2423_in & reg_q2526_in & reg_q2429_in & reg_q882_in & reg_q2409_in & reg_q12_in & reg_q951_in & reg_q949_in & reg_q876_in & reg_q874_in & reg_q960_in & reg_q2064_in & reg_q1411_in & reg_q1409_in & reg_q1920_in & reg_q2407_in & reg_q2405_in & reg_q1389_in & reg_q1387_in & reg_q592_in & reg_q590_in & reg_q2180_in & reg_q2178_in & reg_q2080_in & reg_q2078_in & reg_q1874_in & reg_q2447_in & reg_q2445_in & reg_q2530_in & reg_q2528_in & reg_q522_in & reg_q520_in & reg_q2002_in & reg_q1866_in & reg_q939_in & reg_q937_in & reg_q1217_in & reg_q1215_in & reg_q858_in & reg_q856_in & reg_q791_in & reg_q947_in & reg_q945_in & reg_q526_in & reg_q616_in & reg_q1770_in & reg_q2421_in & reg_q2419_in & reg_q534_in & reg_q532_in & reg_q889_in & reg_q1854_in & reg_q1852_in & reg_q1794_in & reg_q1792_in & reg_q1878_in & reg_q1876_in;

	--coder fullgraph7
with reg_fullgraph7_sel select
reg_fullgraph7_in <=
	"000000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001",
	"000000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010",
	"000000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100",
	"000000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000",
	"000000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000",
	"000000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000",
	"000000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000",
	"000001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000",
	"000001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
	"000001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000",
	"000001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000",
	"000001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000",
	"000001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000",
	"000001110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000",
	"000001111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000",
	"000010000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000",
	"000010001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000",
	"000010010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000",
	"000010011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000",
	"000010100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000",
	"000010101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000",
	"000010110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000",
	"000010111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000",
	"000011000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000",
	"000011001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000",
	"000011010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000",
	"000011011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000",
	"000011100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000",
	"000011101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000",
	"000011110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000",
	"000011111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000",
	"000100000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000",
	"000100001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000",
	"000100010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000",
	"000100011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000",
	"000100100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000",
	"000100101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000",
	"000100110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000",
	"000100111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000",
	"000101000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000",
	"000101001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000",
	"000101010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000",
	"000101011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000",
	"000101100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000",
	"000101101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
	"000101110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000",
	"000101111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000",
	"000110000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000",
	"000110001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000",
	"000110010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000",
	"000110011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000",
	"000110100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000",
	"000110101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000",
	"000110110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000",
	"000110111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000",
	"000111000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000",
	"000111001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000",
	"000111010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000",
	"000111011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000",
	"000111100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000",
	"000111101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000",
	"000111110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000",
	"000111111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000",
	"001000000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000",
	"001000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000",
	"001000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000",
	"001000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000",
	"001000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000",
	"001000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000",
	"001000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000",
	"001000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000",
	"001001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000",
	"001001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000",
	"001001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000",
	"001001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000",
	"001001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001001110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001001111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001010111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001011111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001100111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001101111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001110111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"001111111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010001111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010010111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010011111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010100111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010101111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010110111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"010111111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011001111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011010111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011011111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011100111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011101111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011110111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"011111111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100001111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100010111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100011111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100100111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100101111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100110111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"100111111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000110" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101000111" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001000" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001001" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001010" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001011" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001100" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"101001101" when "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	"000000000" when others;
 --end coder

	p_reg_fullgraph7: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph7 <= reg_fullgraph7_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph7 <= reg_fullgraph7_init;
        else
          reg_fullgraph7 <= reg_fullgraph7_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph7

		reg_q1876 <= '1' when reg_fullgraph7 = "000000001" else '0'; 
		reg_q1878 <= '1' when reg_fullgraph7 = "000000010" else '0'; 
		reg_q1792 <= '1' when reg_fullgraph7 = "000000011" else '0'; 
		reg_q1794 <= '1' when reg_fullgraph7 = "000000100" else '0'; 
		reg_q1852 <= '1' when reg_fullgraph7 = "000000101" else '0'; 
		reg_q1854 <= '1' when reg_fullgraph7 = "000000110" else '0'; 
		reg_q889 <= '1' when reg_fullgraph7 = "000000111" else '0'; 
		reg_q532 <= '1' when reg_fullgraph7 = "000001000" else '0'; 
		reg_q534 <= '1' when reg_fullgraph7 = "000001001" else '0'; 
		reg_q2419 <= '1' when reg_fullgraph7 = "000001010" else '0'; 
		reg_q2421 <= '1' when reg_fullgraph7 = "000001011" else '0'; 
		reg_q1770 <= '1' when reg_fullgraph7 = "000001100" else '0'; 
		reg_q616 <= '1' when reg_fullgraph7 = "000001101" else '0'; 
		reg_q526 <= '1' when reg_fullgraph7 = "000001110" else '0'; 
		reg_q945 <= '1' when reg_fullgraph7 = "000001111" else '0'; 
		reg_q947 <= '1' when reg_fullgraph7 = "000010000" else '0'; 
		reg_q791 <= '1' when reg_fullgraph7 = "000010001" else '0'; 
		reg_q856 <= '1' when reg_fullgraph7 = "000010010" else '0'; 
		reg_q858 <= '1' when reg_fullgraph7 = "000010011" else '0'; 
		reg_q1215 <= '1' when reg_fullgraph7 = "000010100" else '0'; 
		reg_q1217 <= '1' when reg_fullgraph7 = "000010101" else '0'; 
		reg_q937 <= '1' when reg_fullgraph7 = "000010110" else '0'; 
		reg_q939 <= '1' when reg_fullgraph7 = "000010111" else '0'; 
		reg_q1866 <= '1' when reg_fullgraph7 = "000011000" else '0'; 
		reg_q2002 <= '1' when reg_fullgraph7 = "000011001" else '0'; 
		reg_q520 <= '1' when reg_fullgraph7 = "000011010" else '0'; 
		reg_q522 <= '1' when reg_fullgraph7 = "000011011" else '0'; 
		reg_q2528 <= '1' when reg_fullgraph7 = "000011100" else '0'; 
		reg_q2530 <= '1' when reg_fullgraph7 = "000011101" else '0'; 
		reg_q2445 <= '1' when reg_fullgraph7 = "000011110" else '0'; 
		reg_q2447 <= '1' when reg_fullgraph7 = "000011111" else '0'; 
		reg_q1874 <= '1' when reg_fullgraph7 = "000100000" else '0'; 
		reg_q2078 <= '1' when reg_fullgraph7 = "000100001" else '0'; 
		reg_q2080 <= '1' when reg_fullgraph7 = "000100010" else '0'; 
		reg_q2178 <= '1' when reg_fullgraph7 = "000100011" else '0'; 
		reg_q2180 <= '1' when reg_fullgraph7 = "000100100" else '0'; 
		reg_q590 <= '1' when reg_fullgraph7 = "000100101" else '0'; 
		reg_q592 <= '1' when reg_fullgraph7 = "000100110" else '0'; 
		reg_q1387 <= '1' when reg_fullgraph7 = "000100111" else '0'; 
		reg_q1389 <= '1' when reg_fullgraph7 = "000101000" else '0'; 
		reg_q2405 <= '1' when reg_fullgraph7 = "000101001" else '0'; 
		reg_q2407 <= '1' when reg_fullgraph7 = "000101010" else '0'; 
		reg_q1920 <= '1' when reg_fullgraph7 = "000101011" else '0'; 
		reg_q1409 <= '1' when reg_fullgraph7 = "000101100" else '0'; 
		reg_q1411 <= '1' when reg_fullgraph7 = "000101101" else '0'; 
		reg_q2064 <= '1' when reg_fullgraph7 = "000101110" else '0'; 
		reg_q960 <= '1' when reg_fullgraph7 = "000101111" else '0'; 
		reg_q874 <= '1' when reg_fullgraph7 = "000110000" else '0'; 
		reg_q876 <= '1' when reg_fullgraph7 = "000110001" else '0'; 
		reg_q949 <= '1' when reg_fullgraph7 = "000110010" else '0'; 
		reg_q951 <= '1' when reg_fullgraph7 = "000110011" else '0'; 
		reg_q12 <= '1' when reg_fullgraph7 = "000110100" else '0'; 
		reg_q2409 <= '1' when reg_fullgraph7 = "000110101" else '0'; 
		reg_q882 <= '1' when reg_fullgraph7 = "000110110" else '0'; 
		reg_q2429 <= '1' when reg_fullgraph7 = "000110111" else '0'; 
		reg_q2526 <= '1' when reg_fullgraph7 = "000111000" else '0'; 
		reg_q2423 <= '1' when reg_fullgraph7 = "000111001" else '0'; 
		reg_q2425 <= '1' when reg_fullgraph7 = "000111010" else '0'; 
		reg_q2196 <= '1' when reg_fullgraph7 = "000111011" else '0'; 
		reg_q2198 <= '1' when reg_fullgraph7 = "000111100" else '0'; 
		reg_q854 <= '1' when reg_fullgraph7 = "000111101" else '0'; 
		reg_q612 <= '1' when reg_fullgraph7 = "000111110" else '0'; 
		reg_q614 <= '1' when reg_fullgraph7 = "000111111" else '0'; 
		reg_q34 <= '1' when reg_fullgraph7 = "001000000" else '0'; 
		reg_q36 <= '1' when reg_fullgraph7 = "001000001" else '0'; 
		reg_q2072 <= '1' when reg_fullgraph7 = "001000010" else '0'; 
		reg_q884 <= '1' when reg_fullgraph7 = "001000011" else '0'; 
		reg_q1207 <= '1' when reg_fullgraph7 = "001000100" else '0'; 
		reg_q1985 <= '1' when reg_fullgraph7 = "001000101" else '0'; 
		reg_q1401 <= '1' when reg_fullgraph7 = "001000110" else '0'; 
		reg_q1403 <= '1' when reg_fullgraph7 = "001000111" else '0'; 
		reg_q38 <= '1' when reg_fullgraph7 = "001001000" else '0'; 
		reg_q1916 <= '1' when reg_fullgraph7 = "001001001" else '0'; 
		reg_q1800 <= '1' when reg_fullgraph7 = "001001010" else '0'; 
		reg_q1226 <= '1' when reg_fullgraph7 = "001001011" else '0'; 
		reg_q2093 <= '1' when reg_fullgraph7 = "001001100" else '0'; 
		reg_q758 <= '1' when reg_fullgraph7 = "001001101" else '0'; 
		reg_q2182 <= '1' when reg_fullgraph7 = "001001110" else '0'; 
		reg_q2184 <= '1' when reg_fullgraph7 = "001001111" else '0'; 
		reg_q598 <= '1' when reg_fullgraph7 = "001010000" else '0'; 
		reg_q600 <= '1' when reg_fullgraph7 = "001010001" else '0'; 
		reg_q1981 <= '1' when reg_fullgraph7 = "001010010" else '0'; 
		reg_q2062 <= '1' when reg_fullgraph7 = "001010011" else '0'; 
		reg_q1393 <= '1' when reg_fullgraph7 = "001010100" else '0'; 
		reg_q474 <= '1' when reg_fullgraph7 = "001010101" else '0'; 
		reg_q476 <= '1' when reg_fullgraph7 = "001010110" else '0'; 
		reg_q2395 <= '1' when reg_fullgraph7 = "001010111" else '0'; 
		reg_q2397 <= '1' when reg_fullgraph7 = "001011000" else '0'; 
		reg_q1205 <= '1' when reg_fullgraph7 = "001011001" else '0'; 
		reg_q1924 <= '1' when reg_fullgraph7 = "001011010" else '0'; 
		reg_q2439 <= '1' when reg_fullgraph7 = "001011011" else '0'; 
		reg_q2441 <= '1' when reg_fullgraph7 = "001011100" else '0'; 
		reg_q630 <= '1' when reg_fullgraph7 = "001011101" else '0'; 
		reg_q1850 <= '1' when reg_fullgraph7 = "001011110" else '0'; 
		reg_q1888 <= '1' when reg_fullgraph7 = "001011111" else '0'; 
		reg_q1890 <= '1' when reg_fullgraph7 = "001100000" else '0'; 
		reg_q528 <= '1' when reg_fullgraph7 = "001100001" else '0'; 
		reg_q530 <= '1' when reg_fullgraph7 = "001100010" else '0'; 
		reg_q606 <= '1' when reg_fullgraph7 = "001100011" else '0'; 
		reg_q608 <= '1' when reg_fullgraph7 = "001100100" else '0'; 
		reg_q2431 <= '1' when reg_fullgraph7 = "001100101" else '0'; 
		reg_q2433 <= '1' when reg_fullgraph7 = "001100110" else '0'; 
		reg_q1987 <= '1' when reg_fullgraph7 = "001100111" else '0'; 
		reg_q1989 <= '1' when reg_fullgraph7 = "001101000" else '0'; 
		reg_q1832 <= '1' when reg_fullgraph7 = "001101001" else '0'; 
		reg_q1834 <= '1' when reg_fullgraph7 = "001101010" else '0'; 
		reg_q799 <= '1' when reg_fullgraph7 = "001101011" else '0'; 
		reg_q801 <= '1' when reg_fullgraph7 = "001101100" else '0'; 
		reg_q2415 <= '1' when reg_fullgraph7 = "001101101" else '0'; 
		reg_q1910 <= '1' when reg_fullgraph7 = "001101110" else '0'; 
		reg_q1912 <= '1' when reg_fullgraph7 = "001101111" else '0'; 
		reg_q578 <= '1' when reg_fullgraph7 = "001110000" else '0'; 
		reg_q580 <= '1' when reg_fullgraph7 = "001110001" else '0'; 
		reg_q1818 <= '1' when reg_fullgraph7 = "001110010" else '0'; 
		reg_q1820 <= '1' when reg_fullgraph7 = "001110011" else '0'; 
		reg_q1842 <= '1' when reg_fullgraph7 = "001110100" else '0'; 
		reg_q1844 <= '1' when reg_fullgraph7 = "001110101" else '0'; 
		reg_q18 <= '1' when reg_fullgraph7 = "001110110" else '0'; 
		reg_q1646 <= '1' when reg_fullgraph7 = "001110111" else '0'; 
		reg_q506 <= '1' when reg_fullgraph7 = "001111000" else '0'; 
		reg_q508 <= '1' when reg_fullgraph7 = "001111001" else '0'; 
		reg_q628 <= '1' when reg_fullgraph7 = "001111010" else '0'; 
		reg_q131 <= '1' when reg_fullgraph7 = "001111011" else '0'; 
		reg_q1381 <= '1' when reg_fullgraph7 = "001111100" else '0'; 
		reg_q1948 <= '1' when reg_fullgraph7 = "001111101" else '0'; 
		reg_q1950 <= '1' when reg_fullgraph7 = "001111110" else '0'; 
		reg_q1605 <= '1' when reg_fullgraph7 = "001111111" else '0'; 
		reg_q14 <= '1' when reg_fullgraph7 = "010000000" else '0'; 
		reg_q1979 <= '1' when reg_fullgraph7 = "010000001" else '0'; 
		reg_q795 <= '1' when reg_fullgraph7 = "010000010" else '0'; 
		reg_q797 <= '1' when reg_fullgraph7 = "010000011" else '0'; 
		reg_q510 <= '1' when reg_fullgraph7 = "010000100" else '0'; 
		reg_q1814 <= '1' when reg_fullgraph7 = "010000101" else '0'; 
		reg_q562 <= '1' when reg_fullgraph7 = "010000110" else '0'; 
		reg_q564 <= '1' when reg_fullgraph7 = "010000111" else '0'; 
		reg_q943 <= '1' when reg_fullgraph7 = "010001000" else '0'; 
		reg_q1942 <= '1' when reg_fullgraph7 = "010001001" else '0'; 
		reg_q1944 <= '1' when reg_fullgraph7 = "010001010" else '0'; 
		reg_q634 <= '1' when reg_fullgraph7 = "010001011" else '0'; 
		reg_q1213 <= '1' when reg_fullgraph7 = "010001100" else '0'; 
		reg_q1858 <= '1' when reg_fullgraph7 = "010001101" else '0'; 
		reg_q1860 <= '1' when reg_fullgraph7 = "010001110" else '0'; 
		reg_q1836 <= '1' when reg_fullgraph7 = "010001111" else '0'; 
		reg_q1525 <= '1' when reg_fullgraph7 = "010010000" else '0'; 
		reg_q878 <= '1' when reg_fullgraph7 = "010010001" else '0'; 
		reg_q1464 <= '1' when reg_fullgraph7 = "010010010" else '0'; 
		reg_q787 <= '1' when reg_fullgraph7 = "010010011" else '0'; 
		reg_q1862 <= '1' when reg_fullgraph7 = "010010100" else '0'; 
		reg_q1922 <= '1' when reg_fullgraph7 = "010010101" else '0'; 
		reg_q1550 <= '1' when reg_fullgraph7 = "010010110" else '0'; 
		reg_q1870 <= '1' when reg_fullgraph7 = "010010111" else '0'; 
		reg_q1991 <= '1' when reg_fullgraph7 = "010011000" else '0'; 
		reg_q1993 <= '1' when reg_fullgraph7 = "010011001" else '0'; 
		reg_q803 <= '1' when reg_fullgraph7 = "010011010" else '0'; 
		reg_q807 <= '1' when reg_fullgraph7 = "010011011" else '0'; 
		reg_q809 <= '1' when reg_fullgraph7 = "010011100" else '0'; 
		reg_q478 <= '1' when reg_fullgraph7 = "010011101" else '0'; 
		reg_q524 <= '1' when reg_fullgraph7 = "010011110" else '0'; 
		reg_q805 <= '1' when reg_fullgraph7 = "010011111" else '0'; 
		reg_q1219 <= '1' when reg_fullgraph7 = "010100000" else '0'; 
		reg_q1796 <= '1' when reg_fullgraph7 = "010100001" else '0'; 
		reg_q648 <= '1' when reg_fullgraph7 = "010100010" else '0'; 
		reg_q650 <= '1' when reg_fullgraph7 = "010100011" else '0'; 
		reg_q1822 <= '1' when reg_fullgraph7 = "010100100" else '0'; 
		reg_q1824 <= '1' when reg_fullgraph7 = "010100101" else '0'; 
		reg_q2192 <= '1' when reg_fullgraph7 = "010100110" else '0'; 
		reg_q1397 <= '1' when reg_fullgraph7 = "010100111" else '0'; 
		reg_q789 <= '1' when reg_fullgraph7 = "010101000" else '0'; 
		reg_q1830 <= '1' when reg_fullgraph7 = "010101001" else '0'; 
		reg_q1113 <= '1' when reg_fullgraph7 = "010101010" else '0'; 
		reg_q1983 <= '1' when reg_fullgraph7 = "010101011" else '0'; 
		reg_q1872 <= '1' when reg_fullgraph7 = "010101100" else '0'; 
		reg_q2186 <= '1' when reg_fullgraph7 = "010101101" else '0'; 
		reg_q2188 <= '1' when reg_fullgraph7 = "010101110" else '0'; 
		reg_q2162 <= '1' when reg_fullgraph7 = "010101111" else '0'; 
		reg_q1846 <= '1' when reg_fullgraph7 = "010110000" else '0'; 
		reg_q540 <= '1' when reg_fullgraph7 = "010110001" else '0'; 
		reg_q542 <= '1' when reg_fullgraph7 = "010110010" else '0'; 
		reg_q1798 <= '1' when reg_fullgraph7 = "010110011" else '0'; 
		reg_q1936 <= '1' when reg_fullgraph7 = "010110100" else '0'; 
		reg_q2200 <= '1' when reg_fullgraph7 = "010110101" else '0'; 
		reg_q941 <= '1' when reg_fullgraph7 = "010110110" else '0'; 
		reg_q572 <= '1' when reg_fullgraph7 = "010110111" else '0'; 
		reg_q574 <= '1' when reg_fullgraph7 = "010111000" else '0'; 
		reg_q862 <= '1' when reg_fullgraph7 = "010111001" else '0'; 
		reg_q1161 <= '1' when reg_fullgraph7 = "010111010" else '0'; 
		reg_q2524 <= '1' when reg_fullgraph7 = "010111011" else '0'; 
		reg_q638 <= '1' when reg_fullgraph7 = "010111100" else '0'; 
		reg_q640 <= '1' when reg_fullgraph7 = "010111101" else '0'; 
		reg_q594 <= '1' when reg_fullgraph7 = "010111110" else '0'; 
		reg_q32 <= '1' when reg_fullgraph7 = "010111111" else '0'; 
		reg_q872 <= '1' when reg_fullgraph7 = "011000000" else '0'; 
		reg_q2468 <= '1' when reg_fullgraph7 = "011000001" else '0'; 
		reg_q866 <= '1' when reg_fullgraph7 = "011000010" else '0'; 
		reg_q868 <= '1' when reg_fullgraph7 = "011000011" else '0'; 
		reg_q870 <= '1' when reg_fullgraph7 = "011000100" else '0'; 
		reg_q1399 <= '1' when reg_fullgraph7 = "011000101" else '0'; 
		reg_q1928 <= '1' when reg_fullgraph7 = "011000110" else '0'; 
		reg_q642 <= '1' when reg_fullgraph7 = "011000111" else '0'; 
		reg_q644 <= '1' when reg_fullgraph7 = "011001000" else '0'; 
		reg_q2487 <= '1' when reg_fullgraph7 = "011001001" else '0'; 
		reg_q2489 <= '1' when reg_fullgraph7 = "011001010" else '0'; 
		reg_q636 <= '1' when reg_fullgraph7 = "011001011" else '0'; 
		reg_q552 <= '1' when reg_fullgraph7 = "011001100" else '0'; 
		reg_q554 <= '1' when reg_fullgraph7 = "011001101" else '0'; 
		reg_q1365 <= '1' when reg_fullgraph7 = "011001110" else '0'; 
		reg_q1367 <= '1' when reg_fullgraph7 = "011001111" else '0'; 
		reg_q1812 <= '1' when reg_fullgraph7 = "011010000" else '0'; 
		reg_q1371 <= '1' when reg_fullgraph7 = "011010001" else '0'; 
		reg_q2399 <= '1' when reg_fullgraph7 = "011010010" else '0'; 
		reg_q2401 <= '1' when reg_fullgraph7 = "011010011" else '0'; 
		reg_q1908 <= '1' when reg_fullgraph7 = "011010100" else '0'; 
		reg_q584 <= '1' when reg_fullgraph7 = "011010101" else '0'; 
		reg_q586 <= '1' when reg_fullgraph7 = "011010110" else '0'; 
		reg_q576 <= '1' when reg_fullgraph7 = "011010111" else '0'; 
		reg_q20 <= '1' when reg_fullgraph7 = "011011000" else '0'; 
		reg_q2435 <= '1' when reg_fullgraph7 = "011011001" else '0'; 
		reg_q2437 <= '1' when reg_fullgraph7 = "011011010" else '0'; 
		reg_q2413 <= '1' when reg_fullgraph7 = "011011011" else '0'; 
		reg_q560 <= '1' when reg_fullgraph7 = "011011100" else '0'; 
		reg_q1804 <= '1' when reg_fullgraph7 = "011011101" else '0'; 
		reg_q1806 <= '1' when reg_fullgraph7 = "011011110" else '0'; 
		reg_q472 <= '1' when reg_fullgraph7 = "011011111" else '0'; 
		reg_q546 <= '1' when reg_fullgraph7 = "011100000" else '0'; 
		reg_q548 <= '1' when reg_fullgraph7 = "011100001" else '0'; 
		reg_q2493 <= '1' when reg_fullgraph7 = "011100010" else '0'; 
		reg_q582 <= '1' when reg_fullgraph7 = "011100011" else '0'; 
		reg_q492 <= '1' when reg_fullgraph7 = "011100100" else '0'; 
		reg_q494 <= '1' when reg_fullgraph7 = "011100101" else '0'; 
		reg_q602 <= '1' when reg_fullgraph7 = "011100110" else '0'; 
		reg_q2082 <= '1' when reg_fullgraph7 = "011100111" else '0'; 
		reg_q2084 <= '1' when reg_fullgraph7 = "011101000" else '0'; 
		reg_q2190 <= '1' when reg_fullgraph7 = "011101001" else '0'; 
		reg_q1838 <= '1' when reg_fullgraph7 = "011101010" else '0'; 
		reg_q1898 <= '1' when reg_fullgraph7 = "011101011" else '0'; 
		reg_q1900 <= '1' when reg_fullgraph7 = "011101100" else '0'; 
		reg_q8 <= '1' when reg_fullgraph7 = "011101101" else '0'; 
		reg_q496 <= '1' when reg_fullgraph7 = "011101110" else '0'; 
		reg_q498 <= '1' when reg_fullgraph7 = "011101111" else '0'; 
		reg_q462 <= '1' when reg_fullgraph7 = "011110000" else '0'; 
		reg_q464 <= '1' when reg_fullgraph7 = "011110001" else '0'; 
		reg_q568 <= '1' when reg_fullgraph7 = "011110010" else '0'; 
		reg_q1930 <= '1' when reg_fullgraph7 = "011110011" else '0'; 
		reg_q1932 <= '1' when reg_fullgraph7 = "011110100" else '0'; 
		reg_q512 <= '1' when reg_fullgraph7 = "011110101" else '0'; 
		reg_q1914 <= '1' when reg_fullgraph7 = "011110110" else '0'; 
		reg_q1379 <= '1' when reg_fullgraph7 = "011110111" else '0'; 
		reg_q1199 <= '1' when reg_fullgraph7 = "011111000" else '0'; 
		reg_q544 <= '1' when reg_fullgraph7 = "011111001" else '0'; 
		reg_q470 <= '1' when reg_fullgraph7 = "011111010" else '0'; 
		reg_q2508 <= '1' when reg_fullgraph7 = "011111011" else '0'; 
		reg_q480 <= '1' when reg_fullgraph7 = "011111100" else '0'; 
		reg_q482 <= '1' when reg_fullgraph7 = "011111101" else '0'; 
		reg_q500 <= '1' when reg_fullgraph7 = "011111110" else '0'; 
		reg_q1894 <= '1' when reg_fullgraph7 = "011111111" else '0'; 
		reg_q1896 <= '1' when reg_fullgraph7 = "100000000" else '0'; 
		reg_q820 <= '1' when reg_fullgraph7 = "100000001" else '0'; 
		reg_q905 <= '1' when reg_fullgraph7 = "100000010" else '0'; 
		reg_q24 <= '1' when reg_fullgraph7 = "100000011" else '0'; 
		reg_q1856 <= '1' when reg_fullgraph7 = "100000100" else '0'; 
		reg_q1203 <= '1' when reg_fullgraph7 = "100000101" else '0'; 
		reg_q1934 <= '1' when reg_fullgraph7 = "100000110" else '0'; 
		reg_q736 <= '1' when reg_fullgraph7 = "100000111" else '0'; 
		reg_q484 <= '1' when reg_fullgraph7 = "100001000" else '0'; 
		reg_q486 <= '1' when reg_fullgraph7 = "100001001" else '0'; 
		reg_q550 <= '1' when reg_fullgraph7 = "100001010" else '0'; 
		reg_q2086 <= '1' when reg_fullgraph7 = "100001011" else '0'; 
		reg_q2088 <= '1' when reg_fullgraph7 = "100001100" else '0'; 
		reg_q514 <= '1' when reg_fullgraph7 = "100001101" else '0'; 
		reg_q468 <= '1' when reg_fullgraph7 = "100001110" else '0'; 
		reg_q1902 <= '1' when reg_fullgraph7 = "100001111" else '0'; 
		reg_q28 <= '1' when reg_fullgraph7 = "100010000" else '0'; 
		reg_q30 <= '1' when reg_fullgraph7 = "100010001" else '0'; 
		reg_q917 <= '1' when reg_fullgraph7 = "100010010" else '0'; 
		reg_q2443 <= '1' when reg_fullgraph7 = "100010011" else '0'; 
		reg_q1808 <= '1' when reg_fullgraph7 = "100010100" else '0'; 
		reg_q1810 <= '1' when reg_fullgraph7 = "100010101" else '0'; 
		reg_q1369 <= '1' when reg_fullgraph7 = "100010110" else '0'; 
		reg_q588 <= '1' when reg_fullgraph7 = "100010111" else '0'; 
		reg_q1892 <= '1' when reg_fullgraph7 = "100011000" else '0'; 
		reg_q538 <= '1' when reg_fullgraph7 = "100011001" else '0'; 
		reg_q1391 <= '1' when reg_fullgraph7 = "100011010" else '0'; 
		reg_q502 <= '1' when reg_fullgraph7 = "100011011" else '0'; 
		reg_q504 <= '1' when reg_fullgraph7 = "100011100" else '0'; 
		reg_q466 <= '1' when reg_fullgraph7 = "100011101" else '0'; 
		reg_q2463 <= '1' when reg_fullgraph7 = "100011110" else '0'; 
		reg_q2391 <= '1' when reg_fullgraph7 = "100011111" else '0'; 
		reg_q2325 <= '1' when reg_fullgraph7 = "100100000" else '0'; 
		reg_q26 <= '1' when reg_fullgraph7 = "100100001" else '0'; 
		reg_q903 <= '1' when reg_fullgraph7 = "100100010" else '0'; 
		reg_q518 <= '1' when reg_fullgraph7 = "100100011" else '0'; 
		reg_q1840 <= '1' when reg_fullgraph7 = "100100100" else '0'; 
		reg_q624 <= '1' when reg_fullgraph7 = "100100101" else '0'; 
		reg_q626 <= '1' when reg_fullgraph7 = "100100110" else '0'; 
		reg_q516 <= '1' when reg_fullgraph7 = "100100111" else '0'; 
		reg_q1946 <= '1' when reg_fullgraph7 = "100101000" else '0'; 
		reg_q1864 <= '1' when reg_fullgraph7 = "100101001" else '0'; 
		reg_q1940 <= '1' when reg_fullgraph7 = "100101010" else '0'; 
		reg_q42 <= '1' when reg_fullgraph7 = "100101011" else '0'; 
		reg_q44 <= '1' when reg_fullgraph7 = "100101100" else '0'; 
		reg_q2202 <= '1' when reg_fullgraph7 = "100101101" else '0'; 
		reg_q2520 <= '1' when reg_fullgraph7 = "100101110" else '0'; 
		reg_q860 <= '1' when reg_fullgraph7 = "100101111" else '0'; 
		reg_q1031 <= '1' when reg_fullgraph7 = "100110000" else '0'; 
		reg_q2393 <= '1' when reg_fullgraph7 = "100110001" else '0'; 
		reg_q2204 <= '1' when reg_fullgraph7 = "100110010" else '0'; 
		reg_q2206 <= '1' when reg_fullgraph7 = "100110011" else '0'; 
		reg_q646 <= '1' when reg_fullgraph7 = "100110100" else '0'; 
		reg_q2403 <= '1' when reg_fullgraph7 = "100110101" else '0'; 
		reg_q1952 <= '1' when reg_fullgraph7 = "100110110" else '0'; 
		reg_q1405 <= '1' when reg_fullgraph7 = "100110111" else '0'; 
		reg_q1407 <= '1' when reg_fullgraph7 = "100111000" else '0'; 
		reg_q622 <= '1' when reg_fullgraph7 = "100111001" else '0'; 
		reg_q488 <= '1' when reg_fullgraph7 = "100111010" else '0'; 
		reg_q490 <= '1' when reg_fullgraph7 = "100111011" else '0'; 
		reg_q40 <= '1' when reg_fullgraph7 = "100111100" else '0'; 
		reg_q654 <= '1' when reg_fullgraph7 = "100111101" else '0'; 
		reg_q656 <= '1' when reg_fullgraph7 = "100111110" else '0'; 
		reg_q570 <= '1' when reg_fullgraph7 = "100111111" else '0'; 
		reg_q822 <= '1' when reg_fullgraph7 = "101000000" else '0'; 
		reg_q1363 <= '1' when reg_fullgraph7 = "101000001" else '0'; 
		reg_q2522 <= '1' when reg_fullgraph7 = "101000010" else '0'; 
		reg_q652 <= '1' when reg_fullgraph7 = "101000011" else '0'; 
		reg_q1413 <= '1' when reg_fullgraph7 = "101000100" else '0'; 
		reg_q610 <= '1' when reg_fullgraph7 = "101000101" else '0'; 
		reg_q536 <= '1' when reg_fullgraph7 = "101000110" else '0'; 
		reg_q2056 <= '1' when reg_fullgraph7 = "101000111" else '0'; 
		reg_q2058 <= '1' when reg_fullgraph7 = "101001000" else '0'; 
		reg_q660 <= '1' when reg_fullgraph7 = "101001001" else '0'; 
		reg_q662 <= '1' when reg_fullgraph7 = "101001010" else '0'; 
		reg_q2060 <= '1' when reg_fullgraph7 = "101001011" else '0'; 
		reg_q658 <= '1' when reg_fullgraph7 = "101001100" else '0'; 
		reg_q2076 <= '1' when reg_fullgraph7 = "101001101" else '0'; 
--end decoder 

reg_q0_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q0 AND symb_decoder(16#a2#)) OR
 					(reg_q0 AND symb_decoder(16#08#)) OR
 					(reg_q0 AND symb_decoder(16#d3#)) OR
 					(reg_q0 AND symb_decoder(16#79#)) OR
 					(reg_q0 AND symb_decoder(16#6f#)) OR
 					(reg_q0 AND symb_decoder(16#8b#)) OR
 					(reg_q0 AND symb_decoder(16#01#)) OR
 					(reg_q0 AND symb_decoder(16#a5#)) OR
 					(reg_q0 AND symb_decoder(16#9a#)) OR
 					(reg_q0 AND symb_decoder(16#20#)) OR
 					(reg_q0 AND symb_decoder(16#ce#)) OR
 					(reg_q0 AND symb_decoder(16#ee#)) OR
 					(reg_q0 AND symb_decoder(16#46#)) OR
 					(reg_q0 AND symb_decoder(16#90#)) OR
 					(reg_q0 AND symb_decoder(16#68#)) OR
 					(reg_q0 AND symb_decoder(16#73#)) OR
 					(reg_q0 AND symb_decoder(16#c5#)) OR
 					(reg_q0 AND symb_decoder(16#6b#)) OR
 					(reg_q0 AND symb_decoder(16#d1#)) OR
 					(reg_q0 AND symb_decoder(16#85#)) OR
 					(reg_q0 AND symb_decoder(16#2b#)) OR
 					(reg_q0 AND symb_decoder(16#ef#)) OR
 					(reg_q0 AND symb_decoder(16#d5#)) OR
 					(reg_q0 AND symb_decoder(16#2a#)) OR
 					(reg_q0 AND symb_decoder(16#53#)) OR
 					(reg_q0 AND symb_decoder(16#50#)) OR
 					(reg_q0 AND symb_decoder(16#b4#)) OR
 					(reg_q0 AND symb_decoder(16#d4#)) OR
 					(reg_q0 AND symb_decoder(16#2f#)) OR
 					(reg_q0 AND symb_decoder(16#21#)) OR
 					(reg_q0 AND symb_decoder(16#d7#)) OR
 					(reg_q0 AND symb_decoder(16#a1#)) OR
 					(reg_q0 AND symb_decoder(16#69#)) OR
 					(reg_q0 AND symb_decoder(16#4d#)) OR
 					(reg_q0 AND symb_decoder(16#bd#)) OR
 					(reg_q0 AND symb_decoder(16#4a#)) OR
 					(reg_q0 AND symb_decoder(16#71#)) OR
 					(reg_q0 AND symb_decoder(16#19#)) OR
 					(reg_q0 AND symb_decoder(16#f2#)) OR
 					(reg_q0 AND symb_decoder(16#12#)) OR
 					(reg_q0 AND symb_decoder(16#83#)) OR
 					(reg_q0 AND symb_decoder(16#98#)) OR
 					(reg_q0 AND symb_decoder(16#75#)) OR
 					(reg_q0 AND symb_decoder(16#6c#)) OR
 					(reg_q0 AND symb_decoder(16#9f#)) OR
 					(reg_q0 AND symb_decoder(16#cd#)) OR
 					(reg_q0 AND symb_decoder(16#54#)) OR
 					(reg_q0 AND symb_decoder(16#fc#)) OR
 					(reg_q0 AND symb_decoder(16#c8#)) OR
 					(reg_q0 AND symb_decoder(16#57#)) OR
 					(reg_q0 AND symb_decoder(16#33#)) OR
 					(reg_q0 AND symb_decoder(16#c4#)) OR
 					(reg_q0 AND symb_decoder(16#06#)) OR
 					(reg_q0 AND symb_decoder(16#4b#)) OR
 					(reg_q0 AND symb_decoder(16#9b#)) OR
 					(reg_q0 AND symb_decoder(16#32#)) OR
 					(reg_q0 AND symb_decoder(16#5e#)) OR
 					(reg_q0 AND symb_decoder(16#94#)) OR
 					(reg_q0 AND symb_decoder(16#ab#)) OR
 					(reg_q0 AND symb_decoder(16#0a#)) OR
 					(reg_q0 AND symb_decoder(16#09#)) OR
 					(reg_q0 AND symb_decoder(16#d8#)) OR
 					(reg_q0 AND symb_decoder(16#4f#)) OR
 					(reg_q0 AND symb_decoder(16#5c#)) OR
 					(reg_q0 AND symb_decoder(16#dc#)) OR
 					(reg_q0 AND symb_decoder(16#a3#)) OR
 					(reg_q0 AND symb_decoder(16#47#)) OR
 					(reg_q0 AND symb_decoder(16#16#)) OR
 					(reg_q0 AND symb_decoder(16#f9#)) OR
 					(reg_q0 AND symb_decoder(16#4e#)) OR
 					(reg_q0 AND symb_decoder(16#55#)) OR
 					(reg_q0 AND symb_decoder(16#67#)) OR
 					(reg_q0 AND symb_decoder(16#f4#)) OR
 					(reg_q0 AND symb_decoder(16#78#)) OR
 					(reg_q0 AND symb_decoder(16#f8#)) OR
 					(reg_q0 AND symb_decoder(16#b9#)) OR
 					(reg_q0 AND symb_decoder(16#ec#)) OR
 					(reg_q0 AND symb_decoder(16#05#)) OR
 					(reg_q0 AND symb_decoder(16#a9#)) OR
 					(reg_q0 AND symb_decoder(16#fb#)) OR
 					(reg_q0 AND symb_decoder(16#1b#)) OR
 					(reg_q0 AND symb_decoder(16#3d#)) OR
 					(reg_q0 AND symb_decoder(16#d9#)) OR
 					(reg_q0 AND symb_decoder(16#1c#)) OR
 					(reg_q0 AND symb_decoder(16#cb#)) OR
 					(reg_q0 AND symb_decoder(16#58#)) OR
 					(reg_q0 AND symb_decoder(16#0e#)) OR
 					(reg_q0 AND symb_decoder(16#ad#)) OR
 					(reg_q0 AND symb_decoder(16#7e#)) OR
 					(reg_q0 AND symb_decoder(16#ac#)) OR
 					(reg_q0 AND symb_decoder(16#43#)) OR
 					(reg_q0 AND symb_decoder(16#1f#)) OR
 					(reg_q0 AND symb_decoder(16#ca#)) OR
 					(reg_q0 AND symb_decoder(16#02#)) OR
 					(reg_q0 AND symb_decoder(16#e4#)) OR
 					(reg_q0 AND symb_decoder(16#d2#)) OR
 					(reg_q0 AND symb_decoder(16#1a#)) OR
 					(reg_q0 AND symb_decoder(16#c6#)) OR
 					(reg_q0 AND symb_decoder(16#e8#)) OR
 					(reg_q0 AND symb_decoder(16#e0#)) OR
 					(reg_q0 AND symb_decoder(16#f5#)) OR
 					(reg_q0 AND symb_decoder(16#8f#)) OR
 					(reg_q0 AND symb_decoder(16#de#)) OR
 					(reg_q0 AND symb_decoder(16#e1#)) OR
 					(reg_q0 AND symb_decoder(16#f7#)) OR
 					(reg_q0 AND symb_decoder(16#a8#)) OR
 					(reg_q0 AND symb_decoder(16#5f#)) OR
 					(reg_q0 AND symb_decoder(16#3a#)) OR
 					(reg_q0 AND symb_decoder(16#49#)) OR
 					(reg_q0 AND symb_decoder(16#81#)) OR
 					(reg_q0 AND symb_decoder(16#0c#)) OR
 					(reg_q0 AND symb_decoder(16#44#)) OR
 					(reg_q0 AND symb_decoder(16#e6#)) OR
 					(reg_q0 AND symb_decoder(16#af#)) OR
 					(reg_q0 AND symb_decoder(16#11#)) OR
 					(reg_q0 AND symb_decoder(16#9d#)) OR
 					(reg_q0 AND symb_decoder(16#03#)) OR
 					(reg_q0 AND symb_decoder(16#bf#)) OR
 					(reg_q0 AND symb_decoder(16#24#)) OR
 					(reg_q0 AND symb_decoder(16#ba#)) OR
 					(reg_q0 AND symb_decoder(16#36#)) OR
 					(reg_q0 AND symb_decoder(16#6e#)) OR
 					(reg_q0 AND symb_decoder(16#35#)) OR
 					(reg_q0 AND symb_decoder(16#c9#)) OR
 					(reg_q0 AND symb_decoder(16#23#)) OR
 					(reg_q0 AND symb_decoder(16#26#)) OR
 					(reg_q0 AND symb_decoder(16#64#)) OR
 					(reg_q0 AND symb_decoder(16#59#)) OR
 					(reg_q0 AND symb_decoder(16#c7#)) OR
 					(reg_q0 AND symb_decoder(16#3c#)) OR
 					(reg_q0 AND symb_decoder(16#93#)) OR
 					(reg_q0 AND symb_decoder(16#2c#)) OR
 					(reg_q0 AND symb_decoder(16#62#)) OR
 					(reg_q0 AND symb_decoder(16#b7#)) OR
 					(reg_q0 AND symb_decoder(16#87#)) OR
 					(reg_q0 AND symb_decoder(16#7f#)) OR
 					(reg_q0 AND symb_decoder(16#cc#)) OR
 					(reg_q0 AND symb_decoder(16#52#)) OR
 					(reg_q0 AND symb_decoder(16#2e#)) OR
 					(reg_q0 AND symb_decoder(16#f3#)) OR
 					(reg_q0 AND symb_decoder(16#82#)) OR
 					(reg_q0 AND symb_decoder(16#e5#)) OR
 					(reg_q0 AND symb_decoder(16#1e#)) OR
 					(reg_q0 AND symb_decoder(16#cf#)) OR
 					(reg_q0 AND symb_decoder(16#e2#)) OR
 					(reg_q0 AND symb_decoder(16#c1#)) OR
 					(reg_q0 AND symb_decoder(16#10#)) OR
 					(reg_q0 AND symb_decoder(16#a7#)) OR
 					(reg_q0 AND symb_decoder(16#c3#)) OR
 					(reg_q0 AND symb_decoder(16#38#)) OR
 					(reg_q0 AND symb_decoder(16#f1#)) OR
 					(reg_q0 AND symb_decoder(16#29#)) OR
 					(reg_q0 AND symb_decoder(16#76#)) OR
 					(reg_q0 AND symb_decoder(16#8e#)) OR
 					(reg_q0 AND symb_decoder(16#74#)) OR
 					(reg_q0 AND symb_decoder(16#48#)) OR
 					(reg_q0 AND symb_decoder(16#80#)) OR
 					(reg_q0 AND symb_decoder(16#a6#)) OR
 					(reg_q0 AND symb_decoder(16#37#)) OR
 					(reg_q0 AND symb_decoder(16#da#)) OR
 					(reg_q0 AND symb_decoder(16#e3#)) OR
 					(reg_q0 AND symb_decoder(16#c2#)) OR
 					(reg_q0 AND symb_decoder(16#e9#)) OR
 					(reg_q0 AND symb_decoder(16#b5#)) OR
 					(reg_q0 AND symb_decoder(16#99#)) OR
 					(reg_q0 AND symb_decoder(16#31#)) OR
 					(reg_q0 AND symb_decoder(16#28#)) OR
 					(reg_q0 AND symb_decoder(16#3f#)) OR
 					(reg_q0 AND symb_decoder(16#0b#)) OR
 					(reg_q0 AND symb_decoder(16#3e#)) OR
 					(reg_q0 AND symb_decoder(16#22#)) OR
 					(reg_q0 AND symb_decoder(16#4c#)) OR
 					(reg_q0 AND symb_decoder(16#18#)) OR
 					(reg_q0 AND symb_decoder(16#8c#)) OR
 					(reg_q0 AND symb_decoder(16#60#)) OR
 					(reg_q0 AND symb_decoder(16#b3#)) OR
 					(reg_q0 AND symb_decoder(16#ed#)) OR
 					(reg_q0 AND symb_decoder(16#34#)) OR
 					(reg_q0 AND symb_decoder(16#30#)) OR
 					(reg_q0 AND symb_decoder(16#14#)) OR
 					(reg_q0 AND symb_decoder(16#bb#)) OR
 					(reg_q0 AND symb_decoder(16#b6#)) OR
 					(reg_q0 AND symb_decoder(16#aa#)) OR
 					(reg_q0 AND symb_decoder(16#96#)) OR
 					(reg_q0 AND symb_decoder(16#b2#)) OR
 					(reg_q0 AND symb_decoder(16#dd#)) OR
 					(reg_q0 AND symb_decoder(16#d0#)) OR
 					(reg_q0 AND symb_decoder(16#c0#)) OR
 					(reg_q0 AND symb_decoder(16#7d#)) OR
 					(reg_q0 AND symb_decoder(16#fd#)) OR
 					(reg_q0 AND symb_decoder(16#39#)) OR
 					(reg_q0 AND symb_decoder(16#15#)) OR
 					(reg_q0 AND symb_decoder(16#a4#)) OR
 					(reg_q0 AND symb_decoder(16#3b#)) OR
 					(reg_q0 AND symb_decoder(16#89#)) OR
 					(reg_q0 AND symb_decoder(16#ae#)) OR
 					(reg_q0 AND symb_decoder(16#2d#)) OR
 					(reg_q0 AND symb_decoder(16#13#)) OR
 					(reg_q0 AND symb_decoder(16#5d#)) OR
 					(reg_q0 AND symb_decoder(16#91#)) OR
 					(reg_q0 AND symb_decoder(16#5a#)) OR
 					(reg_q0 AND symb_decoder(16#00#)) OR
 					(reg_q0 AND symb_decoder(16#27#)) OR
 					(reg_q0 AND symb_decoder(16#25#)) OR
 					(reg_q0 AND symb_decoder(16#97#)) OR
 					(reg_q0 AND symb_decoder(16#fe#)) OR
 					(reg_q0 AND symb_decoder(16#bc#)) OR
 					(reg_q0 AND symb_decoder(16#9e#)) OR
 					(reg_q0 AND symb_decoder(16#41#)) OR
 					(reg_q0 AND symb_decoder(16#72#)) OR
 					(reg_q0 AND symb_decoder(16#b1#)) OR
 					(reg_q0 AND symb_decoder(16#8a#)) OR
 					(reg_q0 AND symb_decoder(16#88#)) OR
 					(reg_q0 AND symb_decoder(16#ff#)) OR
 					(reg_q0 AND symb_decoder(16#7c#)) OR
 					(reg_q0 AND symb_decoder(16#fa#)) OR
 					(reg_q0 AND symb_decoder(16#66#)) OR
 					(reg_q0 AND symb_decoder(16#7b#)) OR
 					(reg_q0 AND symb_decoder(16#9c#)) OR
 					(reg_q0 AND symb_decoder(16#63#)) OR
 					(reg_q0 AND symb_decoder(16#db#)) OR
 					(reg_q0 AND symb_decoder(16#6d#)) OR
 					(reg_q0 AND symb_decoder(16#eb#)) OR
 					(reg_q0 AND symb_decoder(16#04#)) OR
 					(reg_q0 AND symb_decoder(16#0f#)) OR
 					(reg_q0 AND symb_decoder(16#07#)) OR
 					(reg_q0 AND symb_decoder(16#e7#)) OR
 					(reg_q0 AND symb_decoder(16#17#)) OR
 					(reg_q0 AND symb_decoder(16#95#)) OR
 					(reg_q0 AND symb_decoder(16#0d#)) OR
 					(reg_q0 AND symb_decoder(16#70#)) OR
 					(reg_q0 AND symb_decoder(16#61#)) OR
 					(reg_q0 AND symb_decoder(16#7a#)) OR
 					(reg_q0 AND symb_decoder(16#ea#)) OR
 					(reg_q0 AND symb_decoder(16#a0#)) OR
 					(reg_q0 AND symb_decoder(16#5b#)) OR
 					(reg_q0 AND symb_decoder(16#51#)) OR
 					(reg_q0 AND symb_decoder(16#df#)) OR
 					(reg_q0 AND symb_decoder(16#1d#)) OR
 					(reg_q0 AND symb_decoder(16#45#)) OR
 					(reg_q0 AND symb_decoder(16#8d#)) OR
 					(reg_q0 AND symb_decoder(16#77#)) OR
 					(reg_q0 AND symb_decoder(16#6a#)) OR
 					(reg_q0 AND symb_decoder(16#f6#)) OR
 					(reg_q0 AND symb_decoder(16#f0#)) OR
 					(reg_q0 AND symb_decoder(16#d6#)) OR
 					(reg_q0 AND symb_decoder(16#86#)) OR
 					(reg_q0 AND symb_decoder(16#b8#)) OR
 					(reg_q0 AND symb_decoder(16#92#)) OR
 					(reg_q0 AND symb_decoder(16#56#)) OR
 					(reg_q0 AND symb_decoder(16#84#)) OR
 					(reg_q0 AND symb_decoder(16#42#)) OR
 					(reg_q0 AND symb_decoder(16#b0#)) OR
 					(reg_q0 AND symb_decoder(16#65#)) OR
 					(reg_q0 AND symb_decoder(16#be#)) OR
 					(reg_q0 AND symb_decoder(16#40#));
reg_q0_init <= '0' ;
	p_reg_q0: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q0 <= reg_q0_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q0 <= reg_q0_init;
        else
          reg_q0 <= reg_q0_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q850_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q850 AND symb_decoder(16#a2#)) OR
 					(reg_q850 AND symb_decoder(16#b3#)) OR
 					(reg_q850 AND symb_decoder(16#08#)) OR
 					(reg_q850 AND symb_decoder(16#36#)) OR
 					(reg_q850 AND symb_decoder(16#fb#)) OR
 					(reg_q850 AND symb_decoder(16#a8#)) OR
 					(reg_q850 AND symb_decoder(16#6a#)) OR
 					(reg_q850 AND symb_decoder(16#92#)) OR
 					(reg_q850 AND symb_decoder(16#c7#)) OR
 					(reg_q850 AND symb_decoder(16#32#)) OR
 					(reg_q850 AND symb_decoder(16#70#)) OR
 					(reg_q850 AND symb_decoder(16#cc#)) OR
 					(reg_q850 AND symb_decoder(16#87#)) OR
 					(reg_q850 AND symb_decoder(16#7f#)) OR
 					(reg_q850 AND symb_decoder(16#f5#)) OR
 					(reg_q850 AND symb_decoder(16#3d#)) OR
 					(reg_q850 AND symb_decoder(16#8a#)) OR
 					(reg_q850 AND symb_decoder(16#da#)) OR
 					(reg_q850 AND symb_decoder(16#df#)) OR
 					(reg_q850 AND symb_decoder(16#62#)) OR
 					(reg_q850 AND symb_decoder(16#a5#)) OR
 					(reg_q850 AND symb_decoder(16#9a#)) OR
 					(reg_q850 AND symb_decoder(16#be#)) OR
 					(reg_q850 AND symb_decoder(16#48#)) OR
 					(reg_q850 AND symb_decoder(16#05#)) OR
 					(reg_q850 AND symb_decoder(16#5b#)) OR
 					(reg_q850 AND symb_decoder(16#aa#)) OR
 					(reg_q850 AND symb_decoder(16#f9#)) OR
 					(reg_q850 AND symb_decoder(16#31#)) OR
 					(reg_q850 AND symb_decoder(16#20#)) OR
 					(reg_q850 AND symb_decoder(16#ef#)) OR
 					(reg_q850 AND symb_decoder(16#cb#)) OR
 					(reg_q850 AND symb_decoder(16#9e#)) OR
 					(reg_q850 AND symb_decoder(16#d5#)) OR
 					(reg_q850 AND symb_decoder(16#f3#)) OR
 					(reg_q850 AND symb_decoder(16#d4#)) OR
 					(reg_q850 AND symb_decoder(16#24#)) OR
 					(reg_q850 AND symb_decoder(16#f8#)) OR
 					(reg_q850 AND symb_decoder(16#15#)) OR
 					(reg_q850 AND symb_decoder(16#4d#)) OR
 					(reg_q850 AND symb_decoder(16#8c#)) OR
 					(reg_q850 AND symb_decoder(16#9c#)) OR
 					(reg_q850 AND symb_decoder(16#ad#)) OR
 					(reg_q850 AND symb_decoder(16#c4#)) OR
 					(reg_q850 AND symb_decoder(16#e0#)) OR
 					(reg_q850 AND symb_decoder(16#b1#)) OR
 					(reg_q850 AND symb_decoder(16#17#)) OR
 					(reg_q850 AND symb_decoder(16#39#)) OR
 					(reg_q850 AND symb_decoder(16#23#)) OR
 					(reg_q850 AND symb_decoder(16#3e#)) OR
 					(reg_q850 AND symb_decoder(16#e5#)) OR
 					(reg_q850 AND symb_decoder(16#c6#)) OR
 					(reg_q850 AND symb_decoder(16#a0#)) OR
 					(reg_q850 AND symb_decoder(16#ae#)) OR
 					(reg_q850 AND symb_decoder(16#47#)) OR
 					(reg_q850 AND symb_decoder(16#fe#)) OR
 					(reg_q850 AND symb_decoder(16#33#)) OR
 					(reg_q850 AND symb_decoder(16#29#)) OR
 					(reg_q850 AND symb_decoder(16#ec#)) OR
 					(reg_q850 AND symb_decoder(16#79#)) OR
 					(reg_q850 AND symb_decoder(16#72#)) OR
 					(reg_q850 AND symb_decoder(16#3b#)) OR
 					(reg_q850 AND symb_decoder(16#b8#)) OR
 					(reg_q850 AND symb_decoder(16#f6#)) OR
 					(reg_q850 AND symb_decoder(16#4a#)) OR
 					(reg_q850 AND symb_decoder(16#3c#)) OR
 					(reg_q850 AND symb_decoder(16#56#)) OR
 					(reg_q850 AND symb_decoder(16#07#)) OR
 					(reg_q850 AND symb_decoder(16#d2#)) OR
 					(reg_q850 AND symb_decoder(16#53#)) OR
 					(reg_q850 AND symb_decoder(16#b2#)) OR
 					(reg_q850 AND symb_decoder(16#80#)) OR
 					(reg_q850 AND symb_decoder(16#95#)) OR
 					(reg_q850 AND symb_decoder(16#5e#)) OR
 					(reg_q850 AND symb_decoder(16#ee#)) OR
 					(reg_q850 AND symb_decoder(16#c5#)) OR
 					(reg_q850 AND symb_decoder(16#28#)) OR
 					(reg_q850 AND symb_decoder(16#f0#)) OR
 					(reg_q850 AND symb_decoder(16#a3#)) OR
 					(reg_q850 AND symb_decoder(16#26#)) OR
 					(reg_q850 AND symb_decoder(16#64#)) OR
 					(reg_q850 AND symb_decoder(16#37#)) OR
 					(reg_q850 AND symb_decoder(16#c2#)) OR
 					(reg_q850 AND symb_decoder(16#2f#)) OR
 					(reg_q850 AND symb_decoder(16#94#)) OR
 					(reg_q850 AND symb_decoder(16#7e#)) OR
 					(reg_q850 AND symb_decoder(16#eb#)) OR
 					(reg_q850 AND symb_decoder(16#67#)) OR
 					(reg_q850 AND symb_decoder(16#42#)) OR
 					(reg_q850 AND symb_decoder(16#bb#)) OR
 					(reg_q850 AND symb_decoder(16#ac#)) OR
 					(reg_q850 AND symb_decoder(16#de#)) OR
 					(reg_q850 AND symb_decoder(16#6e#)) OR
 					(reg_q850 AND symb_decoder(16#61#)) OR
 					(reg_q850 AND symb_decoder(16#75#)) OR
 					(reg_q850 AND symb_decoder(16#74#)) OR
 					(reg_q850 AND symb_decoder(16#9d#)) OR
 					(reg_q850 AND symb_decoder(16#5f#)) OR
 					(reg_q850 AND symb_decoder(16#93#)) OR
 					(reg_q850 AND symb_decoder(16#e2#)) OR
 					(reg_q850 AND symb_decoder(16#d1#)) OR
 					(reg_q850 AND symb_decoder(16#b6#)) OR
 					(reg_q850 AND symb_decoder(16#fd#)) OR
 					(reg_q850 AND symb_decoder(16#85#)) OR
 					(reg_q850 AND symb_decoder(16#18#)) OR
 					(reg_q850 AND symb_decoder(16#b5#)) OR
 					(reg_q850 AND symb_decoder(16#bc#)) OR
 					(reg_q850 AND symb_decoder(16#e7#)) OR
 					(reg_q850 AND symb_decoder(16#82#)) OR
 					(reg_q850 AND symb_decoder(16#4e#)) OR
 					(reg_q850 AND symb_decoder(16#e6#)) OR
 					(reg_q850 AND symb_decoder(16#cf#)) OR
 					(reg_q850 AND symb_decoder(16#25#)) OR
 					(reg_q850 AND symb_decoder(16#78#)) OR
 					(reg_q850 AND symb_decoder(16#0f#)) OR
 					(reg_q850 AND symb_decoder(16#58#)) OR
 					(reg_q850 AND symb_decoder(16#e8#)) OR
 					(reg_q850 AND symb_decoder(16#69#)) OR
 					(reg_q850 AND symb_decoder(16#00#)) OR
 					(reg_q850 AND symb_decoder(16#98#)) OR
 					(reg_q850 AND symb_decoder(16#c8#)) OR
 					(reg_q850 AND symb_decoder(16#8f#)) OR
 					(reg_q850 AND symb_decoder(16#44#)) OR
 					(reg_q850 AND symb_decoder(16#55#)) OR
 					(reg_q850 AND symb_decoder(16#a1#)) OR
 					(reg_q850 AND symb_decoder(16#66#)) OR
 					(reg_q850 AND symb_decoder(16#40#)) OR
 					(reg_q850 AND symb_decoder(16#65#)) OR
 					(reg_q850 AND symb_decoder(16#c1#)) OR
 					(reg_q850 AND symb_decoder(16#3a#)) OR
 					(reg_q850 AND symb_decoder(16#2e#)) OR
 					(reg_q850 AND symb_decoder(16#60#)) OR
 					(reg_q850 AND symb_decoder(16#01#)) OR
 					(reg_q850 AND symb_decoder(16#89#)) OR
 					(reg_q850 AND symb_decoder(16#35#)) OR
 					(reg_q850 AND symb_decoder(16#7a#)) OR
 					(reg_q850 AND symb_decoder(16#52#)) OR
 					(reg_q850 AND symb_decoder(16#34#)) OR
 					(reg_q850 AND symb_decoder(16#2c#)) OR
 					(reg_q850 AND symb_decoder(16#0e#)) OR
 					(reg_q850 AND symb_decoder(16#38#)) OR
 					(reg_q850 AND symb_decoder(16#db#)) OR
 					(reg_q850 AND symb_decoder(16#7b#)) OR
 					(reg_q850 AND symb_decoder(16#b4#)) OR
 					(reg_q850 AND symb_decoder(16#06#)) OR
 					(reg_q850 AND symb_decoder(16#bd#)) OR
 					(reg_q850 AND symb_decoder(16#10#)) OR
 					(reg_q850 AND symb_decoder(16#9b#)) OR
 					(reg_q850 AND symb_decoder(16#7c#)) OR
 					(reg_q850 AND symb_decoder(16#7d#)) OR
 					(reg_q850 AND symb_decoder(16#ca#)) OR
 					(reg_q850 AND symb_decoder(16#84#)) OR
 					(reg_q850 AND symb_decoder(16#6d#)) OR
 					(reg_q850 AND symb_decoder(16#6f#)) OR
 					(reg_q850 AND symb_decoder(16#0a#)) OR
 					(reg_q850 AND symb_decoder(16#57#)) OR
 					(reg_q850 AND symb_decoder(16#b7#)) OR
 					(reg_q850 AND symb_decoder(16#1f#)) OR
 					(reg_q850 AND symb_decoder(16#1a#)) OR
 					(reg_q850 AND symb_decoder(16#86#)) OR
 					(reg_q850 AND symb_decoder(16#ab#)) OR
 					(reg_q850 AND symb_decoder(16#96#)) OR
 					(reg_q850 AND symb_decoder(16#77#)) OR
 					(reg_q850 AND symb_decoder(16#27#)) OR
 					(reg_q850 AND symb_decoder(16#2d#)) OR
 					(reg_q850 AND symb_decoder(16#6b#)) OR
 					(reg_q850 AND symb_decoder(16#ea#)) OR
 					(reg_q850 AND symb_decoder(16#4f#)) OR
 					(reg_q850 AND symb_decoder(16#a4#)) OR
 					(reg_q850 AND symb_decoder(16#e9#)) OR
 					(reg_q850 AND symb_decoder(16#68#)) OR
 					(reg_q850 AND symb_decoder(16#22#)) OR
 					(reg_q850 AND symb_decoder(16#41#)) OR
 					(reg_q850 AND symb_decoder(16#ce#)) OR
 					(reg_q850 AND symb_decoder(16#a7#)) OR
 					(reg_q850 AND symb_decoder(16#a6#)) OR
 					(reg_q850 AND symb_decoder(16#0d#)) OR
 					(reg_q850 AND symb_decoder(16#73#)) OR
 					(reg_q850 AND symb_decoder(16#59#)) OR
 					(reg_q850 AND symb_decoder(16#1c#)) OR
 					(reg_q850 AND symb_decoder(16#e1#)) OR
 					(reg_q850 AND symb_decoder(16#09#)) OR
 					(reg_q850 AND symb_decoder(16#d8#)) OR
 					(reg_q850 AND symb_decoder(16#cd#)) OR
 					(reg_q850 AND symb_decoder(16#54#)) OR
 					(reg_q850 AND symb_decoder(16#d0#)) OR
 					(reg_q850 AND symb_decoder(16#b0#)) OR
 					(reg_q850 AND symb_decoder(16#3f#)) OR
 					(reg_q850 AND symb_decoder(16#45#)) OR
 					(reg_q850 AND symb_decoder(16#1e#)) OR
 					(reg_q850 AND symb_decoder(16#1d#)) OR
 					(reg_q850 AND symb_decoder(16#a9#)) OR
 					(reg_q850 AND symb_decoder(16#e3#)) OR
 					(reg_q850 AND symb_decoder(16#97#)) OR
 					(reg_q850 AND symb_decoder(16#f7#)) OR
 					(reg_q850 AND symb_decoder(16#c0#)) OR
 					(reg_q850 AND symb_decoder(16#e4#)) OR
 					(reg_q850 AND symb_decoder(16#f1#)) OR
 					(reg_q850 AND symb_decoder(16#51#)) OR
 					(reg_q850 AND symb_decoder(16#ba#)) OR
 					(reg_q850 AND symb_decoder(16#2a#)) OR
 					(reg_q850 AND symb_decoder(16#88#)) OR
 					(reg_q850 AND symb_decoder(16#83#)) OR
 					(reg_q850 AND symb_decoder(16#12#)) OR
 					(reg_q850 AND symb_decoder(16#6c#)) OR
 					(reg_q850 AND symb_decoder(16#4b#)) OR
 					(reg_q850 AND symb_decoder(16#81#)) OR
 					(reg_q850 AND symb_decoder(16#11#)) OR
 					(reg_q850 AND symb_decoder(16#d3#)) OR
 					(reg_q850 AND symb_decoder(16#b9#)) OR
 					(reg_q850 AND symb_decoder(16#dd#)) OR
 					(reg_q850 AND symb_decoder(16#dc#)) OR
 					(reg_q850 AND symb_decoder(16#76#)) OR
 					(reg_q850 AND symb_decoder(16#21#)) OR
 					(reg_q850 AND symb_decoder(16#d9#)) OR
 					(reg_q850 AND symb_decoder(16#8b#)) OR
 					(reg_q850 AND symb_decoder(16#c3#)) OR
 					(reg_q850 AND symb_decoder(16#ff#)) OR
 					(reg_q850 AND symb_decoder(16#13#)) OR
 					(reg_q850 AND symb_decoder(16#f2#)) OR
 					(reg_q850 AND symb_decoder(16#02#)) OR
 					(reg_q850 AND symb_decoder(16#91#)) OR
 					(reg_q850 AND symb_decoder(16#43#)) OR
 					(reg_q850 AND symb_decoder(16#c9#)) OR
 					(reg_q850 AND symb_decoder(16#16#)) OR
 					(reg_q850 AND symb_decoder(16#63#)) OR
 					(reg_q850 AND symb_decoder(16#50#)) OR
 					(reg_q850 AND symb_decoder(16#5d#)) OR
 					(reg_q850 AND symb_decoder(16#1b#)) OR
 					(reg_q850 AND symb_decoder(16#fc#)) OR
 					(reg_q850 AND symb_decoder(16#71#)) OR
 					(reg_q850 AND symb_decoder(16#90#)) OR
 					(reg_q850 AND symb_decoder(16#8e#)) OR
 					(reg_q850 AND symb_decoder(16#0c#)) OR
 					(reg_q850 AND symb_decoder(16#5c#)) OR
 					(reg_q850 AND symb_decoder(16#bf#)) OR
 					(reg_q850 AND symb_decoder(16#2b#)) OR
 					(reg_q850 AND symb_decoder(16#04#)) OR
 					(reg_q850 AND symb_decoder(16#f4#)) OR
 					(reg_q850 AND symb_decoder(16#14#)) OR
 					(reg_q850 AND symb_decoder(16#30#)) OR
 					(reg_q850 AND symb_decoder(16#0b#)) OR
 					(reg_q850 AND symb_decoder(16#5a#)) OR
 					(reg_q850 AND symb_decoder(16#af#)) OR
 					(reg_q850 AND symb_decoder(16#ed#)) OR
 					(reg_q850 AND symb_decoder(16#19#)) OR
 					(reg_q850 AND symb_decoder(16#4c#)) OR
 					(reg_q850 AND symb_decoder(16#99#)) OR
 					(reg_q850 AND symb_decoder(16#46#)) OR
 					(reg_q850 AND symb_decoder(16#8d#)) OR
 					(reg_q850 AND symb_decoder(16#fa#)) OR
 					(reg_q850 AND symb_decoder(16#d7#)) OR
 					(reg_q850 AND symb_decoder(16#d6#)) OR
 					(reg_q850 AND symb_decoder(16#03#)) OR
 					(reg_q850 AND symb_decoder(16#9f#)) OR
 					(reg_q850 AND symb_decoder(16#49#));
reg_q850_init <= '0' ;
	p_reg_q850: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q850 <= reg_q850_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q850 <= reg_q850_init;
        else
          reg_q850 <= reg_q850_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph10

reg_q2615_in <= (reg_q2579 AND symb_decoder(16#79#)) OR
 					(reg_q2579 AND symb_decoder(16#62#)) OR
 					(reg_q2579 AND symb_decoder(16#7d#)) OR
 					(reg_q2579 AND symb_decoder(16#3a#)) OR
 					(reg_q2579 AND symb_decoder(16#b0#)) OR
 					(reg_q2579 AND symb_decoder(16#ca#)) OR
 					(reg_q2579 AND symb_decoder(16#ec#)) OR
 					(reg_q2579 AND symb_decoder(16#55#)) OR
 					(reg_q2579 AND symb_decoder(16#77#)) OR
 					(reg_q2579 AND symb_decoder(16#66#)) OR
 					(reg_q2579 AND symb_decoder(16#bb#)) OR
 					(reg_q2579 AND symb_decoder(16#4c#)) OR
 					(reg_q2579 AND symb_decoder(16#c6#)) OR
 					(reg_q2579 AND symb_decoder(16#ac#)) OR
 					(reg_q2579 AND symb_decoder(16#c2#)) OR
 					(reg_q2579 AND symb_decoder(16#27#)) OR
 					(reg_q2579 AND symb_decoder(16#a9#)) OR
 					(reg_q2579 AND symb_decoder(16#5c#)) OR
 					(reg_q2579 AND symb_decoder(16#d1#)) OR
 					(reg_q2579 AND symb_decoder(16#da#)) OR
 					(reg_q2579 AND symb_decoder(16#8a#)) OR
 					(reg_q2579 AND symb_decoder(16#5b#)) OR
 					(reg_q2579 AND symb_decoder(16#c8#)) OR
 					(reg_q2579 AND symb_decoder(16#1a#)) OR
 					(reg_q2579 AND symb_decoder(16#e0#)) OR
 					(reg_q2579 AND symb_decoder(16#09#)) OR
 					(reg_q2579 AND symb_decoder(16#06#)) OR
 					(reg_q2579 AND symb_decoder(16#64#)) OR
 					(reg_q2579 AND symb_decoder(16#30#)) OR
 					(reg_q2579 AND symb_decoder(16#8e#)) OR
 					(reg_q2579 AND symb_decoder(16#10#)) OR
 					(reg_q2579 AND symb_decoder(16#cb#)) OR
 					(reg_q2579 AND symb_decoder(16#a2#)) OR
 					(reg_q2579 AND symb_decoder(16#57#)) OR
 					(reg_q2579 AND symb_decoder(16#c5#)) OR
 					(reg_q2579 AND symb_decoder(16#28#)) OR
 					(reg_q2579 AND symb_decoder(16#36#)) OR
 					(reg_q2579 AND symb_decoder(16#61#)) OR
 					(reg_q2579 AND symb_decoder(16#c0#)) OR
 					(reg_q2579 AND symb_decoder(16#b9#)) OR
 					(reg_q2579 AND symb_decoder(16#7a#)) OR
 					(reg_q2579 AND symb_decoder(16#19#)) OR
 					(reg_q2579 AND symb_decoder(16#ce#)) OR
 					(reg_q2579 AND symb_decoder(16#04#)) OR
 					(reg_q2579 AND symb_decoder(16#41#)) OR
 					(reg_q2579 AND symb_decoder(16#42#)) OR
 					(reg_q2579 AND symb_decoder(16#ab#)) OR
 					(reg_q2579 AND symb_decoder(16#13#)) OR
 					(reg_q2579 AND symb_decoder(16#db#)) OR
 					(reg_q2579 AND symb_decoder(16#48#)) OR
 					(reg_q2579 AND symb_decoder(16#aa#)) OR
 					(reg_q2579 AND symb_decoder(16#17#)) OR
 					(reg_q2579 AND symb_decoder(16#dd#)) OR
 					(reg_q2579 AND symb_decoder(16#03#)) OR
 					(reg_q2579 AND symb_decoder(16#2c#)) OR
 					(reg_q2579 AND symb_decoder(16#6d#)) OR
 					(reg_q2579 AND symb_decoder(16#ef#)) OR
 					(reg_q2579 AND symb_decoder(16#e1#)) OR
 					(reg_q2579 AND symb_decoder(16#9c#)) OR
 					(reg_q2579 AND symb_decoder(16#8c#)) OR
 					(reg_q2579 AND symb_decoder(16#3f#)) OR
 					(reg_q2579 AND symb_decoder(16#d2#)) OR
 					(reg_q2579 AND symb_decoder(16#33#)) OR
 					(reg_q2579 AND symb_decoder(16#bd#)) OR
 					(reg_q2579 AND symb_decoder(16#58#)) OR
 					(reg_q2579 AND symb_decoder(16#ad#)) OR
 					(reg_q2579 AND symb_decoder(16#3c#)) OR
 					(reg_q2579 AND symb_decoder(16#81#)) OR
 					(reg_q2579 AND symb_decoder(16#b1#)) OR
 					(reg_q2579 AND symb_decoder(16#fd#)) OR
 					(reg_q2579 AND symb_decoder(16#fe#)) OR
 					(reg_q2579 AND symb_decoder(16#08#)) OR
 					(reg_q2579 AND symb_decoder(16#98#)) OR
 					(reg_q2579 AND symb_decoder(16#fa#)) OR
 					(reg_q2579 AND symb_decoder(16#e3#)) OR
 					(reg_q2579 AND symb_decoder(16#54#)) OR
 					(reg_q2579 AND symb_decoder(16#cd#)) OR
 					(reg_q2579 AND symb_decoder(16#e4#)) OR
 					(reg_q2579 AND symb_decoder(16#f4#)) OR
 					(reg_q2579 AND symb_decoder(16#72#)) OR
 					(reg_q2579 AND symb_decoder(16#2f#)) OR
 					(reg_q2579 AND symb_decoder(16#6a#)) OR
 					(reg_q2579 AND symb_decoder(16#a8#)) OR
 					(reg_q2579 AND symb_decoder(16#e8#)) OR
 					(reg_q2579 AND symb_decoder(16#52#)) OR
 					(reg_q2579 AND symb_decoder(16#ba#)) OR
 					(reg_q2579 AND symb_decoder(16#0e#)) OR
 					(reg_q2579 AND symb_decoder(16#92#)) OR
 					(reg_q2579 AND symb_decoder(16#47#)) OR
 					(reg_q2579 AND symb_decoder(16#7b#)) OR
 					(reg_q2579 AND symb_decoder(16#b5#)) OR
 					(reg_q2579 AND symb_decoder(16#e7#)) OR
 					(reg_q2579 AND symb_decoder(16#6b#)) OR
 					(reg_q2579 AND symb_decoder(16#7e#)) OR
 					(reg_q2579 AND symb_decoder(16#9a#)) OR
 					(reg_q2579 AND symb_decoder(16#26#)) OR
 					(reg_q2579 AND symb_decoder(16#3d#)) OR
 					(reg_q2579 AND symb_decoder(16#69#)) OR
 					(reg_q2579 AND symb_decoder(16#83#)) OR
 					(reg_q2579 AND symb_decoder(16#2e#)) OR
 					(reg_q2579 AND symb_decoder(16#2d#)) OR
 					(reg_q2579 AND symb_decoder(16#7c#)) OR
 					(reg_q2579 AND symb_decoder(16#d3#)) OR
 					(reg_q2579 AND symb_decoder(16#5d#)) OR
 					(reg_q2579 AND symb_decoder(16#b7#)) OR
 					(reg_q2579 AND symb_decoder(16#94#)) OR
 					(reg_q2579 AND symb_decoder(16#d5#)) OR
 					(reg_q2579 AND symb_decoder(16#a3#)) OR
 					(reg_q2579 AND symb_decoder(16#20#)) OR
 					(reg_q2579 AND symb_decoder(16#9e#)) OR
 					(reg_q2579 AND symb_decoder(16#39#)) OR
 					(reg_q2579 AND symb_decoder(16#31#)) OR
 					(reg_q2579 AND symb_decoder(16#35#)) OR
 					(reg_q2579 AND symb_decoder(16#1f#)) OR
 					(reg_q2579 AND symb_decoder(16#85#)) OR
 					(reg_q2579 AND symb_decoder(16#73#)) OR
 					(reg_q2579 AND symb_decoder(16#a6#)) OR
 					(reg_q2579 AND symb_decoder(16#d4#)) OR
 					(reg_q2579 AND symb_decoder(16#82#)) OR
 					(reg_q2579 AND symb_decoder(16#de#)) OR
 					(reg_q2579 AND symb_decoder(16#b3#)) OR
 					(reg_q2579 AND symb_decoder(16#f2#)) OR
 					(reg_q2579 AND symb_decoder(16#8b#)) OR
 					(reg_q2579 AND symb_decoder(16#d9#)) OR
 					(reg_q2579 AND symb_decoder(16#0c#)) OR
 					(reg_q2579 AND symb_decoder(16#dc#)) OR
 					(reg_q2579 AND symb_decoder(16#45#)) OR
 					(reg_q2579 AND symb_decoder(16#e5#)) OR
 					(reg_q2579 AND symb_decoder(16#8f#)) OR
 					(reg_q2579 AND symb_decoder(16#e2#)) OR
 					(reg_q2579 AND symb_decoder(16#6e#)) OR
 					(reg_q2579 AND symb_decoder(16#70#)) OR
 					(reg_q2579 AND symb_decoder(16#f0#)) OR
 					(reg_q2579 AND symb_decoder(16#f7#)) OR
 					(reg_q2579 AND symb_decoder(16#ed#)) OR
 					(reg_q2579 AND symb_decoder(16#3e#)) OR
 					(reg_q2579 AND symb_decoder(16#f3#)) OR
 					(reg_q2579 AND symb_decoder(16#6c#)) OR
 					(reg_q2579 AND symb_decoder(16#86#)) OR
 					(reg_q2579 AND symb_decoder(16#38#)) OR
 					(reg_q2579 AND symb_decoder(16#29#)) OR
 					(reg_q2579 AND symb_decoder(16#c7#)) OR
 					(reg_q2579 AND symb_decoder(16#1d#)) OR
 					(reg_q2579 AND symb_decoder(16#75#)) OR
 					(reg_q2579 AND symb_decoder(16#97#)) OR
 					(reg_q2579 AND symb_decoder(16#78#)) OR
 					(reg_q2579 AND symb_decoder(16#9b#)) OR
 					(reg_q2579 AND symb_decoder(16#d0#)) OR
 					(reg_q2579 AND symb_decoder(16#22#)) OR
 					(reg_q2579 AND symb_decoder(16#63#)) OR
 					(reg_q2579 AND symb_decoder(16#b6#)) OR
 					(reg_q2579 AND symb_decoder(16#01#)) OR
 					(reg_q2579 AND symb_decoder(16#91#)) OR
 					(reg_q2579 AND symb_decoder(16#49#)) OR
 					(reg_q2579 AND symb_decoder(16#bc#)) OR
 					(reg_q2579 AND symb_decoder(16#43#)) OR
 					(reg_q2579 AND symb_decoder(16#76#)) OR
 					(reg_q2579 AND symb_decoder(16#37#)) OR
 					(reg_q2579 AND symb_decoder(16#6f#)) OR
 					(reg_q2579 AND symb_decoder(16#51#)) OR
 					(reg_q2579 AND symb_decoder(16#0b#)) OR
 					(reg_q2579 AND symb_decoder(16#c4#)) OR
 					(reg_q2579 AND symb_decoder(16#56#)) OR
 					(reg_q2579 AND symb_decoder(16#df#)) OR
 					(reg_q2579 AND symb_decoder(16#65#)) OR
 					(reg_q2579 AND symb_decoder(16#40#)) OR
 					(reg_q2579 AND symb_decoder(16#5f#)) OR
 					(reg_q2579 AND symb_decoder(16#b2#)) OR
 					(reg_q2579 AND symb_decoder(16#89#)) OR
 					(reg_q2579 AND symb_decoder(16#ff#)) OR
 					(reg_q2579 AND symb_decoder(16#f6#)) OR
 					(reg_q2579 AND symb_decoder(16#c9#)) OR
 					(reg_q2579 AND symb_decoder(16#3b#)) OR
 					(reg_q2579 AND symb_decoder(16#fb#)) OR
 					(reg_q2579 AND symb_decoder(16#f1#)) OR
 					(reg_q2579 AND symb_decoder(16#18#)) OR
 					(reg_q2579 AND symb_decoder(16#f8#)) OR
 					(reg_q2579 AND symb_decoder(16#ae#)) OR
 					(reg_q2579 AND symb_decoder(16#f5#)) OR
 					(reg_q2579 AND symb_decoder(16#4e#)) OR
 					(reg_q2579 AND symb_decoder(16#1b#)) OR
 					(reg_q2579 AND symb_decoder(16#74#)) OR
 					(reg_q2579 AND symb_decoder(16#d7#)) OR
 					(reg_q2579 AND symb_decoder(16#a5#)) OR
 					(reg_q2579 AND symb_decoder(16#44#)) OR
 					(reg_q2579 AND symb_decoder(16#5a#)) OR
 					(reg_q2579 AND symb_decoder(16#1c#)) OR
 					(reg_q2579 AND symb_decoder(16#99#)) OR
 					(reg_q2579 AND symb_decoder(16#68#)) OR
 					(reg_q2579 AND symb_decoder(16#05#)) OR
 					(reg_q2579 AND symb_decoder(16#c3#)) OR
 					(reg_q2579 AND symb_decoder(16#e6#)) OR
 					(reg_q2579 AND symb_decoder(16#af#)) OR
 					(reg_q2579 AND symb_decoder(16#4a#)) OR
 					(reg_q2579 AND symb_decoder(16#15#)) OR
 					(reg_q2579 AND symb_decoder(16#1e#)) OR
 					(reg_q2579 AND symb_decoder(16#93#)) OR
 					(reg_q2579 AND symb_decoder(16#d6#)) OR
 					(reg_q2579 AND symb_decoder(16#4f#)) OR
 					(reg_q2579 AND symb_decoder(16#12#)) OR
 					(reg_q2579 AND symb_decoder(16#53#)) OR
 					(reg_q2579 AND symb_decoder(16#02#)) OR
 					(reg_q2579 AND symb_decoder(16#21#)) OR
 					(reg_q2579 AND symb_decoder(16#16#)) OR
 					(reg_q2579 AND symb_decoder(16#cc#)) OR
 					(reg_q2579 AND symb_decoder(16#eb#)) OR
 					(reg_q2579 AND symb_decoder(16#b8#)) OR
 					(reg_q2579 AND symb_decoder(16#7f#)) OR
 					(reg_q2579 AND symb_decoder(16#8d#)) OR
 					(reg_q2579 AND symb_decoder(16#a1#)) OR
 					(reg_q2579 AND symb_decoder(16#f9#)) OR
 					(reg_q2579 AND symb_decoder(16#46#)) OR
 					(reg_q2579 AND symb_decoder(16#14#)) OR
 					(reg_q2579 AND symb_decoder(16#87#)) OR
 					(reg_q2579 AND symb_decoder(16#0f#)) OR
 					(reg_q2579 AND symb_decoder(16#67#)) OR
 					(reg_q2579 AND symb_decoder(16#71#)) OR
 					(reg_q2579 AND symb_decoder(16#4b#)) OR
 					(reg_q2579 AND symb_decoder(16#e9#)) OR
 					(reg_q2579 AND symb_decoder(16#fc#)) OR
 					(reg_q2579 AND symb_decoder(16#a0#)) OR
 					(reg_q2579 AND symb_decoder(16#a7#)) OR
 					(reg_q2579 AND symb_decoder(16#4d#)) OR
 					(reg_q2579 AND symb_decoder(16#cf#)) OR
 					(reg_q2579 AND symb_decoder(16#84#)) OR
 					(reg_q2579 AND symb_decoder(16#07#)) OR
 					(reg_q2579 AND symb_decoder(16#ea#)) OR
 					(reg_q2579 AND symb_decoder(16#d8#)) OR
 					(reg_q2579 AND symb_decoder(16#95#)) OR
 					(reg_q2579 AND symb_decoder(16#00#)) OR
 					(reg_q2579 AND symb_decoder(16#80#)) OR
 					(reg_q2579 AND symb_decoder(16#60#)) OR
 					(reg_q2579 AND symb_decoder(16#11#)) OR
 					(reg_q2579 AND symb_decoder(16#c1#)) OR
 					(reg_q2579 AND symb_decoder(16#34#)) OR
 					(reg_q2579 AND symb_decoder(16#59#)) OR
 					(reg_q2579 AND symb_decoder(16#24#)) OR
 					(reg_q2579 AND symb_decoder(16#23#)) OR
 					(reg_q2579 AND symb_decoder(16#a4#)) OR
 					(reg_q2579 AND symb_decoder(16#25#)) OR
 					(reg_q2579 AND symb_decoder(16#ee#)) OR
 					(reg_q2579 AND symb_decoder(16#50#)) OR
 					(reg_q2579 AND symb_decoder(16#2a#)) OR
 					(reg_q2579 AND symb_decoder(16#90#)) OR
 					(reg_q2579 AND symb_decoder(16#be#)) OR
 					(reg_q2579 AND symb_decoder(16#9f#)) OR
 					(reg_q2579 AND symb_decoder(16#5e#)) OR
 					(reg_q2579 AND symb_decoder(16#b4#)) OR
 					(reg_q2579 AND symb_decoder(16#bf#)) OR
 					(reg_q2579 AND symb_decoder(16#96#)) OR
 					(reg_q2579 AND symb_decoder(16#88#)) OR
 					(reg_q2579 AND symb_decoder(16#2b#)) OR
 					(reg_q2579 AND symb_decoder(16#32#)) OR
 					(reg_q2579 AND symb_decoder(16#9d#)) OR
 					(reg_q2615 AND symb_decoder(16#a9#)) OR
 					(reg_q2615 AND symb_decoder(16#78#)) OR
 					(reg_q2615 AND symb_decoder(16#b7#)) OR
 					(reg_q2615 AND symb_decoder(16#e1#)) OR
 					(reg_q2615 AND symb_decoder(16#4f#)) OR
 					(reg_q2615 AND symb_decoder(16#34#)) OR
 					(reg_q2615 AND symb_decoder(16#d9#)) OR
 					(reg_q2615 AND symb_decoder(16#b5#)) OR
 					(reg_q2615 AND symb_decoder(16#3d#)) OR
 					(reg_q2615 AND symb_decoder(16#21#)) OR
 					(reg_q2615 AND symb_decoder(16#3c#)) OR
 					(reg_q2615 AND symb_decoder(16#a1#)) OR
 					(reg_q2615 AND symb_decoder(16#9d#)) OR
 					(reg_q2615 AND symb_decoder(16#11#)) OR
 					(reg_q2615 AND symb_decoder(16#ee#)) OR
 					(reg_q2615 AND symb_decoder(16#af#)) OR
 					(reg_q2615 AND symb_decoder(16#8d#)) OR
 					(reg_q2615 AND symb_decoder(16#1c#)) OR
 					(reg_q2615 AND symb_decoder(16#fc#)) OR
 					(reg_q2615 AND symb_decoder(16#4d#)) OR
 					(reg_q2615 AND symb_decoder(16#01#)) OR
 					(reg_q2615 AND symb_decoder(16#02#)) OR
 					(reg_q2615 AND symb_decoder(16#c8#)) OR
 					(reg_q2615 AND symb_decoder(16#95#)) OR
 					(reg_q2615 AND symb_decoder(16#b1#)) OR
 					(reg_q2615 AND symb_decoder(16#bd#)) OR
 					(reg_q2615 AND symb_decoder(16#5c#)) OR
 					(reg_q2615 AND symb_decoder(16#59#)) OR
 					(reg_q2615 AND symb_decoder(16#15#)) OR
 					(reg_q2615 AND symb_decoder(16#52#)) OR
 					(reg_q2615 AND symb_decoder(16#82#)) OR
 					(reg_q2615 AND symb_decoder(16#ae#)) OR
 					(reg_q2615 AND symb_decoder(16#b4#)) OR
 					(reg_q2615 AND symb_decoder(16#61#)) OR
 					(reg_q2615 AND symb_decoder(16#f0#)) OR
 					(reg_q2615 AND symb_decoder(16#2d#)) OR
 					(reg_q2615 AND symb_decoder(16#44#)) OR
 					(reg_q2615 AND symb_decoder(16#7e#)) OR
 					(reg_q2615 AND symb_decoder(16#41#)) OR
 					(reg_q2615 AND symb_decoder(16#31#)) OR
 					(reg_q2615 AND symb_decoder(16#5e#)) OR
 					(reg_q2615 AND symb_decoder(16#85#)) OR
 					(reg_q2615 AND symb_decoder(16#72#)) OR
 					(reg_q2615 AND symb_decoder(16#75#)) OR
 					(reg_q2615 AND symb_decoder(16#d4#)) OR
 					(reg_q2615 AND symb_decoder(16#6b#)) OR
 					(reg_q2615 AND symb_decoder(16#9e#)) OR
 					(reg_q2615 AND symb_decoder(16#28#)) OR
 					(reg_q2615 AND symb_decoder(16#cf#)) OR
 					(reg_q2615 AND symb_decoder(16#4a#)) OR
 					(reg_q2615 AND symb_decoder(16#e2#)) OR
 					(reg_q2615 AND symb_decoder(16#1f#)) OR
 					(reg_q2615 AND symb_decoder(16#9b#)) OR
 					(reg_q2615 AND symb_decoder(16#f2#)) OR
 					(reg_q2615 AND symb_decoder(16#bc#)) OR
 					(reg_q2615 AND symb_decoder(16#26#)) OR
 					(reg_q2615 AND symb_decoder(16#4e#)) OR
 					(reg_q2615 AND symb_decoder(16#2e#)) OR
 					(reg_q2615 AND symb_decoder(16#f8#)) OR
 					(reg_q2615 AND symb_decoder(16#67#)) OR
 					(reg_q2615 AND symb_decoder(16#3a#)) OR
 					(reg_q2615 AND symb_decoder(16#83#)) OR
 					(reg_q2615 AND symb_decoder(16#12#)) OR
 					(reg_q2615 AND symb_decoder(16#b6#)) OR
 					(reg_q2615 AND symb_decoder(16#e8#)) OR
 					(reg_q2615 AND symb_decoder(16#0f#)) OR
 					(reg_q2615 AND symb_decoder(16#94#)) OR
 					(reg_q2615 AND symb_decoder(16#1e#)) OR
 					(reg_q2615 AND symb_decoder(16#2f#)) OR
 					(reg_q2615 AND symb_decoder(16#98#)) OR
 					(reg_q2615 AND symb_decoder(16#42#)) OR
 					(reg_q2615 AND symb_decoder(16#0e#)) OR
 					(reg_q2615 AND symb_decoder(16#ff#)) OR
 					(reg_q2615 AND symb_decoder(16#c4#)) OR
 					(reg_q2615 AND symb_decoder(16#2a#)) OR
 					(reg_q2615 AND symb_decoder(16#6c#)) OR
 					(reg_q2615 AND symb_decoder(16#09#)) OR
 					(reg_q2615 AND symb_decoder(16#5f#)) OR
 					(reg_q2615 AND symb_decoder(16#91#)) OR
 					(reg_q2615 AND symb_decoder(16#00#)) OR
 					(reg_q2615 AND symb_decoder(16#6a#)) OR
 					(reg_q2615 AND symb_decoder(16#43#)) OR
 					(reg_q2615 AND symb_decoder(16#03#)) OR
 					(reg_q2615 AND symb_decoder(16#8f#)) OR
 					(reg_q2615 AND symb_decoder(16#ea#)) OR
 					(reg_q2615 AND symb_decoder(16#87#)) OR
 					(reg_q2615 AND symb_decoder(16#d5#)) OR
 					(reg_q2615 AND symb_decoder(16#25#)) OR
 					(reg_q2615 AND symb_decoder(16#e5#)) OR
 					(reg_q2615 AND symb_decoder(16#3b#)) OR
 					(reg_q2615 AND symb_decoder(16#e3#)) OR
 					(reg_q2615 AND symb_decoder(16#23#)) OR
 					(reg_q2615 AND symb_decoder(16#77#)) OR
 					(reg_q2615 AND symb_decoder(16#b3#)) OR
 					(reg_q2615 AND symb_decoder(16#18#)) OR
 					(reg_q2615 AND symb_decoder(16#46#)) OR
 					(reg_q2615 AND symb_decoder(16#37#)) OR
 					(reg_q2615 AND symb_decoder(16#a0#)) OR
 					(reg_q2615 AND symb_decoder(16#a2#)) OR
 					(reg_q2615 AND symb_decoder(16#8b#)) OR
 					(reg_q2615 AND symb_decoder(16#69#)) OR
 					(reg_q2615 AND symb_decoder(16#0b#)) OR
 					(reg_q2615 AND symb_decoder(16#ed#)) OR
 					(reg_q2615 AND symb_decoder(16#c1#)) OR
 					(reg_q2615 AND symb_decoder(16#30#)) OR
 					(reg_q2615 AND symb_decoder(16#db#)) OR
 					(reg_q2615 AND symb_decoder(16#48#)) OR
 					(reg_q2615 AND symb_decoder(16#a4#)) OR
 					(reg_q2615 AND symb_decoder(16#13#)) OR
 					(reg_q2615 AND symb_decoder(16#e4#)) OR
 					(reg_q2615 AND symb_decoder(16#17#)) OR
 					(reg_q2615 AND symb_decoder(16#89#)) OR
 					(reg_q2615 AND symb_decoder(16#7a#)) OR
 					(reg_q2615 AND symb_decoder(16#d6#)) OR
 					(reg_q2615 AND symb_decoder(16#36#)) OR
 					(reg_q2615 AND symb_decoder(16#5b#)) OR
 					(reg_q2615 AND symb_decoder(16#32#)) OR
 					(reg_q2615 AND symb_decoder(16#05#)) OR
 					(reg_q2615 AND symb_decoder(16#8a#)) OR
 					(reg_q2615 AND symb_decoder(16#20#)) OR
 					(reg_q2615 AND symb_decoder(16#5d#)) OR
 					(reg_q2615 AND symb_decoder(16#b9#)) OR
 					(reg_q2615 AND symb_decoder(16#3e#)) OR
 					(reg_q2615 AND symb_decoder(16#53#)) OR
 					(reg_q2615 AND symb_decoder(16#64#)) OR
 					(reg_q2615 AND symb_decoder(16#99#)) OR
 					(reg_q2615 AND symb_decoder(16#51#)) OR
 					(reg_q2615 AND symb_decoder(16#fd#)) OR
 					(reg_q2615 AND symb_decoder(16#f4#)) OR
 					(reg_q2615 AND symb_decoder(16#62#)) OR
 					(reg_q2615 AND symb_decoder(16#92#)) OR
 					(reg_q2615 AND symb_decoder(16#35#)) OR
 					(reg_q2615 AND symb_decoder(16#50#)) OR
 					(reg_q2615 AND symb_decoder(16#c6#)) OR
 					(reg_q2615 AND symb_decoder(16#33#)) OR
 					(reg_q2615 AND symb_decoder(16#60#)) OR
 					(reg_q2615 AND symb_decoder(16#97#)) OR
 					(reg_q2615 AND symb_decoder(16#f6#)) OR
 					(reg_q2615 AND symb_decoder(16#b2#)) OR
 					(reg_q2615 AND symb_decoder(16#55#)) OR
 					(reg_q2615 AND symb_decoder(16#d1#)) OR
 					(reg_q2615 AND symb_decoder(16#66#)) OR
 					(reg_q2615 AND symb_decoder(16#b0#)) OR
 					(reg_q2615 AND symb_decoder(16#04#)) OR
 					(reg_q2615 AND symb_decoder(16#d7#)) OR
 					(reg_q2615 AND symb_decoder(16#70#)) OR
 					(reg_q2615 AND symb_decoder(16#2b#)) OR
 					(reg_q2615 AND symb_decoder(16#63#)) OR
 					(reg_q2615 AND symb_decoder(16#d0#)) OR
 					(reg_q2615 AND symb_decoder(16#8e#)) OR
 					(reg_q2615 AND symb_decoder(16#7c#)) OR
 					(reg_q2615 AND symb_decoder(16#7d#)) OR
 					(reg_q2615 AND symb_decoder(16#4b#)) OR
 					(reg_q2615 AND symb_decoder(16#10#)) OR
 					(reg_q2615 AND symb_decoder(16#79#)) OR
 					(reg_q2615 AND symb_decoder(16#9f#)) OR
 					(reg_q2615 AND symb_decoder(16#e7#)) OR
 					(reg_q2615 AND symb_decoder(16#fa#)) OR
 					(reg_q2615 AND symb_decoder(16#6d#)) OR
 					(reg_q2615 AND symb_decoder(16#d2#)) OR
 					(reg_q2615 AND symb_decoder(16#08#)) OR
 					(reg_q2615 AND symb_decoder(16#e6#)) OR
 					(reg_q2615 AND symb_decoder(16#38#)) OR
 					(reg_q2615 AND symb_decoder(16#56#)) OR
 					(reg_q2615 AND symb_decoder(16#86#)) OR
 					(reg_q2615 AND symb_decoder(16#dd#)) OR
 					(reg_q2615 AND symb_decoder(16#ba#)) OR
 					(reg_q2615 AND symb_decoder(16#47#)) OR
 					(reg_q2615 AND symb_decoder(16#39#)) OR
 					(reg_q2615 AND symb_decoder(16#a6#)) OR
 					(reg_q2615 AND symb_decoder(16#07#)) OR
 					(reg_q2615 AND symb_decoder(16#9a#)) OR
 					(reg_q2615 AND symb_decoder(16#73#)) OR
 					(reg_q2615 AND symb_decoder(16#c7#)) OR
 					(reg_q2615 AND symb_decoder(16#d8#)) OR
 					(reg_q2615 AND symb_decoder(16#bb#)) OR
 					(reg_q2615 AND symb_decoder(16#06#)) OR
 					(reg_q2615 AND symb_decoder(16#90#)) OR
 					(reg_q2615 AND symb_decoder(16#80#)) OR
 					(reg_q2615 AND symb_decoder(16#2c#)) OR
 					(reg_q2615 AND symb_decoder(16#29#)) OR
 					(reg_q2615 AND symb_decoder(16#b8#)) OR
 					(reg_q2615 AND symb_decoder(16#96#)) OR
 					(reg_q2615 AND symb_decoder(16#c3#)) OR
 					(reg_q2615 AND symb_decoder(16#c0#)) OR
 					(reg_q2615 AND symb_decoder(16#eb#)) OR
 					(reg_q2615 AND symb_decoder(16#9c#)) OR
 					(reg_q2615 AND symb_decoder(16#d3#)) OR
 					(reg_q2615 AND symb_decoder(16#0c#)) OR
 					(reg_q2615 AND symb_decoder(16#5a#)) OR
 					(reg_q2615 AND symb_decoder(16#58#)) OR
 					(reg_q2615 AND symb_decoder(16#ef#)) OR
 					(reg_q2615 AND symb_decoder(16#76#)) OR
 					(reg_q2615 AND symb_decoder(16#45#)) OR
 					(reg_q2615 AND symb_decoder(16#e0#)) OR
 					(reg_q2615 AND symb_decoder(16#de#)) OR
 					(reg_q2615 AND symb_decoder(16#1d#)) OR
 					(reg_q2615 AND symb_decoder(16#df#)) OR
 					(reg_q2615 AND symb_decoder(16#cb#)) OR
 					(reg_q2615 AND symb_decoder(16#7f#)) OR
 					(reg_q2615 AND symb_decoder(16#c5#)) OR
 					(reg_q2615 AND symb_decoder(16#71#)) OR
 					(reg_q2615 AND symb_decoder(16#40#)) OR
 					(reg_q2615 AND symb_decoder(16#8c#)) OR
 					(reg_q2615 AND symb_decoder(16#16#)) OR
 					(reg_q2615 AND symb_decoder(16#6e#)) OR
 					(reg_q2615 AND symb_decoder(16#fe#)) OR
 					(reg_q2615 AND symb_decoder(16#ec#)) OR
 					(reg_q2615 AND symb_decoder(16#88#)) OR
 					(reg_q2615 AND symb_decoder(16#1a#)) OR
 					(reg_q2615 AND symb_decoder(16#81#)) OR
 					(reg_q2615 AND symb_decoder(16#ca#)) OR
 					(reg_q2615 AND symb_decoder(16#7b#)) OR
 					(reg_q2615 AND symb_decoder(16#f7#)) OR
 					(reg_q2615 AND symb_decoder(16#a3#)) OR
 					(reg_q2615 AND symb_decoder(16#aa#)) OR
 					(reg_q2615 AND symb_decoder(16#a5#)) OR
 					(reg_q2615 AND symb_decoder(16#a7#)) OR
 					(reg_q2615 AND symb_decoder(16#1b#)) OR
 					(reg_q2615 AND symb_decoder(16#ce#)) OR
 					(reg_q2615 AND symb_decoder(16#84#)) OR
 					(reg_q2615 AND symb_decoder(16#dc#)) OR
 					(reg_q2615 AND symb_decoder(16#ac#)) OR
 					(reg_q2615 AND symb_decoder(16#24#)) OR
 					(reg_q2615 AND symb_decoder(16#f1#)) OR
 					(reg_q2615 AND symb_decoder(16#f3#)) OR
 					(reg_q2615 AND symb_decoder(16#4c#)) OR
 					(reg_q2615 AND symb_decoder(16#f5#)) OR
 					(reg_q2615 AND symb_decoder(16#f9#)) OR
 					(reg_q2615 AND symb_decoder(16#3f#)) OR
 					(reg_q2615 AND symb_decoder(16#74#)) OR
 					(reg_q2615 AND symb_decoder(16#27#)) OR
 					(reg_q2615 AND symb_decoder(16#49#)) OR
 					(reg_q2615 AND symb_decoder(16#14#)) OR
 					(reg_q2615 AND symb_decoder(16#bf#)) OR
 					(reg_q2615 AND symb_decoder(16#6f#)) OR
 					(reg_q2615 AND symb_decoder(16#65#)) OR
 					(reg_q2615 AND symb_decoder(16#c2#)) OR
 					(reg_q2615 AND symb_decoder(16#cc#)) OR
 					(reg_q2615 AND symb_decoder(16#e9#)) OR
 					(reg_q2615 AND symb_decoder(16#da#)) OR
 					(reg_q2615 AND symb_decoder(16#ad#)) OR
 					(reg_q2615 AND symb_decoder(16#93#)) OR
 					(reg_q2615 AND symb_decoder(16#c9#)) OR
 					(reg_q2615 AND symb_decoder(16#68#)) OR
 					(reg_q2615 AND symb_decoder(16#fb#)) OR
 					(reg_q2615 AND symb_decoder(16#be#)) OR
 					(reg_q2615 AND symb_decoder(16#cd#)) OR
 					(reg_q2615 AND symb_decoder(16#54#)) OR
 					(reg_q2615 AND symb_decoder(16#a8#)) OR
 					(reg_q2615 AND symb_decoder(16#57#)) OR
 					(reg_q2615 AND symb_decoder(16#19#)) OR
 					(reg_q2615 AND symb_decoder(16#22#)) OR
 					(reg_q2615 AND symb_decoder(16#ab#));
reg_q1112_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1111 AND symb_decoder(16#0a#)) OR
 					(reg_q1111 AND symb_decoder(16#0d#));
reg_q953_in <= (reg_q951 AND symb_decoder(16#00#));
reg_q2504_in <= (reg_q2502 AND symb_decoder(16#50#));
reg_q2506_in <= (reg_q2504 AND symb_decoder(16#4f#));
reg_q2510_in <= (reg_q2508 AND symb_decoder(16#54#));
reg_q2491_in <= (reg_q2489 AND symb_decoder(16#52#));
reg_q2485_in <= (reg_q2695 AND symb_decoder(16#2a#));
reg_fullgraph10_init <= "0000";

reg_fullgraph10_sel <= "00000000" & reg_q2485_in & reg_q2491_in & reg_q2510_in & reg_q2506_in & reg_q2504_in & reg_q953_in & reg_q1112_in & reg_q2615_in;

	--coder fullgraph10
with reg_fullgraph10_sel select
reg_fullgraph10_in <=
	"0001" when "0000000000000001",
	"0010" when "0000000000000010",
	"0011" when "0000000000000100",
	"0100" when "0000000000001000",
	"0101" when "0000000000010000",
	"0110" when "0000000000100000",
	"0111" when "0000000001000000",
	"1000" when "0000000010000000",
	"0000" when others;
 --end coder

	p_reg_fullgraph10: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph10 <= reg_fullgraph10_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph10 <= reg_fullgraph10_init;
        else
          reg_fullgraph10 <= reg_fullgraph10_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph10

		reg_q2615 <= '1' when reg_fullgraph10 = "0001" else '0'; 
		reg_q1112 <= '1' when reg_fullgraph10 = "0010" else '0'; 
		reg_q953 <= '1' when reg_fullgraph10 = "0011" else '0'; 
		reg_q2504 <= '1' when reg_fullgraph10 = "0100" else '0'; 
		reg_q2506 <= '1' when reg_fullgraph10 = "0101" else '0'; 
		reg_q2510 <= '1' when reg_fullgraph10 = "0110" else '0'; 
		reg_q2491 <= '1' when reg_fullgraph10 = "0111" else '0'; 
		reg_q2485 <= '1' when reg_fullgraph10 = "1000" else '0'; 
--end decoder 

reg_q1359_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1359 AND symb_decoder(16#47#)) OR
 					(reg_q1359 AND symb_decoder(16#54#)) OR
 					(reg_q1359 AND symb_decoder(16#cd#)) OR
 					(reg_q1359 AND symb_decoder(16#46#)) OR
 					(reg_q1359 AND symb_decoder(16#a3#)) OR
 					(reg_q1359 AND symb_decoder(16#de#)) OR
 					(reg_q1359 AND symb_decoder(16#3f#)) OR
 					(reg_q1359 AND symb_decoder(16#37#)) OR
 					(reg_q1359 AND symb_decoder(16#f0#)) OR
 					(reg_q1359 AND symb_decoder(16#ef#)) OR
 					(reg_q1359 AND symb_decoder(16#25#)) OR
 					(reg_q1359 AND symb_decoder(16#3b#)) OR
 					(reg_q1359 AND symb_decoder(16#ac#)) OR
 					(reg_q1359 AND symb_decoder(16#48#)) OR
 					(reg_q1359 AND symb_decoder(16#bb#)) OR
 					(reg_q1359 AND symb_decoder(16#c0#)) OR
 					(reg_q1359 AND symb_decoder(16#68#)) OR
 					(reg_q1359 AND symb_decoder(16#a4#)) OR
 					(reg_q1359 AND symb_decoder(16#79#)) OR
 					(reg_q1359 AND symb_decoder(16#8f#)) OR
 					(reg_q1359 AND symb_decoder(16#19#)) OR
 					(reg_q1359 AND symb_decoder(16#d9#)) OR
 					(reg_q1359 AND symb_decoder(16#b8#)) OR
 					(reg_q1359 AND symb_decoder(16#27#)) OR
 					(reg_q1359 AND symb_decoder(16#94#)) OR
 					(reg_q1359 AND symb_decoder(16#d5#)) OR
 					(reg_q1359 AND symb_decoder(16#ff#)) OR
 					(reg_q1359 AND symb_decoder(16#ae#)) OR
 					(reg_q1359 AND symb_decoder(16#7d#)) OR
 					(reg_q1359 AND symb_decoder(16#b4#)) OR
 					(reg_q1359 AND symb_decoder(16#5e#)) OR
 					(reg_q1359 AND symb_decoder(16#92#)) OR
 					(reg_q1359 AND symb_decoder(16#b7#)) OR
 					(reg_q1359 AND symb_decoder(16#dd#)) OR
 					(reg_q1359 AND symb_decoder(16#01#)) OR
 					(reg_q1359 AND symb_decoder(16#23#)) OR
 					(reg_q1359 AND symb_decoder(16#f3#)) OR
 					(reg_q1359 AND symb_decoder(16#99#)) OR
 					(reg_q1359 AND symb_decoder(16#da#)) OR
 					(reg_q1359 AND symb_decoder(16#61#)) OR
 					(reg_q1359 AND symb_decoder(16#41#)) OR
 					(reg_q1359 AND symb_decoder(16#29#)) OR
 					(reg_q1359 AND symb_decoder(16#60#)) OR
 					(reg_q1359 AND symb_decoder(16#07#)) OR
 					(reg_q1359 AND symb_decoder(16#ba#)) OR
 					(reg_q1359 AND symb_decoder(16#12#)) OR
 					(reg_q1359 AND symb_decoder(16#d2#)) OR
 					(reg_q1359 AND symb_decoder(16#8c#)) OR
 					(reg_q1359 AND symb_decoder(16#cb#)) OR
 					(reg_q1359 AND symb_decoder(16#4a#)) OR
 					(reg_q1359 AND symb_decoder(16#11#)) OR
 					(reg_q1359 AND symb_decoder(16#95#)) OR
 					(reg_q1359 AND symb_decoder(16#2a#)) OR
 					(reg_q1359 AND symb_decoder(16#d6#)) OR
 					(reg_q1359 AND symb_decoder(16#9e#)) OR
 					(reg_q1359 AND symb_decoder(16#dc#)) OR
 					(reg_q1359 AND symb_decoder(16#ed#)) OR
 					(reg_q1359 AND symb_decoder(16#50#)) OR
 					(reg_q1359 AND symb_decoder(16#3d#)) OR
 					(reg_q1359 AND symb_decoder(16#1f#)) OR
 					(reg_q1359 AND symb_decoder(16#38#)) OR
 					(reg_q1359 AND symb_decoder(16#fd#)) OR
 					(reg_q1359 AND symb_decoder(16#d4#)) OR
 					(reg_q1359 AND symb_decoder(16#d8#)) OR
 					(reg_q1359 AND symb_decoder(16#ec#)) OR
 					(reg_q1359 AND symb_decoder(16#13#)) OR
 					(reg_q1359 AND symb_decoder(16#f2#)) OR
 					(reg_q1359 AND symb_decoder(16#aa#)) OR
 					(reg_q1359 AND symb_decoder(16#7e#)) OR
 					(reg_q1359 AND symb_decoder(16#4b#)) OR
 					(reg_q1359 AND symb_decoder(16#fc#)) OR
 					(reg_q1359 AND symb_decoder(16#17#)) OR
 					(reg_q1359 AND symb_decoder(16#78#)) OR
 					(reg_q1359 AND symb_decoder(16#0d#)) OR
 					(reg_q1359 AND symb_decoder(16#7c#)) OR
 					(reg_q1359 AND symb_decoder(16#6b#)) OR
 					(reg_q1359 AND symb_decoder(16#52#)) OR
 					(reg_q1359 AND symb_decoder(16#03#)) OR
 					(reg_q1359 AND symb_decoder(16#9d#)) OR
 					(reg_q1359 AND symb_decoder(16#88#)) OR
 					(reg_q1359 AND symb_decoder(16#e6#)) OR
 					(reg_q1359 AND symb_decoder(16#ad#)) OR
 					(reg_q1359 AND symb_decoder(16#e1#)) OR
 					(reg_q1359 AND symb_decoder(16#2b#)) OR
 					(reg_q1359 AND symb_decoder(16#b0#)) OR
 					(reg_q1359 AND symb_decoder(16#f5#)) OR
 					(reg_q1359 AND symb_decoder(16#28#)) OR
 					(reg_q1359 AND symb_decoder(16#9f#)) OR
 					(reg_q1359 AND symb_decoder(16#e9#)) OR
 					(reg_q1359 AND symb_decoder(16#db#)) OR
 					(reg_q1359 AND symb_decoder(16#f1#)) OR
 					(reg_q1359 AND symb_decoder(16#c4#)) OR
 					(reg_q1359 AND symb_decoder(16#c7#)) OR
 					(reg_q1359 AND symb_decoder(16#5d#)) OR
 					(reg_q1359 AND symb_decoder(16#85#)) OR
 					(reg_q1359 AND symb_decoder(16#82#)) OR
 					(reg_q1359 AND symb_decoder(16#f7#)) OR
 					(reg_q1359 AND symb_decoder(16#bc#)) OR
 					(reg_q1359 AND symb_decoder(16#f9#)) OR
 					(reg_q1359 AND symb_decoder(16#14#)) OR
 					(reg_q1359 AND symb_decoder(16#93#)) OR
 					(reg_q1359 AND symb_decoder(16#ea#)) OR
 					(reg_q1359 AND symb_decoder(16#1a#)) OR
 					(reg_q1359 AND symb_decoder(16#cc#)) OR
 					(reg_q1359 AND symb_decoder(16#fb#)) OR
 					(reg_q1359 AND symb_decoder(16#96#)) OR
 					(reg_q1359 AND symb_decoder(16#af#)) OR
 					(reg_q1359 AND symb_decoder(16#9b#)) OR
 					(reg_q1359 AND symb_decoder(16#1b#)) OR
 					(reg_q1359 AND symb_decoder(16#56#)) OR
 					(reg_q1359 AND symb_decoder(16#5b#)) OR
 					(reg_q1359 AND symb_decoder(16#f6#)) OR
 					(reg_q1359 AND symb_decoder(16#44#)) OR
 					(reg_q1359 AND symb_decoder(16#b5#)) OR
 					(reg_q1359 AND symb_decoder(16#72#)) OR
 					(reg_q1359 AND symb_decoder(16#08#)) OR
 					(reg_q1359 AND symb_decoder(16#31#)) OR
 					(reg_q1359 AND symb_decoder(16#4c#)) OR
 					(reg_q1359 AND symb_decoder(16#9c#)) OR
 					(reg_q1359 AND symb_decoder(16#87#)) OR
 					(reg_q1359 AND symb_decoder(16#65#)) OR
 					(reg_q1359 AND symb_decoder(16#3c#)) OR
 					(reg_q1359 AND symb_decoder(16#bd#)) OR
 					(reg_q1359 AND symb_decoder(16#2c#)) OR
 					(reg_q1359 AND symb_decoder(16#84#)) OR
 					(reg_q1359 AND symb_decoder(16#5f#)) OR
 					(reg_q1359 AND symb_decoder(16#8a#)) OR
 					(reg_q1359 AND symb_decoder(16#04#)) OR
 					(reg_q1359 AND symb_decoder(16#cf#)) OR
 					(reg_q1359 AND symb_decoder(16#c6#)) OR
 					(reg_q1359 AND symb_decoder(16#73#)) OR
 					(reg_q1359 AND symb_decoder(16#e0#)) OR
 					(reg_q1359 AND symb_decoder(16#0f#)) OR
 					(reg_q1359 AND symb_decoder(16#1c#)) OR
 					(reg_q1359 AND symb_decoder(16#6a#)) OR
 					(reg_q1359 AND symb_decoder(16#4d#)) OR
 					(reg_q1359 AND symb_decoder(16#a5#)) OR
 					(reg_q1359 AND symb_decoder(16#8b#)) OR
 					(reg_q1359 AND symb_decoder(16#c3#)) OR
 					(reg_q1359 AND symb_decoder(16#f4#)) OR
 					(reg_q1359 AND symb_decoder(16#74#)) OR
 					(reg_q1359 AND symb_decoder(16#7f#)) OR
 					(reg_q1359 AND symb_decoder(16#ce#)) OR
 					(reg_q1359 AND symb_decoder(16#b1#)) OR
 					(reg_q1359 AND symb_decoder(16#b3#)) OR
 					(reg_q1359 AND symb_decoder(16#66#)) OR
 					(reg_q1359 AND symb_decoder(16#6e#)) OR
 					(reg_q1359 AND symb_decoder(16#e5#)) OR
 					(reg_q1359 AND symb_decoder(16#81#)) OR
 					(reg_q1359 AND symb_decoder(16#df#)) OR
 					(reg_q1359 AND symb_decoder(16#71#)) OR
 					(reg_q1359 AND symb_decoder(16#0b#)) OR
 					(reg_q1359 AND symb_decoder(16#15#)) OR
 					(reg_q1359 AND symb_decoder(16#d7#)) OR
 					(reg_q1359 AND symb_decoder(16#e7#)) OR
 					(reg_q1359 AND symb_decoder(16#00#)) OR
 					(reg_q1359 AND symb_decoder(16#22#)) OR
 					(reg_q1359 AND symb_decoder(16#20#)) OR
 					(reg_q1359 AND symb_decoder(16#80#)) OR
 					(reg_q1359 AND symb_decoder(16#fe#)) OR
 					(reg_q1359 AND symb_decoder(16#e8#)) OR
 					(reg_q1359 AND symb_decoder(16#c1#)) OR
 					(reg_q1359 AND symb_decoder(16#77#)) OR
 					(reg_q1359 AND symb_decoder(16#5c#)) OR
 					(reg_q1359 AND symb_decoder(16#3a#)) OR
 					(reg_q1359 AND symb_decoder(16#a7#)) OR
 					(reg_q1359 AND symb_decoder(16#63#)) OR
 					(reg_q1359 AND symb_decoder(16#0c#)) OR
 					(reg_q1359 AND symb_decoder(16#1e#)) OR
 					(reg_q1359 AND symb_decoder(16#a9#)) OR
 					(reg_q1359 AND symb_decoder(16#89#)) OR
 					(reg_q1359 AND symb_decoder(16#a8#)) OR
 					(reg_q1359 AND symb_decoder(16#f8#)) OR
 					(reg_q1359 AND symb_decoder(16#49#)) OR
 					(reg_q1359 AND symb_decoder(16#32#)) OR
 					(reg_q1359 AND symb_decoder(16#33#)) OR
 					(reg_q1359 AND symb_decoder(16#6f#)) OR
 					(reg_q1359 AND symb_decoder(16#c8#)) OR
 					(reg_q1359 AND symb_decoder(16#67#)) OR
 					(reg_q1359 AND symb_decoder(16#e3#)) OR
 					(reg_q1359 AND symb_decoder(16#b2#)) OR
 					(reg_q1359 AND symb_decoder(16#86#)) OR
 					(reg_q1359 AND symb_decoder(16#2f#)) OR
 					(reg_q1359 AND symb_decoder(16#42#)) OR
 					(reg_q1359 AND symb_decoder(16#58#)) OR
 					(reg_q1359 AND symb_decoder(16#eb#)) OR
 					(reg_q1359 AND symb_decoder(16#26#)) OR
 					(reg_q1359 AND symb_decoder(16#16#)) OR
 					(reg_q1359 AND symb_decoder(16#59#)) OR
 					(reg_q1359 AND symb_decoder(16#62#)) OR
 					(reg_q1359 AND symb_decoder(16#45#)) OR
 					(reg_q1359 AND symb_decoder(16#8e#)) OR
 					(reg_q1359 AND symb_decoder(16#2e#)) OR
 					(reg_q1359 AND symb_decoder(16#64#)) OR
 					(reg_q1359 AND symb_decoder(16#98#)) OR
 					(reg_q1359 AND symb_decoder(16#4e#)) OR
 					(reg_q1359 AND symb_decoder(16#57#)) OR
 					(reg_q1359 AND symb_decoder(16#9a#)) OR
 					(reg_q1359 AND symb_decoder(16#ca#)) OR
 					(reg_q1359 AND symb_decoder(16#bf#)) OR
 					(reg_q1359 AND symb_decoder(16#06#)) OR
 					(reg_q1359 AND symb_decoder(16#70#)) OR
 					(reg_q1359 AND symb_decoder(16#34#)) OR
 					(reg_q1359 AND symb_decoder(16#91#)) OR
 					(reg_q1359 AND symb_decoder(16#43#)) OR
 					(reg_q1359 AND symb_decoder(16#0a#)) OR
 					(reg_q1359 AND symb_decoder(16#c5#)) OR
 					(reg_q1359 AND symb_decoder(16#b6#)) OR
 					(reg_q1359 AND symb_decoder(16#8d#)) OR
 					(reg_q1359 AND symb_decoder(16#6d#)) OR
 					(reg_q1359 AND symb_decoder(16#be#)) OR
 					(reg_q1359 AND symb_decoder(16#ee#)) OR
 					(reg_q1359 AND symb_decoder(16#a6#)) OR
 					(reg_q1359 AND symb_decoder(16#fa#)) OR
 					(reg_q1359 AND symb_decoder(16#39#)) OR
 					(reg_q1359 AND symb_decoder(16#d3#)) OR
 					(reg_q1359 AND symb_decoder(16#75#)) OR
 					(reg_q1359 AND symb_decoder(16#55#)) OR
 					(reg_q1359 AND symb_decoder(16#6c#)) OR
 					(reg_q1359 AND symb_decoder(16#a2#)) OR
 					(reg_q1359 AND symb_decoder(16#1d#)) OR
 					(reg_q1359 AND symb_decoder(16#02#)) OR
 					(reg_q1359 AND symb_decoder(16#24#)) OR
 					(reg_q1359 AND symb_decoder(16#10#)) OR
 					(reg_q1359 AND symb_decoder(16#0e#)) OR
 					(reg_q1359 AND symb_decoder(16#7a#)) OR
 					(reg_q1359 AND symb_decoder(16#e2#)) OR
 					(reg_q1359 AND symb_decoder(16#83#)) OR
 					(reg_q1359 AND symb_decoder(16#90#)) OR
 					(reg_q1359 AND symb_decoder(16#05#)) OR
 					(reg_q1359 AND symb_decoder(16#ab#)) OR
 					(reg_q1359 AND symb_decoder(16#5a#)) OR
 					(reg_q1359 AND symb_decoder(16#7b#)) OR
 					(reg_q1359 AND symb_decoder(16#97#)) OR
 					(reg_q1359 AND symb_decoder(16#d1#)) OR
 					(reg_q1359 AND symb_decoder(16#51#)) OR
 					(reg_q1359 AND symb_decoder(16#09#)) OR
 					(reg_q1359 AND symb_decoder(16#c9#)) OR
 					(reg_q1359 AND symb_decoder(16#69#)) OR
 					(reg_q1359 AND symb_decoder(16#4f#)) OR
 					(reg_q1359 AND symb_decoder(16#3e#)) OR
 					(reg_q1359 AND symb_decoder(16#c2#)) OR
 					(reg_q1359 AND symb_decoder(16#40#)) OR
 					(reg_q1359 AND symb_decoder(16#d0#)) OR
 					(reg_q1359 AND symb_decoder(16#53#)) OR
 					(reg_q1359 AND symb_decoder(16#18#)) OR
 					(reg_q1359 AND symb_decoder(16#35#)) OR
 					(reg_q1359 AND symb_decoder(16#30#)) OR
 					(reg_q1359 AND symb_decoder(16#e4#)) OR
 					(reg_q1359 AND symb_decoder(16#a0#)) OR
 					(reg_q1359 AND symb_decoder(16#2d#)) OR
 					(reg_q1359 AND symb_decoder(16#b9#)) OR
 					(reg_q1359 AND symb_decoder(16#76#)) OR
 					(reg_q1359 AND symb_decoder(16#36#)) OR
 					(reg_q1359 AND symb_decoder(16#a1#)) OR
 					(reg_q1359 AND symb_decoder(16#21#));
reg_q1359_init <= '0' ;
	p_reg_q1359: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1359 <= reg_q1359_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1359 <= reg_q1359_init;
        else
          reg_q1359 <= reg_q1359_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2618_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2618 AND symb_decoder(16#09#)) OR
 					(reg_q2618 AND symb_decoder(16#0f#)) OR
 					(reg_q2618 AND symb_decoder(16#3f#)) OR
 					(reg_q2618 AND symb_decoder(16#59#)) OR
 					(reg_q2618 AND symb_decoder(16#87#)) OR
 					(reg_q2618 AND symb_decoder(16#98#)) OR
 					(reg_q2618 AND symb_decoder(16#24#)) OR
 					(reg_q2618 AND symb_decoder(16#39#)) OR
 					(reg_q2618 AND symb_decoder(16#ea#)) OR
 					(reg_q2618 AND symb_decoder(16#d4#)) OR
 					(reg_q2618 AND symb_decoder(16#0e#)) OR
 					(reg_q2618 AND symb_decoder(16#5e#)) OR
 					(reg_q2618 AND symb_decoder(16#8f#)) OR
 					(reg_q2618 AND symb_decoder(16#19#)) OR
 					(reg_q2618 AND symb_decoder(16#31#)) OR
 					(reg_q2618 AND symb_decoder(16#f6#)) OR
 					(reg_q2618 AND symb_decoder(16#30#)) OR
 					(reg_q2618 AND symb_decoder(16#82#)) OR
 					(reg_q2618 AND symb_decoder(16#a4#)) OR
 					(reg_q2618 AND symb_decoder(16#c9#)) OR
 					(reg_q2618 AND symb_decoder(16#40#)) OR
 					(reg_q2618 AND symb_decoder(16#9c#)) OR
 					(reg_q2618 AND symb_decoder(16#23#)) OR
 					(reg_q2618 AND symb_decoder(16#bc#)) OR
 					(reg_q2618 AND symb_decoder(16#06#)) OR
 					(reg_q2618 AND symb_decoder(16#b6#)) OR
 					(reg_q2618 AND symb_decoder(16#75#)) OR
 					(reg_q2618 AND symb_decoder(16#52#)) OR
 					(reg_q2618 AND symb_decoder(16#86#)) OR
 					(reg_q2618 AND symb_decoder(16#4f#)) OR
 					(reg_q2618 AND symb_decoder(16#d6#)) OR
 					(reg_q2618 AND symb_decoder(16#89#)) OR
 					(reg_q2618 AND symb_decoder(16#a2#)) OR
 					(reg_q2618 AND symb_decoder(16#28#)) OR
 					(reg_q2618 AND symb_decoder(16#1e#)) OR
 					(reg_q2618 AND symb_decoder(16#5f#)) OR
 					(reg_q2618 AND symb_decoder(16#8b#)) OR
 					(reg_q2618 AND symb_decoder(16#e9#)) OR
 					(reg_q2618 AND symb_decoder(16#ab#)) OR
 					(reg_q2618 AND symb_decoder(16#dd#)) OR
 					(reg_q2618 AND symb_decoder(16#3d#)) OR
 					(reg_q2618 AND symb_decoder(16#65#)) OR
 					(reg_q2618 AND symb_decoder(16#51#)) OR
 					(reg_q2618 AND symb_decoder(16#4b#)) OR
 					(reg_q2618 AND symb_decoder(16#1a#)) OR
 					(reg_q2618 AND symb_decoder(16#53#)) OR
 					(reg_q2618 AND symb_decoder(16#90#)) OR
 					(reg_q2618 AND symb_decoder(16#92#)) OR
 					(reg_q2618 AND symb_decoder(16#04#)) OR
 					(reg_q2618 AND symb_decoder(16#b0#)) OR
 					(reg_q2618 AND symb_decoder(16#e2#)) OR
 					(reg_q2618 AND symb_decoder(16#db#)) OR
 					(reg_q2618 AND symb_decoder(16#94#)) OR
 					(reg_q2618 AND symb_decoder(16#4a#)) OR
 					(reg_q2618 AND symb_decoder(16#34#)) OR
 					(reg_q2618 AND symb_decoder(16#d2#)) OR
 					(reg_q2618 AND symb_decoder(16#80#)) OR
 					(reg_q2618 AND symb_decoder(16#47#)) OR
 					(reg_q2618 AND symb_decoder(16#f0#)) OR
 					(reg_q2618 AND symb_decoder(16#07#)) OR
 					(reg_q2618 AND symb_decoder(16#ae#)) OR
 					(reg_q2618 AND symb_decoder(16#b3#)) OR
 					(reg_q2618 AND symb_decoder(16#46#)) OR
 					(reg_q2618 AND symb_decoder(16#ce#)) OR
 					(reg_q2618 AND symb_decoder(16#33#)) OR
 					(reg_q2618 AND symb_decoder(16#d3#)) OR
 					(reg_q2618 AND symb_decoder(16#d1#)) OR
 					(reg_q2618 AND symb_decoder(16#fb#)) OR
 					(reg_q2618 AND symb_decoder(16#05#)) OR
 					(reg_q2618 AND symb_decoder(16#6a#)) OR
 					(reg_q2618 AND symb_decoder(16#f7#)) OR
 					(reg_q2618 AND symb_decoder(16#ad#)) OR
 					(reg_q2618 AND symb_decoder(16#42#)) OR
 					(reg_q2618 AND symb_decoder(16#ac#)) OR
 					(reg_q2618 AND symb_decoder(16#be#)) OR
 					(reg_q2618 AND symb_decoder(16#1b#)) OR
 					(reg_q2618 AND symb_decoder(16#de#)) OR
 					(reg_q2618 AND symb_decoder(16#ec#)) OR
 					(reg_q2618 AND symb_decoder(16#18#)) OR
 					(reg_q2618 AND symb_decoder(16#96#)) OR
 					(reg_q2618 AND symb_decoder(16#97#)) OR
 					(reg_q2618 AND symb_decoder(16#ef#)) OR
 					(reg_q2618 AND symb_decoder(16#ba#)) OR
 					(reg_q2618 AND symb_decoder(16#54#)) OR
 					(reg_q2618 AND symb_decoder(16#cd#)) OR
 					(reg_q2618 AND symb_decoder(16#66#)) OR
 					(reg_q2618 AND symb_decoder(16#bd#)) OR
 					(reg_q2618 AND symb_decoder(16#64#)) OR
 					(reg_q2618 AND symb_decoder(16#eb#)) OR
 					(reg_q2618 AND symb_decoder(16#6f#)) OR
 					(reg_q2618 AND symb_decoder(16#b1#)) OR
 					(reg_q2618 AND symb_decoder(16#9b#)) OR
 					(reg_q2618 AND symb_decoder(16#b5#)) OR
 					(reg_q2618 AND symb_decoder(16#63#)) OR
 					(reg_q2618 AND symb_decoder(16#f3#)) OR
 					(reg_q2618 AND symb_decoder(16#55#)) OR
 					(reg_q2618 AND symb_decoder(16#8e#)) OR
 					(reg_q2618 AND symb_decoder(16#af#)) OR
 					(reg_q2618 AND symb_decoder(16#61#)) OR
 					(reg_q2618 AND symb_decoder(16#72#)) OR
 					(reg_q2618 AND symb_decoder(16#b8#)) OR
 					(reg_q2618 AND symb_decoder(16#a1#)) OR
 					(reg_q2618 AND symb_decoder(16#5c#)) OR
 					(reg_q2618 AND symb_decoder(16#b7#)) OR
 					(reg_q2618 AND symb_decoder(16#5d#)) OR
 					(reg_q2618 AND symb_decoder(16#6c#)) OR
 					(reg_q2618 AND symb_decoder(16#3e#)) OR
 					(reg_q2618 AND symb_decoder(16#5a#)) OR
 					(reg_q2618 AND symb_decoder(16#0b#)) OR
 					(reg_q2618 AND symb_decoder(16#1f#)) OR
 					(reg_q2618 AND symb_decoder(16#7d#)) OR
 					(reg_q2618 AND symb_decoder(16#7b#)) OR
 					(reg_q2618 AND symb_decoder(16#71#)) OR
 					(reg_q2618 AND symb_decoder(16#29#)) OR
 					(reg_q2618 AND symb_decoder(16#fa#)) OR
 					(reg_q2618 AND symb_decoder(16#69#)) OR
 					(reg_q2618 AND symb_decoder(16#14#)) OR
 					(reg_q2618 AND symb_decoder(16#02#)) OR
 					(reg_q2618 AND symb_decoder(16#8d#)) OR
 					(reg_q2618 AND symb_decoder(16#f9#)) OR
 					(reg_q2618 AND symb_decoder(16#bf#)) OR
 					(reg_q2618 AND symb_decoder(16#fc#)) OR
 					(reg_q2618 AND symb_decoder(16#e5#)) OR
 					(reg_q2618 AND symb_decoder(16#e3#)) OR
 					(reg_q2618 AND symb_decoder(16#88#)) OR
 					(reg_q2618 AND symb_decoder(16#01#)) OR
 					(reg_q2618 AND symb_decoder(16#78#)) OR
 					(reg_q2618 AND symb_decoder(16#d7#)) OR
 					(reg_q2618 AND symb_decoder(16#cb#)) OR
 					(reg_q2618 AND symb_decoder(16#fe#)) OR
 					(reg_q2618 AND symb_decoder(16#9f#)) OR
 					(reg_q2618 AND symb_decoder(16#44#)) OR
 					(reg_q2618 AND symb_decoder(16#68#)) OR
 					(reg_q2618 AND symb_decoder(16#4c#)) OR
 					(reg_q2618 AND symb_decoder(16#cc#)) OR
 					(reg_q2618 AND symb_decoder(16#a7#)) OR
 					(reg_q2618 AND symb_decoder(16#83#)) OR
 					(reg_q2618 AND symb_decoder(16#32#)) OR
 					(reg_q2618 AND symb_decoder(16#56#)) OR
 					(reg_q2618 AND symb_decoder(16#62#)) OR
 					(reg_q2618 AND symb_decoder(16#aa#)) OR
 					(reg_q2618 AND symb_decoder(16#58#)) OR
 					(reg_q2618 AND symb_decoder(16#ff#)) OR
 					(reg_q2618 AND symb_decoder(16#b9#)) OR
 					(reg_q2618 AND symb_decoder(16#0c#)) OR
 					(reg_q2618 AND symb_decoder(16#4e#)) OR
 					(reg_q2618 AND symb_decoder(16#c2#)) OR
 					(reg_q2618 AND symb_decoder(16#67#)) OR
 					(reg_q2618 AND symb_decoder(16#15#)) OR
 					(reg_q2618 AND symb_decoder(16#a0#)) OR
 					(reg_q2618 AND symb_decoder(16#0a#)) OR
 					(reg_q2618 AND symb_decoder(16#c3#)) OR
 					(reg_q2618 AND symb_decoder(16#e6#)) OR
 					(reg_q2618 AND symb_decoder(16#f2#)) OR
 					(reg_q2618 AND symb_decoder(16#2e#)) OR
 					(reg_q2618 AND symb_decoder(16#16#)) OR
 					(reg_q2618 AND symb_decoder(16#00#)) OR
 					(reg_q2618 AND symb_decoder(16#7c#)) OR
 					(reg_q2618 AND symb_decoder(16#27#)) OR
 					(reg_q2618 AND symb_decoder(16#11#)) OR
 					(reg_q2618 AND symb_decoder(16#c1#)) OR
 					(reg_q2618 AND symb_decoder(16#ca#)) OR
 					(reg_q2618 AND symb_decoder(16#8a#)) OR
 					(reg_q2618 AND symb_decoder(16#e4#)) OR
 					(reg_q2618 AND symb_decoder(16#99#)) OR
 					(reg_q2618 AND symb_decoder(16#f1#)) OR
 					(reg_q2618 AND symb_decoder(16#93#)) OR
 					(reg_q2618 AND symb_decoder(16#4d#)) OR
 					(reg_q2618 AND symb_decoder(16#dc#)) OR
 					(reg_q2618 AND symb_decoder(16#c0#)) OR
 					(reg_q2618 AND symb_decoder(16#95#)) OR
 					(reg_q2618 AND symb_decoder(16#ed#)) OR
 					(reg_q2618 AND symb_decoder(16#03#)) OR
 					(reg_q2618 AND symb_decoder(16#f4#)) OR
 					(reg_q2618 AND symb_decoder(16#f8#)) OR
 					(reg_q2618 AND symb_decoder(16#0d#)) OR
 					(reg_q2618 AND symb_decoder(16#b2#)) OR
 					(reg_q2618 AND symb_decoder(16#c4#)) OR
 					(reg_q2618 AND symb_decoder(16#12#)) OR
 					(reg_q2618 AND symb_decoder(16#73#)) OR
 					(reg_q2618 AND symb_decoder(16#17#)) OR
 					(reg_q2618 AND symb_decoder(16#60#)) OR
 					(reg_q2618 AND symb_decoder(16#b4#)) OR
 					(reg_q2618 AND symb_decoder(16#22#)) OR
 					(reg_q2618 AND symb_decoder(16#e8#)) OR
 					(reg_q2618 AND symb_decoder(16#37#)) OR
 					(reg_q2618 AND symb_decoder(16#3b#)) OR
 					(reg_q2618 AND symb_decoder(16#84#)) OR
 					(reg_q2618 AND symb_decoder(16#10#)) OR
 					(reg_q2618 AND symb_decoder(16#70#)) OR
 					(reg_q2618 AND symb_decoder(16#43#)) OR
 					(reg_q2618 AND symb_decoder(16#20#)) OR
 					(reg_q2618 AND symb_decoder(16#45#)) OR
 					(reg_q2618 AND symb_decoder(16#d9#)) OR
 					(reg_q2618 AND symb_decoder(16#a8#)) OR
 					(reg_q2618 AND symb_decoder(16#cf#)) OR
 					(reg_q2618 AND symb_decoder(16#26#)) OR
 					(reg_q2618 AND symb_decoder(16#9a#)) OR
 					(reg_q2618 AND symb_decoder(16#df#)) OR
 					(reg_q2618 AND symb_decoder(16#1c#)) OR
 					(reg_q2618 AND symb_decoder(16#9d#)) OR
 					(reg_q2618 AND symb_decoder(16#13#)) OR
 					(reg_q2618 AND symb_decoder(16#6e#)) OR
 					(reg_q2618 AND symb_decoder(16#91#)) OR
 					(reg_q2618 AND symb_decoder(16#57#)) OR
 					(reg_q2618 AND symb_decoder(16#77#)) OR
 					(reg_q2618 AND symb_decoder(16#3c#)) OR
 					(reg_q2618 AND symb_decoder(16#41#)) OR
 					(reg_q2618 AND symb_decoder(16#9e#)) OR
 					(reg_q2618 AND symb_decoder(16#6b#)) OR
 					(reg_q2618 AND symb_decoder(16#81#)) OR
 					(reg_q2618 AND symb_decoder(16#2c#)) OR
 					(reg_q2618 AND symb_decoder(16#c7#)) OR
 					(reg_q2618 AND symb_decoder(16#da#)) OR
 					(reg_q2618 AND symb_decoder(16#a3#)) OR
 					(reg_q2618 AND symb_decoder(16#ee#)) OR
 					(reg_q2618 AND symb_decoder(16#49#)) OR
 					(reg_q2618 AND symb_decoder(16#e0#)) OR
 					(reg_q2618 AND symb_decoder(16#85#)) OR
 					(reg_q2618 AND symb_decoder(16#bb#)) OR
 					(reg_q2618 AND symb_decoder(16#50#)) OR
 					(reg_q2618 AND symb_decoder(16#e7#)) OR
 					(reg_q2618 AND symb_decoder(16#7f#)) OR
 					(reg_q2618 AND symb_decoder(16#d8#)) OR
 					(reg_q2618 AND symb_decoder(16#7e#)) OR
 					(reg_q2618 AND symb_decoder(16#1d#)) OR
 					(reg_q2618 AND symb_decoder(16#fd#)) OR
 					(reg_q2618 AND symb_decoder(16#a6#)) OR
 					(reg_q2618 AND symb_decoder(16#c5#)) OR
 					(reg_q2618 AND symb_decoder(16#d0#)) OR
 					(reg_q2618 AND symb_decoder(16#38#)) OR
 					(reg_q2618 AND symb_decoder(16#36#)) OR
 					(reg_q2618 AND symb_decoder(16#c6#)) OR
 					(reg_q2618 AND symb_decoder(16#48#)) OR
 					(reg_q2618 AND symb_decoder(16#6d#)) OR
 					(reg_q2618 AND symb_decoder(16#74#)) OR
 					(reg_q2618 AND symb_decoder(16#5b#)) OR
 					(reg_q2618 AND symb_decoder(16#3a#)) OR
 					(reg_q2618 AND symb_decoder(16#25#)) OR
 					(reg_q2618 AND symb_decoder(16#a9#)) OR
 					(reg_q2618 AND symb_decoder(16#f5#)) OR
 					(reg_q2618 AND symb_decoder(16#76#)) OR
 					(reg_q2618 AND symb_decoder(16#d5#)) OR
 					(reg_q2618 AND symb_decoder(16#2b#)) OR
 					(reg_q2618 AND symb_decoder(16#21#)) OR
 					(reg_q2618 AND symb_decoder(16#c8#)) OR
 					(reg_q2618 AND symb_decoder(16#79#)) OR
 					(reg_q2618 AND symb_decoder(16#2f#)) OR
 					(reg_q2618 AND symb_decoder(16#e1#)) OR
 					(reg_q2618 AND symb_decoder(16#08#)) OR
 					(reg_q2618 AND symb_decoder(16#2d#)) OR
 					(reg_q2618 AND symb_decoder(16#35#)) OR
 					(reg_q2618 AND symb_decoder(16#7a#)) OR
 					(reg_q2618 AND symb_decoder(16#8c#)) OR
 					(reg_q2618 AND symb_decoder(16#2a#)) OR
 					(reg_q2618 AND symb_decoder(16#a5#));
reg_q2618_init <= '0' ;
	p_reg_q2618: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2618 <= reg_q2618_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2618 <= reg_q2618_init;
        else
          reg_q2618 <= reg_q2618_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1742_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1742 AND symb_decoder(16#1b#)) OR
 					(reg_q1742 AND symb_decoder(16#6e#)) OR
 					(reg_q1742 AND symb_decoder(16#bb#)) OR
 					(reg_q1742 AND symb_decoder(16#76#)) OR
 					(reg_q1742 AND symb_decoder(16#25#)) OR
 					(reg_q1742 AND symb_decoder(16#5c#)) OR
 					(reg_q1742 AND symb_decoder(16#cd#)) OR
 					(reg_q1742 AND symb_decoder(16#54#)) OR
 					(reg_q1742 AND symb_decoder(16#cc#)) OR
 					(reg_q1742 AND symb_decoder(16#88#)) OR
 					(reg_q1742 AND symb_decoder(16#99#)) OR
 					(reg_q1742 AND symb_decoder(16#2b#)) OR
 					(reg_q1742 AND symb_decoder(16#c9#)) OR
 					(reg_q1742 AND symb_decoder(16#75#)) OR
 					(reg_q1742 AND symb_decoder(16#28#)) OR
 					(reg_q1742 AND symb_decoder(16#05#)) OR
 					(reg_q1742 AND symb_decoder(16#fe#)) OR
 					(reg_q1742 AND symb_decoder(16#e9#)) OR
 					(reg_q1742 AND symb_decoder(16#ea#)) OR
 					(reg_q1742 AND symb_decoder(16#7a#)) OR
 					(reg_q1742 AND symb_decoder(16#2d#)) OR
 					(reg_q1742 AND symb_decoder(16#ce#)) OR
 					(reg_q1742 AND symb_decoder(16#80#)) OR
 					(reg_q1742 AND symb_decoder(16#e2#)) OR
 					(reg_q1742 AND symb_decoder(16#cb#)) OR
 					(reg_q1742 AND symb_decoder(16#d6#)) OR
 					(reg_q1742 AND symb_decoder(16#0e#)) OR
 					(reg_q1742 AND symb_decoder(16#7f#)) OR
 					(reg_q1742 AND symb_decoder(16#0b#)) OR
 					(reg_q1742 AND symb_decoder(16#0a#)) OR
 					(reg_q1742 AND symb_decoder(16#8e#)) OR
 					(reg_q1742 AND symb_decoder(16#0d#)) OR
 					(reg_q1742 AND symb_decoder(16#9f#)) OR
 					(reg_q1742 AND symb_decoder(16#3a#)) OR
 					(reg_q1742 AND symb_decoder(16#bc#)) OR
 					(reg_q1742 AND symb_decoder(16#d3#)) OR
 					(reg_q1742 AND symb_decoder(16#7c#)) OR
 					(reg_q1742 AND symb_decoder(16#32#)) OR
 					(reg_q1742 AND symb_decoder(16#1d#)) OR
 					(reg_q1742 AND symb_decoder(16#12#)) OR
 					(reg_q1742 AND symb_decoder(16#62#)) OR
 					(reg_q1742 AND symb_decoder(16#4a#)) OR
 					(reg_q1742 AND symb_decoder(16#22#)) OR
 					(reg_q1742 AND symb_decoder(16#fc#)) OR
 					(reg_q1742 AND symb_decoder(16#ef#)) OR
 					(reg_q1742 AND symb_decoder(16#3c#)) OR
 					(reg_q1742 AND symb_decoder(16#ff#)) OR
 					(reg_q1742 AND symb_decoder(16#56#)) OR
 					(reg_q1742 AND symb_decoder(16#94#)) OR
 					(reg_q1742 AND symb_decoder(16#b5#)) OR
 					(reg_q1742 AND symb_decoder(16#52#)) OR
 					(reg_q1742 AND symb_decoder(16#ad#)) OR
 					(reg_q1742 AND symb_decoder(16#16#)) OR
 					(reg_q1742 AND symb_decoder(16#e8#)) OR
 					(reg_q1742 AND symb_decoder(16#84#)) OR
 					(reg_q1742 AND symb_decoder(16#38#)) OR
 					(reg_q1742 AND symb_decoder(16#92#)) OR
 					(reg_q1742 AND symb_decoder(16#30#)) OR
 					(reg_q1742 AND symb_decoder(16#ac#)) OR
 					(reg_q1742 AND symb_decoder(16#e4#)) OR
 					(reg_q1742 AND symb_decoder(16#44#)) OR
 					(reg_q1742 AND symb_decoder(16#b6#)) OR
 					(reg_q1742 AND symb_decoder(16#14#)) OR
 					(reg_q1742 AND symb_decoder(16#9b#)) OR
 					(reg_q1742 AND symb_decoder(16#a2#)) OR
 					(reg_q1742 AND symb_decoder(16#67#)) OR
 					(reg_q1742 AND symb_decoder(16#35#)) OR
 					(reg_q1742 AND symb_decoder(16#af#)) OR
 					(reg_q1742 AND symb_decoder(16#0f#)) OR
 					(reg_q1742 AND symb_decoder(16#61#)) OR
 					(reg_q1742 AND symb_decoder(16#23#)) OR
 					(reg_q1742 AND symb_decoder(16#ab#)) OR
 					(reg_q1742 AND symb_decoder(16#41#)) OR
 					(reg_q1742 AND symb_decoder(16#7d#)) OR
 					(reg_q1742 AND symb_decoder(16#06#)) OR
 					(reg_q1742 AND symb_decoder(16#77#)) OR
 					(reg_q1742 AND symb_decoder(16#0c#)) OR
 					(reg_q1742 AND symb_decoder(16#10#)) OR
 					(reg_q1742 AND symb_decoder(16#b1#)) OR
 					(reg_q1742 AND symb_decoder(16#f6#)) OR
 					(reg_q1742 AND symb_decoder(16#37#)) OR
 					(reg_q1742 AND symb_decoder(16#8b#)) OR
 					(reg_q1742 AND symb_decoder(16#11#)) OR
 					(reg_q1742 AND symb_decoder(16#83#)) OR
 					(reg_q1742 AND symb_decoder(16#42#)) OR
 					(reg_q1742 AND symb_decoder(16#c2#)) OR
 					(reg_q1742 AND symb_decoder(16#d5#)) OR
 					(reg_q1742 AND symb_decoder(16#39#)) OR
 					(reg_q1742 AND symb_decoder(16#69#)) OR
 					(reg_q1742 AND symb_decoder(16#b0#)) OR
 					(reg_q1742 AND symb_decoder(16#a8#)) OR
 					(reg_q1742 AND symb_decoder(16#1f#)) OR
 					(reg_q1742 AND symb_decoder(16#5e#)) OR
 					(reg_q1742 AND symb_decoder(16#a9#)) OR
 					(reg_q1742 AND symb_decoder(16#d9#)) OR
 					(reg_q1742 AND symb_decoder(16#f0#)) OR
 					(reg_q1742 AND symb_decoder(16#4e#)) OR
 					(reg_q1742 AND symb_decoder(16#40#)) OR
 					(reg_q1742 AND symb_decoder(16#a7#)) OR
 					(reg_q1742 AND symb_decoder(16#02#)) OR
 					(reg_q1742 AND symb_decoder(16#01#)) OR
 					(reg_q1742 AND symb_decoder(16#d0#)) OR
 					(reg_q1742 AND symb_decoder(16#db#)) OR
 					(reg_q1742 AND symb_decoder(16#86#)) OR
 					(reg_q1742 AND symb_decoder(16#09#)) OR
 					(reg_q1742 AND symb_decoder(16#a1#)) OR
 					(reg_q1742 AND symb_decoder(16#2f#)) OR
 					(reg_q1742 AND symb_decoder(16#9a#)) OR
 					(reg_q1742 AND symb_decoder(16#6a#)) OR
 					(reg_q1742 AND symb_decoder(16#5a#)) OR
 					(reg_q1742 AND symb_decoder(16#66#)) OR
 					(reg_q1742 AND symb_decoder(16#46#)) OR
 					(reg_q1742 AND symb_decoder(16#7b#)) OR
 					(reg_q1742 AND symb_decoder(16#fd#)) OR
 					(reg_q1742 AND symb_decoder(16#81#)) OR
 					(reg_q1742 AND symb_decoder(16#d8#)) OR
 					(reg_q1742 AND symb_decoder(16#6f#)) OR
 					(reg_q1742 AND symb_decoder(16#6b#)) OR
 					(reg_q1742 AND symb_decoder(16#df#)) OR
 					(reg_q1742 AND symb_decoder(16#ec#)) OR
 					(reg_q1742 AND symb_decoder(16#48#)) OR
 					(reg_q1742 AND symb_decoder(16#50#)) OR
 					(reg_q1742 AND symb_decoder(16#a3#)) OR
 					(reg_q1742 AND symb_decoder(16#47#)) OR
 					(reg_q1742 AND symb_decoder(16#91#)) OR
 					(reg_q1742 AND symb_decoder(16#27#)) OR
 					(reg_q1742 AND symb_decoder(16#e5#)) OR
 					(reg_q1742 AND symb_decoder(16#ed#)) OR
 					(reg_q1742 AND symb_decoder(16#e1#)) OR
 					(reg_q1742 AND symb_decoder(16#f9#)) OR
 					(reg_q1742 AND symb_decoder(16#bd#)) OR
 					(reg_q1742 AND symb_decoder(16#29#)) OR
 					(reg_q1742 AND symb_decoder(16#a6#)) OR
 					(reg_q1742 AND symb_decoder(16#aa#)) OR
 					(reg_q1742 AND symb_decoder(16#4b#)) OR
 					(reg_q1742 AND symb_decoder(16#fa#)) OR
 					(reg_q1742 AND symb_decoder(16#45#)) OR
 					(reg_q1742 AND symb_decoder(16#18#)) OR
 					(reg_q1742 AND symb_decoder(16#65#)) OR
 					(reg_q1742 AND symb_decoder(16#ca#)) OR
 					(reg_q1742 AND symb_decoder(16#13#)) OR
 					(reg_q1742 AND symb_decoder(16#43#)) OR
 					(reg_q1742 AND symb_decoder(16#4c#)) OR
 					(reg_q1742 AND symb_decoder(16#5b#)) OR
 					(reg_q1742 AND symb_decoder(16#6c#)) OR
 					(reg_q1742 AND symb_decoder(16#3f#)) OR
 					(reg_q1742 AND symb_decoder(16#da#)) OR
 					(reg_q1742 AND symb_decoder(16#90#)) OR
 					(reg_q1742 AND symb_decoder(16#95#)) OR
 					(reg_q1742 AND symb_decoder(16#53#)) OR
 					(reg_q1742 AND symb_decoder(16#19#)) OR
 					(reg_q1742 AND symb_decoder(16#f2#)) OR
 					(reg_q1742 AND symb_decoder(16#c5#)) OR
 					(reg_q1742 AND symb_decoder(16#03#)) OR
 					(reg_q1742 AND symb_decoder(16#72#)) OR
 					(reg_q1742 AND symb_decoder(16#8d#)) OR
 					(reg_q1742 AND symb_decoder(16#7e#)) OR
 					(reg_q1742 AND symb_decoder(16#1c#)) OR
 					(reg_q1742 AND symb_decoder(16#e3#)) OR
 					(reg_q1742 AND symb_decoder(16#6d#)) OR
 					(reg_q1742 AND symb_decoder(16#97#)) OR
 					(reg_q1742 AND symb_decoder(16#e0#)) OR
 					(reg_q1742 AND symb_decoder(16#15#)) OR
 					(reg_q1742 AND symb_decoder(16#5d#)) OR
 					(reg_q1742 AND symb_decoder(16#ee#)) OR
 					(reg_q1742 AND symb_decoder(16#d1#)) OR
 					(reg_q1742 AND symb_decoder(16#f1#)) OR
 					(reg_q1742 AND symb_decoder(16#c8#)) OR
 					(reg_q1742 AND symb_decoder(16#e7#)) OR
 					(reg_q1742 AND symb_decoder(16#70#)) OR
 					(reg_q1742 AND symb_decoder(16#60#)) OR
 					(reg_q1742 AND symb_decoder(16#31#)) OR
 					(reg_q1742 AND symb_decoder(16#f7#)) OR
 					(reg_q1742 AND symb_decoder(16#98#)) OR
 					(reg_q1742 AND symb_decoder(16#2a#)) OR
 					(reg_q1742 AND symb_decoder(16#93#)) OR
 					(reg_q1742 AND symb_decoder(16#20#)) OR
 					(reg_q1742 AND symb_decoder(16#a4#)) OR
 					(reg_q1742 AND symb_decoder(16#34#)) OR
 					(reg_q1742 AND symb_decoder(16#51#)) OR
 					(reg_q1742 AND symb_decoder(16#96#)) OR
 					(reg_q1742 AND symb_decoder(16#4d#)) OR
 					(reg_q1742 AND symb_decoder(16#b2#)) OR
 					(reg_q1742 AND symb_decoder(16#33#)) OR
 					(reg_q1742 AND symb_decoder(16#b8#)) OR
 					(reg_q1742 AND symb_decoder(16#58#)) OR
 					(reg_q1742 AND symb_decoder(16#59#)) OR
 					(reg_q1742 AND symb_decoder(16#c7#)) OR
 					(reg_q1742 AND symb_decoder(16#9d#)) OR
 					(reg_q1742 AND symb_decoder(16#d2#)) OR
 					(reg_q1742 AND symb_decoder(16#dd#)) OR
 					(reg_q1742 AND symb_decoder(16#e6#)) OR
 					(reg_q1742 AND symb_decoder(16#3b#)) OR
 					(reg_q1742 AND symb_decoder(16#00#)) OR
 					(reg_q1742 AND symb_decoder(16#8f#)) OR
 					(reg_q1742 AND symb_decoder(16#fb#)) OR
 					(reg_q1742 AND symb_decoder(16#1a#)) OR
 					(reg_q1742 AND symb_decoder(16#f3#)) OR
 					(reg_q1742 AND symb_decoder(16#63#)) OR
 					(reg_q1742 AND symb_decoder(16#64#)) OR
 					(reg_q1742 AND symb_decoder(16#de#)) OR
 					(reg_q1742 AND symb_decoder(16#36#)) OR
 					(reg_q1742 AND symb_decoder(16#57#)) OR
 					(reg_q1742 AND symb_decoder(16#b3#)) OR
 					(reg_q1742 AND symb_decoder(16#85#)) OR
 					(reg_q1742 AND symb_decoder(16#ba#)) OR
 					(reg_q1742 AND symb_decoder(16#21#)) OR
 					(reg_q1742 AND symb_decoder(16#b7#)) OR
 					(reg_q1742 AND symb_decoder(16#3d#)) OR
 					(reg_q1742 AND symb_decoder(16#24#)) OR
 					(reg_q1742 AND symb_decoder(16#cf#)) OR
 					(reg_q1742 AND symb_decoder(16#d7#)) OR
 					(reg_q1742 AND symb_decoder(16#f8#)) OR
 					(reg_q1742 AND symb_decoder(16#9c#)) OR
 					(reg_q1742 AND symb_decoder(16#bf#)) OR
 					(reg_q1742 AND symb_decoder(16#74#)) OR
 					(reg_q1742 AND symb_decoder(16#26#)) OR
 					(reg_q1742 AND symb_decoder(16#07#)) OR
 					(reg_q1742 AND symb_decoder(16#d4#)) OR
 					(reg_q1742 AND symb_decoder(16#c0#)) OR
 					(reg_q1742 AND symb_decoder(16#78#)) OR
 					(reg_q1742 AND symb_decoder(16#c6#)) OR
 					(reg_q1742 AND symb_decoder(16#3e#)) OR
 					(reg_q1742 AND symb_decoder(16#8a#)) OR
 					(reg_q1742 AND symb_decoder(16#04#)) OR
 					(reg_q1742 AND symb_decoder(16#c4#)) OR
 					(reg_q1742 AND symb_decoder(16#73#)) OR
 					(reg_q1742 AND symb_decoder(16#1e#)) OR
 					(reg_q1742 AND symb_decoder(16#9e#)) OR
 					(reg_q1742 AND symb_decoder(16#2e#)) OR
 					(reg_q1742 AND symb_decoder(16#8c#)) OR
 					(reg_q1742 AND symb_decoder(16#79#)) OR
 					(reg_q1742 AND symb_decoder(16#f5#)) OR
 					(reg_q1742 AND symb_decoder(16#ae#)) OR
 					(reg_q1742 AND symb_decoder(16#4f#)) OR
 					(reg_q1742 AND symb_decoder(16#17#)) OR
 					(reg_q1742 AND symb_decoder(16#b9#)) OR
 					(reg_q1742 AND symb_decoder(16#a5#)) OR
 					(reg_q1742 AND symb_decoder(16#08#)) OR
 					(reg_q1742 AND symb_decoder(16#eb#)) OR
 					(reg_q1742 AND symb_decoder(16#71#)) OR
 					(reg_q1742 AND symb_decoder(16#c3#)) OR
 					(reg_q1742 AND symb_decoder(16#5f#)) OR
 					(reg_q1742 AND symb_decoder(16#dc#)) OR
 					(reg_q1742 AND symb_decoder(16#2c#)) OR
 					(reg_q1742 AND symb_decoder(16#55#)) OR
 					(reg_q1742 AND symb_decoder(16#f4#)) OR
 					(reg_q1742 AND symb_decoder(16#b4#)) OR
 					(reg_q1742 AND symb_decoder(16#a0#)) OR
 					(reg_q1742 AND symb_decoder(16#c1#)) OR
 					(reg_q1742 AND symb_decoder(16#89#)) OR
 					(reg_q1742 AND symb_decoder(16#82#)) OR
 					(reg_q1742 AND symb_decoder(16#be#)) OR
 					(reg_q1742 AND symb_decoder(16#87#)) OR
 					(reg_q1742 AND symb_decoder(16#49#)) OR
 					(reg_q1742 AND symb_decoder(16#68#));
reg_q1742_init <= '0' ;
	p_reg_q1742: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1742 <= reg_q1742_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1742 <= reg_q1742_init;
        else
          reg_q1742 <= reg_q1742_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2383_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2383 AND symb_decoder(16#f4#)) OR
 					(reg_q2383 AND symb_decoder(16#38#)) OR
 					(reg_q2383 AND symb_decoder(16#4d#)) OR
 					(reg_q2383 AND symb_decoder(16#ce#)) OR
 					(reg_q2383 AND symb_decoder(16#09#)) OR
 					(reg_q2383 AND symb_decoder(16#79#)) OR
 					(reg_q2383 AND symb_decoder(16#5b#)) OR
 					(reg_q2383 AND symb_decoder(16#3f#)) OR
 					(reg_q2383 AND symb_decoder(16#04#)) OR
 					(reg_q2383 AND symb_decoder(16#a9#)) OR
 					(reg_q2383 AND symb_decoder(16#4c#)) OR
 					(reg_q2383 AND symb_decoder(16#63#)) OR
 					(reg_q2383 AND symb_decoder(16#2c#)) OR
 					(reg_q2383 AND symb_decoder(16#85#)) OR
 					(reg_q2383 AND symb_decoder(16#c4#)) OR
 					(reg_q2383 AND symb_decoder(16#fd#)) OR
 					(reg_q2383 AND symb_decoder(16#0e#)) OR
 					(reg_q2383 AND symb_decoder(16#e2#)) OR
 					(reg_q2383 AND symb_decoder(16#e7#)) OR
 					(reg_q2383 AND symb_decoder(16#ab#)) OR
 					(reg_q2383 AND symb_decoder(16#08#)) OR
 					(reg_q2383 AND symb_decoder(16#94#)) OR
 					(reg_q2383 AND symb_decoder(16#e0#)) OR
 					(reg_q2383 AND symb_decoder(16#7f#)) OR
 					(reg_q2383 AND symb_decoder(16#06#)) OR
 					(reg_q2383 AND symb_decoder(16#de#)) OR
 					(reg_q2383 AND symb_decoder(16#d5#)) OR
 					(reg_q2383 AND symb_decoder(16#70#)) OR
 					(reg_q2383 AND symb_decoder(16#2e#)) OR
 					(reg_q2383 AND symb_decoder(16#2b#)) OR
 					(reg_q2383 AND symb_decoder(16#05#)) OR
 					(reg_q2383 AND symb_decoder(16#25#)) OR
 					(reg_q2383 AND symb_decoder(16#78#)) OR
 					(reg_q2383 AND symb_decoder(16#c2#)) OR
 					(reg_q2383 AND symb_decoder(16#dd#)) OR
 					(reg_q2383 AND symb_decoder(16#27#)) OR
 					(reg_q2383 AND symb_decoder(16#d8#)) OR
 					(reg_q2383 AND symb_decoder(16#cc#)) OR
 					(reg_q2383 AND symb_decoder(16#48#)) OR
 					(reg_q2383 AND symb_decoder(16#8b#)) OR
 					(reg_q2383 AND symb_decoder(16#16#)) OR
 					(reg_q2383 AND symb_decoder(16#29#)) OR
 					(reg_q2383 AND symb_decoder(16#90#)) OR
 					(reg_q2383 AND symb_decoder(16#5c#)) OR
 					(reg_q2383 AND symb_decoder(16#ec#)) OR
 					(reg_q2383 AND symb_decoder(16#98#)) OR
 					(reg_q2383 AND symb_decoder(16#3b#)) OR
 					(reg_q2383 AND symb_decoder(16#6b#)) OR
 					(reg_q2383 AND symb_decoder(16#ff#)) OR
 					(reg_q2383 AND symb_decoder(16#80#)) OR
 					(reg_q2383 AND symb_decoder(16#37#)) OR
 					(reg_q2383 AND symb_decoder(16#74#)) OR
 					(reg_q2383 AND symb_decoder(16#54#)) OR
 					(reg_q2383 AND symb_decoder(16#cd#)) OR
 					(reg_q2383 AND symb_decoder(16#a4#)) OR
 					(reg_q2383 AND symb_decoder(16#01#)) OR
 					(reg_q2383 AND symb_decoder(16#8c#)) OR
 					(reg_q2383 AND symb_decoder(16#6e#)) OR
 					(reg_q2383 AND symb_decoder(16#43#)) OR
 					(reg_q2383 AND symb_decoder(16#76#)) OR
 					(reg_q2383 AND symb_decoder(16#67#)) OR
 					(reg_q2383 AND symb_decoder(16#ea#)) OR
 					(reg_q2383 AND symb_decoder(16#eb#)) OR
 					(reg_q2383 AND symb_decoder(16#b2#)) OR
 					(reg_q2383 AND symb_decoder(16#28#)) OR
 					(reg_q2383 AND symb_decoder(16#81#)) OR
 					(reg_q2383 AND symb_decoder(16#9d#)) OR
 					(reg_q2383 AND symb_decoder(16#17#)) OR
 					(reg_q2383 AND symb_decoder(16#14#)) OR
 					(reg_q2383 AND symb_decoder(16#e5#)) OR
 					(reg_q2383 AND symb_decoder(16#1e#)) OR
 					(reg_q2383 AND symb_decoder(16#c3#)) OR
 					(reg_q2383 AND symb_decoder(16#97#)) OR
 					(reg_q2383 AND symb_decoder(16#83#)) OR
 					(reg_q2383 AND symb_decoder(16#b1#)) OR
 					(reg_q2383 AND symb_decoder(16#1b#)) OR
 					(reg_q2383 AND symb_decoder(16#7d#)) OR
 					(reg_q2383 AND symb_decoder(16#9f#)) OR
 					(reg_q2383 AND symb_decoder(16#1d#)) OR
 					(reg_q2383 AND symb_decoder(16#d2#)) OR
 					(reg_q2383 AND symb_decoder(16#db#)) OR
 					(reg_q2383 AND symb_decoder(16#d4#)) OR
 					(reg_q2383 AND symb_decoder(16#6d#)) OR
 					(reg_q2383 AND symb_decoder(16#a2#)) OR
 					(reg_q2383 AND symb_decoder(16#3c#)) OR
 					(reg_q2383 AND symb_decoder(16#6a#)) OR
 					(reg_q2383 AND symb_decoder(16#0c#)) OR
 					(reg_q2383 AND symb_decoder(16#ef#)) OR
 					(reg_q2383 AND symb_decoder(16#b9#)) OR
 					(reg_q2383 AND symb_decoder(16#41#)) OR
 					(reg_q2383 AND symb_decoder(16#2a#)) OR
 					(reg_q2383 AND symb_decoder(16#57#)) OR
 					(reg_q2383 AND symb_decoder(16#9a#)) OR
 					(reg_q2383 AND symb_decoder(16#89#)) OR
 					(reg_q2383 AND symb_decoder(16#13#)) OR
 					(reg_q2383 AND symb_decoder(16#d7#)) OR
 					(reg_q2383 AND symb_decoder(16#36#)) OR
 					(reg_q2383 AND symb_decoder(16#e6#)) OR
 					(reg_q2383 AND symb_decoder(16#c5#)) OR
 					(reg_q2383 AND symb_decoder(16#f0#)) OR
 					(reg_q2383 AND symb_decoder(16#b6#)) OR
 					(reg_q2383 AND symb_decoder(16#65#)) OR
 					(reg_q2383 AND symb_decoder(16#47#)) OR
 					(reg_q2383 AND symb_decoder(16#61#)) OR
 					(reg_q2383 AND symb_decoder(16#fb#)) OR
 					(reg_q2383 AND symb_decoder(16#7a#)) OR
 					(reg_q2383 AND symb_decoder(16#53#)) OR
 					(reg_q2383 AND symb_decoder(16#03#)) OR
 					(reg_q2383 AND symb_decoder(16#aa#)) OR
 					(reg_q2383 AND symb_decoder(16#42#)) OR
 					(reg_q2383 AND symb_decoder(16#b3#)) OR
 					(reg_q2383 AND symb_decoder(16#73#)) OR
 					(reg_q2383 AND symb_decoder(16#c1#)) OR
 					(reg_q2383 AND symb_decoder(16#c8#)) OR
 					(reg_q2383 AND symb_decoder(16#f2#)) OR
 					(reg_q2383 AND symb_decoder(16#e3#)) OR
 					(reg_q2383 AND symb_decoder(16#56#)) OR
 					(reg_q2383 AND symb_decoder(16#2d#)) OR
 					(reg_q2383 AND symb_decoder(16#9b#)) OR
 					(reg_q2383 AND symb_decoder(16#a7#)) OR
 					(reg_q2383 AND symb_decoder(16#1c#)) OR
 					(reg_q2383 AND symb_decoder(16#a5#)) OR
 					(reg_q2383 AND symb_decoder(16#50#)) OR
 					(reg_q2383 AND symb_decoder(16#23#)) OR
 					(reg_q2383 AND symb_decoder(16#64#)) OR
 					(reg_q2383 AND symb_decoder(16#ca#)) OR
 					(reg_q2383 AND symb_decoder(16#df#)) OR
 					(reg_q2383 AND symb_decoder(16#f3#)) OR
 					(reg_q2383 AND symb_decoder(16#b0#)) OR
 					(reg_q2383 AND symb_decoder(16#a0#)) OR
 					(reg_q2383 AND symb_decoder(16#bf#)) OR
 					(reg_q2383 AND symb_decoder(16#bd#)) OR
 					(reg_q2383 AND symb_decoder(16#51#)) OR
 					(reg_q2383 AND symb_decoder(16#4f#)) OR
 					(reg_q2383 AND symb_decoder(16#7e#)) OR
 					(reg_q2383 AND symb_decoder(16#af#)) OR
 					(reg_q2383 AND symb_decoder(16#6f#)) OR
 					(reg_q2383 AND symb_decoder(16#c6#)) OR
 					(reg_q2383 AND symb_decoder(16#88#)) OR
 					(reg_q2383 AND symb_decoder(16#35#)) OR
 					(reg_q2383 AND symb_decoder(16#4a#)) OR
 					(reg_q2383 AND symb_decoder(16#f9#)) OR
 					(reg_q2383 AND symb_decoder(16#7b#)) OR
 					(reg_q2383 AND symb_decoder(16#00#)) OR
 					(reg_q2383 AND symb_decoder(16#58#)) OR
 					(reg_q2383 AND symb_decoder(16#3a#)) OR
 					(reg_q2383 AND symb_decoder(16#77#)) OR
 					(reg_q2383 AND symb_decoder(16#e4#)) OR
 					(reg_q2383 AND symb_decoder(16#9c#)) OR
 					(reg_q2383 AND symb_decoder(16#92#)) OR
 					(reg_q2383 AND symb_decoder(16#f8#)) OR
 					(reg_q2383 AND symb_decoder(16#5d#)) OR
 					(reg_q2383 AND symb_decoder(16#c0#)) OR
 					(reg_q2383 AND symb_decoder(16#d6#)) OR
 					(reg_q2383 AND symb_decoder(16#30#)) OR
 					(reg_q2383 AND symb_decoder(16#11#)) OR
 					(reg_q2383 AND symb_decoder(16#a3#)) OR
 					(reg_q2383 AND symb_decoder(16#ed#)) OR
 					(reg_q2383 AND symb_decoder(16#d0#)) OR
 					(reg_q2383 AND symb_decoder(16#72#)) OR
 					(reg_q2383 AND symb_decoder(16#cf#)) OR
 					(reg_q2383 AND symb_decoder(16#ac#)) OR
 					(reg_q2383 AND symb_decoder(16#55#)) OR
 					(reg_q2383 AND symb_decoder(16#da#)) OR
 					(reg_q2383 AND symb_decoder(16#fa#)) OR
 					(reg_q2383 AND symb_decoder(16#ba#)) OR
 					(reg_q2383 AND symb_decoder(16#d1#)) OR
 					(reg_q2383 AND symb_decoder(16#40#)) OR
 					(reg_q2383 AND symb_decoder(16#46#)) OR
 					(reg_q2383 AND symb_decoder(16#b4#)) OR
 					(reg_q2383 AND symb_decoder(16#5e#)) OR
 					(reg_q2383 AND symb_decoder(16#99#)) OR
 					(reg_q2383 AND symb_decoder(16#33#)) OR
 					(reg_q2383 AND symb_decoder(16#fe#)) OR
 					(reg_q2383 AND symb_decoder(16#69#)) OR
 					(reg_q2383 AND symb_decoder(16#26#)) OR
 					(reg_q2383 AND symb_decoder(16#66#)) OR
 					(reg_q2383 AND symb_decoder(16#34#)) OR
 					(reg_q2383 AND symb_decoder(16#e9#)) OR
 					(reg_q2383 AND symb_decoder(16#18#)) OR
 					(reg_q2383 AND symb_decoder(16#dc#)) OR
 					(reg_q2383 AND symb_decoder(16#a6#)) OR
 					(reg_q2383 AND symb_decoder(16#8e#)) OR
 					(reg_q2383 AND symb_decoder(16#87#)) OR
 					(reg_q2383 AND symb_decoder(16#95#)) OR
 					(reg_q2383 AND symb_decoder(16#84#)) OR
 					(reg_q2383 AND symb_decoder(16#f1#)) OR
 					(reg_q2383 AND symb_decoder(16#21#)) OR
 					(reg_q2383 AND symb_decoder(16#f5#)) OR
 					(reg_q2383 AND symb_decoder(16#c9#)) OR
 					(reg_q2383 AND symb_decoder(16#31#)) OR
 					(reg_q2383 AND symb_decoder(16#62#)) OR
 					(reg_q2383 AND symb_decoder(16#5f#)) OR
 					(reg_q2383 AND symb_decoder(16#e1#)) OR
 					(reg_q2383 AND symb_decoder(16#b7#)) OR
 					(reg_q2383 AND symb_decoder(16#0f#)) OR
 					(reg_q2383 AND symb_decoder(16#a8#)) OR
 					(reg_q2383 AND symb_decoder(16#8f#)) OR
 					(reg_q2383 AND symb_decoder(16#19#)) OR
 					(reg_q2383 AND symb_decoder(16#6c#)) OR
 					(reg_q2383 AND symb_decoder(16#bb#)) OR
 					(reg_q2383 AND symb_decoder(16#10#)) OR
 					(reg_q2383 AND symb_decoder(16#22#)) OR
 					(reg_q2383 AND symb_decoder(16#ee#)) OR
 					(reg_q2383 AND symb_decoder(16#3e#)) OR
 					(reg_q2383 AND symb_decoder(16#93#)) OR
 					(reg_q2383 AND symb_decoder(16#d9#)) OR
 					(reg_q2383 AND symb_decoder(16#bc#)) OR
 					(reg_q2383 AND symb_decoder(16#fc#)) OR
 					(reg_q2383 AND symb_decoder(16#1f#)) OR
 					(reg_q2383 AND symb_decoder(16#0d#)) OR
 					(reg_q2383 AND symb_decoder(16#68#)) OR
 					(reg_q2383 AND symb_decoder(16#32#)) OR
 					(reg_q2383 AND symb_decoder(16#02#)) OR
 					(reg_q2383 AND symb_decoder(16#c7#)) OR
 					(reg_q2383 AND symb_decoder(16#8a#)) OR
 					(reg_q2383 AND symb_decoder(16#b5#)) OR
 					(reg_q2383 AND symb_decoder(16#2f#)) OR
 					(reg_q2383 AND symb_decoder(16#44#)) OR
 					(reg_q2383 AND symb_decoder(16#8d#)) OR
 					(reg_q2383 AND symb_decoder(16#91#)) OR
 					(reg_q2383 AND symb_decoder(16#1a#)) OR
 					(reg_q2383 AND symb_decoder(16#b8#)) OR
 					(reg_q2383 AND symb_decoder(16#59#)) OR
 					(reg_q2383 AND symb_decoder(16#ae#)) OR
 					(reg_q2383 AND symb_decoder(16#39#)) OR
 					(reg_q2383 AND symb_decoder(16#0a#)) OR
 					(reg_q2383 AND symb_decoder(16#5a#)) OR
 					(reg_q2383 AND symb_decoder(16#0b#)) OR
 					(reg_q2383 AND symb_decoder(16#82#)) OR
 					(reg_q2383 AND symb_decoder(16#cb#)) OR
 					(reg_q2383 AND symb_decoder(16#4e#)) OR
 					(reg_q2383 AND symb_decoder(16#d3#)) OR
 					(reg_q2383 AND symb_decoder(16#20#)) OR
 					(reg_q2383 AND symb_decoder(16#52#)) OR
 					(reg_q2383 AND symb_decoder(16#75#)) OR
 					(reg_q2383 AND symb_decoder(16#a1#)) OR
 					(reg_q2383 AND symb_decoder(16#4b#)) OR
 					(reg_q2383 AND symb_decoder(16#49#)) OR
 					(reg_q2383 AND symb_decoder(16#86#)) OR
 					(reg_q2383 AND symb_decoder(16#12#)) OR
 					(reg_q2383 AND symb_decoder(16#7c#)) OR
 					(reg_q2383 AND symb_decoder(16#60#)) OR
 					(reg_q2383 AND symb_decoder(16#e8#)) OR
 					(reg_q2383 AND symb_decoder(16#9e#)) OR
 					(reg_q2383 AND symb_decoder(16#ad#)) OR
 					(reg_q2383 AND symb_decoder(16#24#)) OR
 					(reg_q2383 AND symb_decoder(16#f7#)) OR
 					(reg_q2383 AND symb_decoder(16#45#)) OR
 					(reg_q2383 AND symb_decoder(16#15#)) OR
 					(reg_q2383 AND symb_decoder(16#3d#)) OR
 					(reg_q2383 AND symb_decoder(16#f6#)) OR
 					(reg_q2383 AND symb_decoder(16#be#)) OR
 					(reg_q2383 AND symb_decoder(16#07#)) OR
 					(reg_q2383 AND symb_decoder(16#71#)) OR
 					(reg_q2383 AND symb_decoder(16#96#));
reg_q2383_init <= '0' ;
	p_reg_q2383: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2383 <= reg_q2383_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2383 <= reg_q2383_init;
        else
          reg_q2383 <= reg_q2383_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2124_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2124 AND symb_decoder(16#25#)) OR
 					(reg_q2124 AND symb_decoder(16#f6#)) OR
 					(reg_q2124 AND symb_decoder(16#fc#)) OR
 					(reg_q2124 AND symb_decoder(16#40#)) OR
 					(reg_q2124 AND symb_decoder(16#f4#)) OR
 					(reg_q2124 AND symb_decoder(16#51#)) OR
 					(reg_q2124 AND symb_decoder(16#0f#)) OR
 					(reg_q2124 AND symb_decoder(16#57#)) OR
 					(reg_q2124 AND symb_decoder(16#17#)) OR
 					(reg_q2124 AND symb_decoder(16#2f#)) OR
 					(reg_q2124 AND symb_decoder(16#03#)) OR
 					(reg_q2124 AND symb_decoder(16#22#)) OR
 					(reg_q2124 AND symb_decoder(16#5f#)) OR
 					(reg_q2124 AND symb_decoder(16#cd#)) OR
 					(reg_q2124 AND symb_decoder(16#54#)) OR
 					(reg_q2124 AND symb_decoder(16#8c#)) OR
 					(reg_q2124 AND symb_decoder(16#65#)) OR
 					(reg_q2124 AND symb_decoder(16#e1#)) OR
 					(reg_q2124 AND symb_decoder(16#bc#)) OR
 					(reg_q2124 AND symb_decoder(16#0d#)) OR
 					(reg_q2124 AND symb_decoder(16#bd#)) OR
 					(reg_q2124 AND symb_decoder(16#df#)) OR
 					(reg_q2124 AND symb_decoder(16#5d#)) OR
 					(reg_q2124 AND symb_decoder(16#66#)) OR
 					(reg_q2124 AND symb_decoder(16#ed#)) OR
 					(reg_q2124 AND symb_decoder(16#b9#)) OR
 					(reg_q2124 AND symb_decoder(16#0a#)) OR
 					(reg_q2124 AND symb_decoder(16#30#)) OR
 					(reg_q2124 AND symb_decoder(16#27#)) OR
 					(reg_q2124 AND symb_decoder(16#fb#)) OR
 					(reg_q2124 AND symb_decoder(16#4b#)) OR
 					(reg_q2124 AND symb_decoder(16#15#)) OR
 					(reg_q2124 AND symb_decoder(16#23#)) OR
 					(reg_q2124 AND symb_decoder(16#12#)) OR
 					(reg_q2124 AND symb_decoder(16#18#)) OR
 					(reg_q2124 AND symb_decoder(16#47#)) OR
 					(reg_q2124 AND symb_decoder(16#04#)) OR
 					(reg_q2124 AND symb_decoder(16#81#)) OR
 					(reg_q2124 AND symb_decoder(16#ec#)) OR
 					(reg_q2124 AND symb_decoder(16#9a#)) OR
 					(reg_q2124 AND symb_decoder(16#44#)) OR
 					(reg_q2124 AND symb_decoder(16#d0#)) OR
 					(reg_q2124 AND symb_decoder(16#97#)) OR
 					(reg_q2124 AND symb_decoder(16#9c#)) OR
 					(reg_q2124 AND symb_decoder(16#eb#)) OR
 					(reg_q2124 AND symb_decoder(16#1e#)) OR
 					(reg_q2124 AND symb_decoder(16#6a#)) OR
 					(reg_q2124 AND symb_decoder(16#7c#)) OR
 					(reg_q2124 AND symb_decoder(16#6e#)) OR
 					(reg_q2124 AND symb_decoder(16#2c#)) OR
 					(reg_q2124 AND symb_decoder(16#e5#)) OR
 					(reg_q2124 AND symb_decoder(16#ab#)) OR
 					(reg_q2124 AND symb_decoder(16#2d#)) OR
 					(reg_q2124 AND symb_decoder(16#09#)) OR
 					(reg_q2124 AND symb_decoder(16#ce#)) OR
 					(reg_q2124 AND symb_decoder(16#cb#)) OR
 					(reg_q2124 AND symb_decoder(16#16#)) OR
 					(reg_q2124 AND symb_decoder(16#46#)) OR
 					(reg_q2124 AND symb_decoder(16#4e#)) OR
 					(reg_q2124 AND symb_decoder(16#f1#)) OR
 					(reg_q2124 AND symb_decoder(16#41#)) OR
 					(reg_q2124 AND symb_decoder(16#76#)) OR
 					(reg_q2124 AND symb_decoder(16#cf#)) OR
 					(reg_q2124 AND symb_decoder(16#c1#)) OR
 					(reg_q2124 AND symb_decoder(16#c5#)) OR
 					(reg_q2124 AND symb_decoder(16#0c#)) OR
 					(reg_q2124 AND symb_decoder(16#b6#)) OR
 					(reg_q2124 AND symb_decoder(16#87#)) OR
 					(reg_q2124 AND symb_decoder(16#9b#)) OR
 					(reg_q2124 AND symb_decoder(16#d4#)) OR
 					(reg_q2124 AND symb_decoder(16#ca#)) OR
 					(reg_q2124 AND symb_decoder(16#11#)) OR
 					(reg_q2124 AND symb_decoder(16#b0#)) OR
 					(reg_q2124 AND symb_decoder(16#9d#)) OR
 					(reg_q2124 AND symb_decoder(16#2a#)) OR
 					(reg_q2124 AND symb_decoder(16#43#)) OR
 					(reg_q2124 AND symb_decoder(16#b5#)) OR
 					(reg_q2124 AND symb_decoder(16#c8#)) OR
 					(reg_q2124 AND symb_decoder(16#b7#)) OR
 					(reg_q2124 AND symb_decoder(16#ba#)) OR
 					(reg_q2124 AND symb_decoder(16#e2#)) OR
 					(reg_q2124 AND symb_decoder(16#37#)) OR
 					(reg_q2124 AND symb_decoder(16#fd#)) OR
 					(reg_q2124 AND symb_decoder(16#60#)) OR
 					(reg_q2124 AND symb_decoder(16#a1#)) OR
 					(reg_q2124 AND symb_decoder(16#cc#)) OR
 					(reg_q2124 AND symb_decoder(16#7d#)) OR
 					(reg_q2124 AND symb_decoder(16#ea#)) OR
 					(reg_q2124 AND symb_decoder(16#f8#)) OR
 					(reg_q2124 AND symb_decoder(16#84#)) OR
 					(reg_q2124 AND symb_decoder(16#8a#)) OR
 					(reg_q2124 AND symb_decoder(16#75#)) OR
 					(reg_q2124 AND symb_decoder(16#f2#)) OR
 					(reg_q2124 AND symb_decoder(16#e0#)) OR
 					(reg_q2124 AND symb_decoder(16#82#)) OR
 					(reg_q2124 AND symb_decoder(16#ee#)) OR
 					(reg_q2124 AND symb_decoder(16#53#)) OR
 					(reg_q2124 AND symb_decoder(16#55#)) OR
 					(reg_q2124 AND symb_decoder(16#6b#)) OR
 					(reg_q2124 AND symb_decoder(16#d2#)) OR
 					(reg_q2124 AND symb_decoder(16#34#)) OR
 					(reg_q2124 AND symb_decoder(16#67#)) OR
 					(reg_q2124 AND symb_decoder(16#a0#)) OR
 					(reg_q2124 AND symb_decoder(16#62#)) OR
 					(reg_q2124 AND symb_decoder(16#d9#)) OR
 					(reg_q2124 AND symb_decoder(16#8e#)) OR
 					(reg_q2124 AND symb_decoder(16#88#)) OR
 					(reg_q2124 AND symb_decoder(16#e7#)) OR
 					(reg_q2124 AND symb_decoder(16#aa#)) OR
 					(reg_q2124 AND symb_decoder(16#fa#)) OR
 					(reg_q2124 AND symb_decoder(16#f5#)) OR
 					(reg_q2124 AND symb_decoder(16#f7#)) OR
 					(reg_q2124 AND symb_decoder(16#92#)) OR
 					(reg_q2124 AND symb_decoder(16#21#)) OR
 					(reg_q2124 AND symb_decoder(16#bb#)) OR
 					(reg_q2124 AND symb_decoder(16#4d#)) OR
 					(reg_q2124 AND symb_decoder(16#d3#)) OR
 					(reg_q2124 AND symb_decoder(16#35#)) OR
 					(reg_q2124 AND symb_decoder(16#e3#)) OR
 					(reg_q2124 AND symb_decoder(16#6c#)) OR
 					(reg_q2124 AND symb_decoder(16#85#)) OR
 					(reg_q2124 AND symb_decoder(16#89#)) OR
 					(reg_q2124 AND symb_decoder(16#c6#)) OR
 					(reg_q2124 AND symb_decoder(16#8b#)) OR
 					(reg_q2124 AND symb_decoder(16#32#)) OR
 					(reg_q2124 AND symb_decoder(16#73#)) OR
 					(reg_q2124 AND symb_decoder(16#4c#)) OR
 					(reg_q2124 AND symb_decoder(16#c2#)) OR
 					(reg_q2124 AND symb_decoder(16#9e#)) OR
 					(reg_q2124 AND symb_decoder(16#a5#)) OR
 					(reg_q2124 AND symb_decoder(16#19#)) OR
 					(reg_q2124 AND symb_decoder(16#8f#)) OR
 					(reg_q2124 AND symb_decoder(16#86#)) OR
 					(reg_q2124 AND symb_decoder(16#69#)) OR
 					(reg_q2124 AND symb_decoder(16#5c#)) OR
 					(reg_q2124 AND symb_decoder(16#07#)) OR
 					(reg_q2124 AND symb_decoder(16#13#)) OR
 					(reg_q2124 AND symb_decoder(16#7f#)) OR
 					(reg_q2124 AND symb_decoder(16#3d#)) OR
 					(reg_q2124 AND symb_decoder(16#2e#)) OR
 					(reg_q2124 AND symb_decoder(16#ff#)) OR
 					(reg_q2124 AND symb_decoder(16#36#)) OR
 					(reg_q2124 AND symb_decoder(16#48#)) OR
 					(reg_q2124 AND symb_decoder(16#72#)) OR
 					(reg_q2124 AND symb_decoder(16#91#)) OR
 					(reg_q2124 AND symb_decoder(16#c3#)) OR
 					(reg_q2124 AND symb_decoder(16#98#)) OR
 					(reg_q2124 AND symb_decoder(16#3a#)) OR
 					(reg_q2124 AND symb_decoder(16#b3#)) OR
 					(reg_q2124 AND symb_decoder(16#3b#)) OR
 					(reg_q2124 AND symb_decoder(16#a9#)) OR
 					(reg_q2124 AND symb_decoder(16#a8#)) OR
 					(reg_q2124 AND symb_decoder(16#38#)) OR
 					(reg_q2124 AND symb_decoder(16#e8#)) OR
 					(reg_q2124 AND symb_decoder(16#56#)) OR
 					(reg_q2124 AND symb_decoder(16#1a#)) OR
 					(reg_q2124 AND symb_decoder(16#49#)) OR
 					(reg_q2124 AND symb_decoder(16#77#)) OR
 					(reg_q2124 AND symb_decoder(16#fe#)) OR
 					(reg_q2124 AND symb_decoder(16#de#)) OR
 					(reg_q2124 AND symb_decoder(16#e4#)) OR
 					(reg_q2124 AND symb_decoder(16#b8#)) OR
 					(reg_q2124 AND symb_decoder(16#2b#)) OR
 					(reg_q2124 AND symb_decoder(16#4f#)) OR
 					(reg_q2124 AND symb_decoder(16#7b#)) OR
 					(reg_q2124 AND symb_decoder(16#a3#)) OR
 					(reg_q2124 AND symb_decoder(16#d8#)) OR
 					(reg_q2124 AND symb_decoder(16#71#)) OR
 					(reg_q2124 AND symb_decoder(16#5e#)) OR
 					(reg_q2124 AND symb_decoder(16#31#)) OR
 					(reg_q2124 AND symb_decoder(16#b1#)) OR
 					(reg_q2124 AND symb_decoder(16#7e#)) OR
 					(reg_q2124 AND symb_decoder(16#0e#)) OR
 					(reg_q2124 AND symb_decoder(16#28#)) OR
 					(reg_q2124 AND symb_decoder(16#20#)) OR
 					(reg_q2124 AND symb_decoder(16#05#)) OR
 					(reg_q2124 AND symb_decoder(16#a7#)) OR
 					(reg_q2124 AND symb_decoder(16#d5#)) OR
 					(reg_q2124 AND symb_decoder(16#af#)) OR
 					(reg_q2124 AND symb_decoder(16#39#)) OR
 					(reg_q2124 AND symb_decoder(16#29#)) OR
 					(reg_q2124 AND symb_decoder(16#79#)) OR
 					(reg_q2124 AND symb_decoder(16#bf#)) OR
 					(reg_q2124 AND symb_decoder(16#5a#)) OR
 					(reg_q2124 AND symb_decoder(16#78#)) OR
 					(reg_q2124 AND symb_decoder(16#83#)) OR
 					(reg_q2124 AND symb_decoder(16#4a#)) OR
 					(reg_q2124 AND symb_decoder(16#c9#)) OR
 					(reg_q2124 AND symb_decoder(16#be#)) OR
 					(reg_q2124 AND symb_decoder(16#02#)) OR
 					(reg_q2124 AND symb_decoder(16#00#)) OR
 					(reg_q2124 AND symb_decoder(16#b4#)) OR
 					(reg_q2124 AND symb_decoder(16#01#)) OR
 					(reg_q2124 AND symb_decoder(16#6d#)) OR
 					(reg_q2124 AND symb_decoder(16#c4#)) OR
 					(reg_q2124 AND symb_decoder(16#9f#)) OR
 					(reg_q2124 AND symb_decoder(16#64#)) OR
 					(reg_q2124 AND symb_decoder(16#59#)) OR
 					(reg_q2124 AND symb_decoder(16#33#)) OR
 					(reg_q2124 AND symb_decoder(16#1b#)) OR
 					(reg_q2124 AND symb_decoder(16#d6#)) OR
 					(reg_q2124 AND symb_decoder(16#24#)) OR
 					(reg_q2124 AND symb_decoder(16#5b#)) OR
 					(reg_q2124 AND symb_decoder(16#1d#)) OR
 					(reg_q2124 AND symb_decoder(16#e6#)) OR
 					(reg_q2124 AND symb_decoder(16#42#)) OR
 					(reg_q2124 AND symb_decoder(16#06#)) OR
 					(reg_q2124 AND symb_decoder(16#94#)) OR
 					(reg_q2124 AND symb_decoder(16#95#)) OR
 					(reg_q2124 AND symb_decoder(16#61#)) OR
 					(reg_q2124 AND symb_decoder(16#c7#)) OR
 					(reg_q2124 AND symb_decoder(16#70#)) OR
 					(reg_q2124 AND symb_decoder(16#c0#)) OR
 					(reg_q2124 AND symb_decoder(16#a6#)) OR
 					(reg_q2124 AND symb_decoder(16#f3#)) OR
 					(reg_q2124 AND symb_decoder(16#ac#)) OR
 					(reg_q2124 AND symb_decoder(16#ef#)) OR
 					(reg_q2124 AND symb_decoder(16#a2#)) OR
 					(reg_q2124 AND symb_decoder(16#e9#)) OR
 					(reg_q2124 AND symb_decoder(16#ad#)) OR
 					(reg_q2124 AND symb_decoder(16#3f#)) OR
 					(reg_q2124 AND symb_decoder(16#db#)) OR
 					(reg_q2124 AND symb_decoder(16#90#)) OR
 					(reg_q2124 AND symb_decoder(16#d1#)) OR
 					(reg_q2124 AND symb_decoder(16#80#)) OR
 					(reg_q2124 AND symb_decoder(16#ae#)) OR
 					(reg_q2124 AND symb_decoder(16#26#)) OR
 					(reg_q2124 AND symb_decoder(16#99#)) OR
 					(reg_q2124 AND symb_decoder(16#b2#)) OR
 					(reg_q2124 AND symb_decoder(16#63#)) OR
 					(reg_q2124 AND symb_decoder(16#0b#)) OR
 					(reg_q2124 AND symb_decoder(16#50#)) OR
 					(reg_q2124 AND symb_decoder(16#dd#)) OR
 					(reg_q2124 AND symb_decoder(16#52#)) OR
 					(reg_q2124 AND symb_decoder(16#68#)) OR
 					(reg_q2124 AND symb_decoder(16#08#)) OR
 					(reg_q2124 AND symb_decoder(16#93#)) OR
 					(reg_q2124 AND symb_decoder(16#d7#)) OR
 					(reg_q2124 AND symb_decoder(16#3c#)) OR
 					(reg_q2124 AND symb_decoder(16#3e#)) OR
 					(reg_q2124 AND symb_decoder(16#1f#)) OR
 					(reg_q2124 AND symb_decoder(16#f0#)) OR
 					(reg_q2124 AND symb_decoder(16#da#)) OR
 					(reg_q2124 AND symb_decoder(16#6f#)) OR
 					(reg_q2124 AND symb_decoder(16#8d#)) OR
 					(reg_q2124 AND symb_decoder(16#dc#)) OR
 					(reg_q2124 AND symb_decoder(16#58#)) OR
 					(reg_q2124 AND symb_decoder(16#74#)) OR
 					(reg_q2124 AND symb_decoder(16#10#)) OR
 					(reg_q2124 AND symb_decoder(16#1c#)) OR
 					(reg_q2124 AND symb_decoder(16#45#)) OR
 					(reg_q2124 AND symb_decoder(16#96#)) OR
 					(reg_q2124 AND symb_decoder(16#f9#)) OR
 					(reg_q2124 AND symb_decoder(16#7a#)) OR
 					(reg_q2124 AND symb_decoder(16#a4#)) OR
 					(reg_q2124 AND symb_decoder(16#14#));
reg_q2124_init <= '0' ;
	p_reg_q2124: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2124 <= reg_q2124_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2124 <= reg_q2124_init;
        else
          reg_q2124 <= reg_q2124_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1111_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1111 AND symb_decoder(16#bc#)) OR
 					(reg_q1111 AND symb_decoder(16#0a#)) OR
 					(reg_q1111 AND symb_decoder(16#34#)) OR
 					(reg_q1111 AND symb_decoder(16#a8#)) OR
 					(reg_q1111 AND symb_decoder(16#94#)) OR
 					(reg_q1111 AND symb_decoder(16#ca#)) OR
 					(reg_q1111 AND symb_decoder(16#a6#)) OR
 					(reg_q1111 AND symb_decoder(16#b0#)) OR
 					(reg_q1111 AND symb_decoder(16#f2#)) OR
 					(reg_q1111 AND symb_decoder(16#a1#)) OR
 					(reg_q1111 AND symb_decoder(16#31#)) OR
 					(reg_q1111 AND symb_decoder(16#d9#)) OR
 					(reg_q1111 AND symb_decoder(16#62#)) OR
 					(reg_q1111 AND symb_decoder(16#64#)) OR
 					(reg_q1111 AND symb_decoder(16#fa#)) OR
 					(reg_q1111 AND symb_decoder(16#be#)) OR
 					(reg_q1111 AND symb_decoder(16#76#)) OR
 					(reg_q1111 AND symb_decoder(16#b1#)) OR
 					(reg_q1111 AND symb_decoder(16#29#)) OR
 					(reg_q1111 AND symb_decoder(16#18#)) OR
 					(reg_q1111 AND symb_decoder(16#35#)) OR
 					(reg_q1111 AND symb_decoder(16#1c#)) OR
 					(reg_q1111 AND symb_decoder(16#8f#)) OR
 					(reg_q1111 AND symb_decoder(16#24#)) OR
 					(reg_q1111 AND symb_decoder(16#ff#)) OR
 					(reg_q1111 AND symb_decoder(16#11#)) OR
 					(reg_q1111 AND symb_decoder(16#0e#)) OR
 					(reg_q1111 AND symb_decoder(16#86#)) OR
 					(reg_q1111 AND symb_decoder(16#48#)) OR
 					(reg_q1111 AND symb_decoder(16#aa#)) OR
 					(reg_q1111 AND symb_decoder(16#4d#)) OR
 					(reg_q1111 AND symb_decoder(16#8d#)) OR
 					(reg_q1111 AND symb_decoder(16#d0#)) OR
 					(reg_q1111 AND symb_decoder(16#13#)) OR
 					(reg_q1111 AND symb_decoder(16#97#)) OR
 					(reg_q1111 AND symb_decoder(16#69#)) OR
 					(reg_q1111 AND symb_decoder(16#0c#)) OR
 					(reg_q1111 AND symb_decoder(16#c1#)) OR
 					(reg_q1111 AND symb_decoder(16#c8#)) OR
 					(reg_q1111 AND symb_decoder(16#ae#)) OR
 					(reg_q1111 AND symb_decoder(16#55#)) OR
 					(reg_q1111 AND symb_decoder(16#83#)) OR
 					(reg_q1111 AND symb_decoder(16#3f#)) OR
 					(reg_q1111 AND symb_decoder(16#6c#)) OR
 					(reg_q1111 AND symb_decoder(16#50#)) OR
 					(reg_q1111 AND symb_decoder(16#95#)) OR
 					(reg_q1111 AND symb_decoder(16#1e#)) OR
 					(reg_q1111 AND symb_decoder(16#fc#)) OR
 					(reg_q1111 AND symb_decoder(16#1a#)) OR
 					(reg_q1111 AND symb_decoder(16#5f#)) OR
 					(reg_q1111 AND symb_decoder(16#4b#)) OR
 					(reg_q1111 AND symb_decoder(16#10#)) OR
 					(reg_q1111 AND symb_decoder(16#07#)) OR
 					(reg_q1111 AND symb_decoder(16#f6#)) OR
 					(reg_q1111 AND symb_decoder(16#6f#)) OR
 					(reg_q1111 AND symb_decoder(16#ac#)) OR
 					(reg_q1111 AND symb_decoder(16#dc#)) OR
 					(reg_q1111 AND symb_decoder(16#2f#)) OR
 					(reg_q1111 AND symb_decoder(16#38#)) OR
 					(reg_q1111 AND symb_decoder(16#9d#)) OR
 					(reg_q1111 AND symb_decoder(16#1d#)) OR
 					(reg_q1111 AND symb_decoder(16#6a#)) OR
 					(reg_q1111 AND symb_decoder(16#4c#)) OR
 					(reg_q1111 AND symb_decoder(16#a9#)) OR
 					(reg_q1111 AND symb_decoder(16#db#)) OR
 					(reg_q1111 AND symb_decoder(16#a3#)) OR
 					(reg_q1111 AND symb_decoder(16#3e#)) OR
 					(reg_q1111 AND symb_decoder(16#b6#)) OR
 					(reg_q1111 AND symb_decoder(16#cf#)) OR
 					(reg_q1111 AND symb_decoder(16#5a#)) OR
 					(reg_q1111 AND symb_decoder(16#47#)) OR
 					(reg_q1111 AND symb_decoder(16#fe#)) OR
 					(reg_q1111 AND symb_decoder(16#a4#)) OR
 					(reg_q1111 AND symb_decoder(16#12#)) OR
 					(reg_q1111 AND symb_decoder(16#92#)) OR
 					(reg_q1111 AND symb_decoder(16#ef#)) OR
 					(reg_q1111 AND symb_decoder(16#04#)) OR
 					(reg_q1111 AND symb_decoder(16#59#)) OR
 					(reg_q1111 AND symb_decoder(16#bf#)) OR
 					(reg_q1111 AND symb_decoder(16#3d#)) OR
 					(reg_q1111 AND symb_decoder(16#d6#)) OR
 					(reg_q1111 AND symb_decoder(16#9b#)) OR
 					(reg_q1111 AND symb_decoder(16#21#)) OR
 					(reg_q1111 AND symb_decoder(16#cb#)) OR
 					(reg_q1111 AND symb_decoder(16#14#)) OR
 					(reg_q1111 AND symb_decoder(16#b5#)) OR
 					(reg_q1111 AND symb_decoder(16#e9#)) OR
 					(reg_q1111 AND symb_decoder(16#67#)) OR
 					(reg_q1111 AND symb_decoder(16#20#)) OR
 					(reg_q1111 AND symb_decoder(16#9f#)) OR
 					(reg_q1111 AND symb_decoder(16#c3#)) OR
 					(reg_q1111 AND symb_decoder(16#75#)) OR
 					(reg_q1111 AND symb_decoder(16#c0#)) OR
 					(reg_q1111 AND symb_decoder(16#8e#)) OR
 					(reg_q1111 AND symb_decoder(16#2d#)) OR
 					(reg_q1111 AND symb_decoder(16#80#)) OR
 					(reg_q1111 AND symb_decoder(16#0d#)) OR
 					(reg_q1111 AND symb_decoder(16#da#)) OR
 					(reg_q1111 AND symb_decoder(16#30#)) OR
 					(reg_q1111 AND symb_decoder(16#72#)) OR
 					(reg_q1111 AND symb_decoder(16#7a#)) OR
 					(reg_q1111 AND symb_decoder(16#c2#)) OR
 					(reg_q1111 AND symb_decoder(16#17#)) OR
 					(reg_q1111 AND symb_decoder(16#51#)) OR
 					(reg_q1111 AND symb_decoder(16#43#)) OR
 					(reg_q1111 AND symb_decoder(16#c5#)) OR
 					(reg_q1111 AND symb_decoder(16#16#)) OR
 					(reg_q1111 AND symb_decoder(16#e0#)) OR
 					(reg_q1111 AND symb_decoder(16#5c#)) OR
 					(reg_q1111 AND symb_decoder(16#df#)) OR
 					(reg_q1111 AND symb_decoder(16#b3#)) OR
 					(reg_q1111 AND symb_decoder(16#60#)) OR
 					(reg_q1111 AND symb_decoder(16#28#)) OR
 					(reg_q1111 AND symb_decoder(16#03#)) OR
 					(reg_q1111 AND symb_decoder(16#4f#)) OR
 					(reg_q1111 AND symb_decoder(16#b9#)) OR
 					(reg_q1111 AND symb_decoder(16#57#)) OR
 					(reg_q1111 AND symb_decoder(16#ad#)) OR
 					(reg_q1111 AND symb_decoder(16#6d#)) OR
 					(reg_q1111 AND symb_decoder(16#5e#)) OR
 					(reg_q1111 AND symb_decoder(16#99#)) OR
 					(reg_q1111 AND symb_decoder(16#e6#)) OR
 					(reg_q1111 AND symb_decoder(16#96#)) OR
 					(reg_q1111 AND symb_decoder(16#56#)) OR
 					(reg_q1111 AND symb_decoder(16#f9#)) OR
 					(reg_q1111 AND symb_decoder(16#0f#)) OR
 					(reg_q1111 AND symb_decoder(16#ec#)) OR
 					(reg_q1111 AND symb_decoder(16#73#)) OR
 					(reg_q1111 AND symb_decoder(16#19#)) OR
 					(reg_q1111 AND symb_decoder(16#e8#)) OR
 					(reg_q1111 AND symb_decoder(16#5d#)) OR
 					(reg_q1111 AND symb_decoder(16#7f#)) OR
 					(reg_q1111 AND symb_decoder(16#79#)) OR
 					(reg_q1111 AND symb_decoder(16#84#)) OR
 					(reg_q1111 AND symb_decoder(16#7e#)) OR
 					(reg_q1111 AND symb_decoder(16#c7#)) OR
 					(reg_q1111 AND symb_decoder(16#39#)) OR
 					(reg_q1111 AND symb_decoder(16#41#)) OR
 					(reg_q1111 AND symb_decoder(16#91#)) OR
 					(reg_q1111 AND symb_decoder(16#71#)) OR
 					(reg_q1111 AND symb_decoder(16#6e#)) OR
 					(reg_q1111 AND symb_decoder(16#b4#)) OR
 					(reg_q1111 AND symb_decoder(16#f1#)) OR
 					(reg_q1111 AND symb_decoder(16#78#)) OR
 					(reg_q1111 AND symb_decoder(16#d8#)) OR
 					(reg_q1111 AND symb_decoder(16#40#)) OR
 					(reg_q1111 AND symb_decoder(16#32#)) OR
 					(reg_q1111 AND symb_decoder(16#81#)) OR
 					(reg_q1111 AND symb_decoder(16#d7#)) OR
 					(reg_q1111 AND symb_decoder(16#e1#)) OR
 					(reg_q1111 AND symb_decoder(16#f8#)) OR
 					(reg_q1111 AND symb_decoder(16#eb#)) OR
 					(reg_q1111 AND symb_decoder(16#2b#)) OR
 					(reg_q1111 AND symb_decoder(16#0b#)) OR
 					(reg_q1111 AND symb_decoder(16#2e#)) OR
 					(reg_q1111 AND symb_decoder(16#82#)) OR
 					(reg_q1111 AND symb_decoder(16#9e#)) OR
 					(reg_q1111 AND symb_decoder(16#88#)) OR
 					(reg_q1111 AND symb_decoder(16#89#)) OR
 					(reg_q1111 AND symb_decoder(16#3b#)) OR
 					(reg_q1111 AND symb_decoder(16#d4#)) OR
 					(reg_q1111 AND symb_decoder(16#4a#)) OR
 					(reg_q1111 AND symb_decoder(16#c9#)) OR
 					(reg_q1111 AND symb_decoder(16#74#)) OR
 					(reg_q1111 AND symb_decoder(16#42#)) OR
 					(reg_q1111 AND symb_decoder(16#9a#)) OR
 					(reg_q1111 AND symb_decoder(16#f5#)) OR
 					(reg_q1111 AND symb_decoder(16#ee#)) OR
 					(reg_q1111 AND symb_decoder(16#66#)) OR
 					(reg_q1111 AND symb_decoder(16#37#)) OR
 					(reg_q1111 AND symb_decoder(16#cc#)) OR
 					(reg_q1111 AND symb_decoder(16#d1#)) OR
 					(reg_q1111 AND symb_decoder(16#8a#)) OR
 					(reg_q1111 AND symb_decoder(16#00#)) OR
 					(reg_q1111 AND symb_decoder(16#61#)) OR
 					(reg_q1111 AND symb_decoder(16#70#)) OR
 					(reg_q1111 AND symb_decoder(16#ea#)) OR
 					(reg_q1111 AND symb_decoder(16#7c#)) OR
 					(reg_q1111 AND symb_decoder(16#b8#)) OR
 					(reg_q1111 AND symb_decoder(16#a0#)) OR
 					(reg_q1111 AND symb_decoder(16#bb#)) OR
 					(reg_q1111 AND symb_decoder(16#63#)) OR
 					(reg_q1111 AND symb_decoder(16#45#)) OR
 					(reg_q1111 AND symb_decoder(16#54#)) OR
 					(reg_q1111 AND symb_decoder(16#cd#)) OR
 					(reg_q1111 AND symb_decoder(16#98#)) OR
 					(reg_q1111 AND symb_decoder(16#25#)) OR
 					(reg_q1111 AND symb_decoder(16#49#)) OR
 					(reg_q1111 AND symb_decoder(16#fd#)) OR
 					(reg_q1111 AND symb_decoder(16#e5#)) OR
 					(reg_q1111 AND symb_decoder(16#52#)) OR
 					(reg_q1111 AND symb_decoder(16#36#)) OR
 					(reg_q1111 AND symb_decoder(16#22#)) OR
 					(reg_q1111 AND symb_decoder(16#c4#)) OR
 					(reg_q1111 AND symb_decoder(16#4e#)) OR
 					(reg_q1111 AND symb_decoder(16#c6#)) OR
 					(reg_q1111 AND symb_decoder(16#68#)) OR
 					(reg_q1111 AND symb_decoder(16#05#)) OR
 					(reg_q1111 AND symb_decoder(16#9c#)) OR
 					(reg_q1111 AND symb_decoder(16#e2#)) OR
 					(reg_q1111 AND symb_decoder(16#fb#)) OR
 					(reg_q1111 AND symb_decoder(16#a7#)) OR
 					(reg_q1111 AND symb_decoder(16#2c#)) OR
 					(reg_q1111 AND symb_decoder(16#ed#)) OR
 					(reg_q1111 AND symb_decoder(16#3c#)) OR
 					(reg_q1111 AND symb_decoder(16#e3#)) OR
 					(reg_q1111 AND symb_decoder(16#06#)) OR
 					(reg_q1111 AND symb_decoder(16#dd#)) OR
 					(reg_q1111 AND symb_decoder(16#ab#)) OR
 					(reg_q1111 AND symb_decoder(16#27#)) OR
 					(reg_q1111 AND symb_decoder(16#7b#)) OR
 					(reg_q1111 AND symb_decoder(16#8c#)) OR
 					(reg_q1111 AND symb_decoder(16#6b#)) OR
 					(reg_q1111 AND symb_decoder(16#44#)) OR
 					(reg_q1111 AND symb_decoder(16#ce#)) OR
 					(reg_q1111 AND symb_decoder(16#b7#)) OR
 					(reg_q1111 AND symb_decoder(16#d2#)) OR
 					(reg_q1111 AND symb_decoder(16#f3#)) OR
 					(reg_q1111 AND symb_decoder(16#01#)) OR
 					(reg_q1111 AND symb_decoder(16#f7#)) OR
 					(reg_q1111 AND symb_decoder(16#77#)) OR
 					(reg_q1111 AND symb_decoder(16#2a#)) OR
 					(reg_q1111 AND symb_decoder(16#bd#)) OR
 					(reg_q1111 AND symb_decoder(16#33#)) OR
 					(reg_q1111 AND symb_decoder(16#a2#)) OR
 					(reg_q1111 AND symb_decoder(16#58#)) OR
 					(reg_q1111 AND symb_decoder(16#af#)) OR
 					(reg_q1111 AND symb_decoder(16#8b#)) OR
 					(reg_q1111 AND symb_decoder(16#85#)) OR
 					(reg_q1111 AND symb_decoder(16#d5#)) OR
 					(reg_q1111 AND symb_decoder(16#1b#)) OR
 					(reg_q1111 AND symb_decoder(16#de#)) OR
 					(reg_q1111 AND symb_decoder(16#b2#)) OR
 					(reg_q1111 AND symb_decoder(16#93#)) OR
 					(reg_q1111 AND symb_decoder(16#46#)) OR
 					(reg_q1111 AND symb_decoder(16#f4#)) OR
 					(reg_q1111 AND symb_decoder(16#26#)) OR
 					(reg_q1111 AND symb_decoder(16#7d#)) OR
 					(reg_q1111 AND symb_decoder(16#a5#)) OR
 					(reg_q1111 AND symb_decoder(16#53#)) OR
 					(reg_q1111 AND symb_decoder(16#09#)) OR
 					(reg_q1111 AND symb_decoder(16#e4#)) OR
 					(reg_q1111 AND symb_decoder(16#02#)) OR
 					(reg_q1111 AND symb_decoder(16#5b#)) OR
 					(reg_q1111 AND symb_decoder(16#ba#)) OR
 					(reg_q1111 AND symb_decoder(16#23#)) OR
 					(reg_q1111 AND symb_decoder(16#87#)) OR
 					(reg_q1111 AND symb_decoder(16#08#)) OR
 					(reg_q1111 AND symb_decoder(16#3a#)) OR
 					(reg_q1111 AND symb_decoder(16#90#)) OR
 					(reg_q1111 AND symb_decoder(16#e7#)) OR
 					(reg_q1111 AND symb_decoder(16#1f#)) OR
 					(reg_q1111 AND symb_decoder(16#15#)) OR
 					(reg_q1111 AND symb_decoder(16#f0#)) OR
 					(reg_q1111 AND symb_decoder(16#65#)) OR
 					(reg_q1111 AND symb_decoder(16#d3#));
reg_q1111_init <= '0' ;
	p_reg_q1111: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1111 <= reg_q1111_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1111 <= reg_q1111_init;
        else
          reg_q1111 <= reg_q1111_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q556_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q556 AND symb_decoder(16#a5#)) OR
 					(reg_q556 AND symb_decoder(16#5d#)) OR
 					(reg_q556 AND symb_decoder(16#61#)) OR
 					(reg_q556 AND symb_decoder(16#b8#)) OR
 					(reg_q556 AND symb_decoder(16#98#)) OR
 					(reg_q556 AND symb_decoder(16#65#)) OR
 					(reg_q556 AND symb_decoder(16#3b#)) OR
 					(reg_q556 AND symb_decoder(16#a0#)) OR
 					(reg_q556 AND symb_decoder(16#93#)) OR
 					(reg_q556 AND symb_decoder(16#2d#)) OR
 					(reg_q556 AND symb_decoder(16#8e#)) OR
 					(reg_q556 AND symb_decoder(16#0b#)) OR
 					(reg_q556 AND symb_decoder(16#7d#)) OR
 					(reg_q556 AND symb_decoder(16#7f#)) OR
 					(reg_q556 AND symb_decoder(16#52#)) OR
 					(reg_q556 AND symb_decoder(16#70#)) OR
 					(reg_q556 AND symb_decoder(16#e7#)) OR
 					(reg_q556 AND symb_decoder(16#f9#)) OR
 					(reg_q556 AND symb_decoder(16#62#)) OR
 					(reg_q556 AND symb_decoder(16#92#)) OR
 					(reg_q556 AND symb_decoder(16#53#)) OR
 					(reg_q556 AND symb_decoder(16#74#)) OR
 					(reg_q556 AND symb_decoder(16#c3#)) OR
 					(reg_q556 AND symb_decoder(16#24#)) OR
 					(reg_q556 AND symb_decoder(16#8c#)) OR
 					(reg_q556 AND symb_decoder(16#cb#)) OR
 					(reg_q556 AND symb_decoder(16#71#)) OR
 					(reg_q556 AND symb_decoder(16#1c#)) OR
 					(reg_q556 AND symb_decoder(16#ec#)) OR
 					(reg_q556 AND symb_decoder(16#5f#)) OR
 					(reg_q556 AND symb_decoder(16#73#)) OR
 					(reg_q556 AND symb_decoder(16#ff#)) OR
 					(reg_q556 AND symb_decoder(16#57#)) OR
 					(reg_q556 AND symb_decoder(16#16#)) OR
 					(reg_q556 AND symb_decoder(16#21#)) OR
 					(reg_q556 AND symb_decoder(16#d5#)) OR
 					(reg_q556 AND symb_decoder(16#10#)) OR
 					(reg_q556 AND symb_decoder(16#f5#)) OR
 					(reg_q556 AND symb_decoder(16#bd#)) OR
 					(reg_q556 AND symb_decoder(16#44#)) OR
 					(reg_q556 AND symb_decoder(16#05#)) OR
 					(reg_q556 AND symb_decoder(16#33#)) OR
 					(reg_q556 AND symb_decoder(16#e9#)) OR
 					(reg_q556 AND symb_decoder(16#58#)) OR
 					(reg_q556 AND symb_decoder(16#d1#)) OR
 					(reg_q556 AND symb_decoder(16#72#)) OR
 					(reg_q556 AND symb_decoder(16#30#)) OR
 					(reg_q556 AND symb_decoder(16#c8#)) OR
 					(reg_q556 AND symb_decoder(16#e6#)) OR
 					(reg_q556 AND symb_decoder(16#c4#)) OR
 					(reg_q556 AND symb_decoder(16#f2#)) OR
 					(reg_q556 AND symb_decoder(16#3e#)) OR
 					(reg_q556 AND symb_decoder(16#c2#)) OR
 					(reg_q556 AND symb_decoder(16#d2#)) OR
 					(reg_q556 AND symb_decoder(16#b6#)) OR
 					(reg_q556 AND symb_decoder(16#2b#)) OR
 					(reg_q556 AND symb_decoder(16#6a#)) OR
 					(reg_q556 AND symb_decoder(16#db#)) OR
 					(reg_q556 AND symb_decoder(16#be#)) OR
 					(reg_q556 AND symb_decoder(16#b9#)) OR
 					(reg_q556 AND symb_decoder(16#5a#)) OR
 					(reg_q556 AND symb_decoder(16#4d#)) OR
 					(reg_q556 AND symb_decoder(16#00#)) OR
 					(reg_q556 AND symb_decoder(16#14#)) OR
 					(reg_q556 AND symb_decoder(16#c6#)) OR
 					(reg_q556 AND symb_decoder(16#26#)) OR
 					(reg_q556 AND symb_decoder(16#13#)) OR
 					(reg_q556 AND symb_decoder(16#43#)) OR
 					(reg_q556 AND symb_decoder(16#45#)) OR
 					(reg_q556 AND symb_decoder(16#50#)) OR
 					(reg_q556 AND symb_decoder(16#4c#)) OR
 					(reg_q556 AND symb_decoder(16#49#)) OR
 					(reg_q556 AND symb_decoder(16#a4#)) OR
 					(reg_q556 AND symb_decoder(16#8a#)) OR
 					(reg_q556 AND symb_decoder(16#f4#)) OR
 					(reg_q556 AND symb_decoder(16#66#)) OR
 					(reg_q556 AND symb_decoder(16#1a#)) OR
 					(reg_q556 AND symb_decoder(16#94#)) OR
 					(reg_q556 AND symb_decoder(16#85#)) OR
 					(reg_q556 AND symb_decoder(16#3c#)) OR
 					(reg_q556 AND symb_decoder(16#a9#)) OR
 					(reg_q556 AND symb_decoder(16#38#)) OR
 					(reg_q556 AND symb_decoder(16#42#)) OR
 					(reg_q556 AND symb_decoder(16#84#)) OR
 					(reg_q556 AND symb_decoder(16#3d#)) OR
 					(reg_q556 AND symb_decoder(16#59#)) OR
 					(reg_q556 AND symb_decoder(16#88#)) OR
 					(reg_q556 AND symb_decoder(16#6c#)) OR
 					(reg_q556 AND symb_decoder(16#7c#)) OR
 					(reg_q556 AND symb_decoder(16#fb#)) OR
 					(reg_q556 AND symb_decoder(16#6e#)) OR
 					(reg_q556 AND symb_decoder(16#97#)) OR
 					(reg_q556 AND symb_decoder(16#dc#)) OR
 					(reg_q556 AND symb_decoder(16#32#)) OR
 					(reg_q556 AND symb_decoder(16#40#)) OR
 					(reg_q556 AND symb_decoder(16#5e#)) OR
 					(reg_q556 AND symb_decoder(16#60#)) OR
 					(reg_q556 AND symb_decoder(16#6f#)) OR
 					(reg_q556 AND symb_decoder(16#37#)) OR
 					(reg_q556 AND symb_decoder(16#03#)) OR
 					(reg_q556 AND symb_decoder(16#8f#)) OR
 					(reg_q556 AND symb_decoder(16#99#)) OR
 					(reg_q556 AND symb_decoder(16#f7#)) OR
 					(reg_q556 AND symb_decoder(16#46#)) OR
 					(reg_q556 AND symb_decoder(16#d4#)) OR
 					(reg_q556 AND symb_decoder(16#e0#)) OR
 					(reg_q556 AND symb_decoder(16#04#)) OR
 					(reg_q556 AND symb_decoder(16#81#)) OR
 					(reg_q556 AND symb_decoder(16#82#)) OR
 					(reg_q556 AND symb_decoder(16#f3#)) OR
 					(reg_q556 AND symb_decoder(16#4f#)) OR
 					(reg_q556 AND symb_decoder(16#95#)) OR
 					(reg_q556 AND symb_decoder(16#48#)) OR
 					(reg_q556 AND symb_decoder(16#07#)) OR
 					(reg_q556 AND symb_decoder(16#b0#)) OR
 					(reg_q556 AND symb_decoder(16#a1#)) OR
 					(reg_q556 AND symb_decoder(16#87#)) OR
 					(reg_q556 AND symb_decoder(16#6d#)) OR
 					(reg_q556 AND symb_decoder(16#3a#)) OR
 					(reg_q556 AND symb_decoder(16#bc#)) OR
 					(reg_q556 AND symb_decoder(16#ca#)) OR
 					(reg_q556 AND symb_decoder(16#01#)) OR
 					(reg_q556 AND symb_decoder(16#ae#)) OR
 					(reg_q556 AND symb_decoder(16#da#)) OR
 					(reg_q556 AND symb_decoder(16#f1#)) OR
 					(reg_q556 AND symb_decoder(16#54#)) OR
 					(reg_q556 AND symb_decoder(16#cd#)) OR
 					(reg_q556 AND symb_decoder(16#c0#)) OR
 					(reg_q556 AND symb_decoder(16#c7#)) OR
 					(reg_q556 AND symb_decoder(16#d0#)) OR
 					(reg_q556 AND symb_decoder(16#a2#)) OR
 					(reg_q556 AND symb_decoder(16#2a#)) OR
 					(reg_q556 AND symb_decoder(16#b4#)) OR
 					(reg_q556 AND symb_decoder(16#4e#)) OR
 					(reg_q556 AND symb_decoder(16#7b#)) OR
 					(reg_q556 AND symb_decoder(16#c9#)) OR
 					(reg_q556 AND symb_decoder(16#ac#)) OR
 					(reg_q556 AND symb_decoder(16#5c#)) OR
 					(reg_q556 AND symb_decoder(16#d7#)) OR
 					(reg_q556 AND symb_decoder(16#9e#)) OR
 					(reg_q556 AND symb_decoder(16#4b#)) OR
 					(reg_q556 AND symb_decoder(16#02#)) OR
 					(reg_q556 AND symb_decoder(16#76#)) OR
 					(reg_q556 AND symb_decoder(16#ee#)) OR
 					(reg_q556 AND symb_decoder(16#a7#)) OR
 					(reg_q556 AND symb_decoder(16#78#)) OR
 					(reg_q556 AND symb_decoder(16#0a#)) OR
 					(reg_q556 AND symb_decoder(16#d9#)) OR
 					(reg_q556 AND symb_decoder(16#e3#)) OR
 					(reg_q556 AND symb_decoder(16#ed#)) OR
 					(reg_q556 AND symb_decoder(16#2f#)) OR
 					(reg_q556 AND symb_decoder(16#1d#)) OR
 					(reg_q556 AND symb_decoder(16#39#)) OR
 					(reg_q556 AND symb_decoder(16#51#)) OR
 					(reg_q556 AND symb_decoder(16#31#)) OR
 					(reg_q556 AND symb_decoder(16#2e#)) OR
 					(reg_q556 AND symb_decoder(16#09#)) OR
 					(reg_q556 AND symb_decoder(16#ce#)) OR
 					(reg_q556 AND symb_decoder(16#9d#)) OR
 					(reg_q556 AND symb_decoder(16#41#)) OR
 					(reg_q556 AND symb_decoder(16#b2#)) OR
 					(reg_q556 AND symb_decoder(16#bf#)) OR
 					(reg_q556 AND symb_decoder(16#08#)) OR
 					(reg_q556 AND symb_decoder(16#4a#)) OR
 					(reg_q556 AND symb_decoder(16#fa#)) OR
 					(reg_q556 AND symb_decoder(16#17#)) OR
 					(reg_q556 AND symb_decoder(16#ab#)) OR
 					(reg_q556 AND symb_decoder(16#77#)) OR
 					(reg_q556 AND symb_decoder(16#b5#)) OR
 					(reg_q556 AND symb_decoder(16#a3#)) OR
 					(reg_q556 AND symb_decoder(16#06#)) OR
 					(reg_q556 AND symb_decoder(16#9b#)) OR
 					(reg_q556 AND symb_decoder(16#11#)) OR
 					(reg_q556 AND symb_decoder(16#96#)) OR
 					(reg_q556 AND symb_decoder(16#d3#)) OR
 					(reg_q556 AND symb_decoder(16#fd#)) OR
 					(reg_q556 AND symb_decoder(16#67#)) OR
 					(reg_q556 AND symb_decoder(16#a8#)) OR
 					(reg_q556 AND symb_decoder(16#0d#)) OR
 					(reg_q556 AND symb_decoder(16#b1#)) OR
 					(reg_q556 AND symb_decoder(16#1f#)) OR
 					(reg_q556 AND symb_decoder(16#64#)) OR
 					(reg_q556 AND symb_decoder(16#18#)) OR
 					(reg_q556 AND symb_decoder(16#fe#)) OR
 					(reg_q556 AND symb_decoder(16#f8#)) OR
 					(reg_q556 AND symb_decoder(16#d8#)) OR
 					(reg_q556 AND symb_decoder(16#e2#)) OR
 					(reg_q556 AND symb_decoder(16#2c#)) OR
 					(reg_q556 AND symb_decoder(16#27#)) OR
 					(reg_q556 AND symb_decoder(16#28#)) OR
 					(reg_q556 AND symb_decoder(16#c5#)) OR
 					(reg_q556 AND symb_decoder(16#23#)) OR
 					(reg_q556 AND symb_decoder(16#df#)) OR
 					(reg_q556 AND symb_decoder(16#bb#)) OR
 					(reg_q556 AND symb_decoder(16#a6#)) OR
 					(reg_q556 AND symb_decoder(16#56#)) OR
 					(reg_q556 AND symb_decoder(16#1e#)) OR
 					(reg_q556 AND symb_decoder(16#ba#)) OR
 					(reg_q556 AND symb_decoder(16#d6#)) OR
 					(reg_q556 AND symb_decoder(16#8b#)) OR
 					(reg_q556 AND symb_decoder(16#29#)) OR
 					(reg_q556 AND symb_decoder(16#e8#)) OR
 					(reg_q556 AND symb_decoder(16#22#)) OR
 					(reg_q556 AND symb_decoder(16#0e#)) OR
 					(reg_q556 AND symb_decoder(16#cf#)) OR
 					(reg_q556 AND symb_decoder(16#80#)) OR
 					(reg_q556 AND symb_decoder(16#86#)) OR
 					(reg_q556 AND symb_decoder(16#9f#)) OR
 					(reg_q556 AND symb_decoder(16#cc#)) OR
 					(reg_q556 AND symb_decoder(16#ef#)) OR
 					(reg_q556 AND symb_decoder(16#15#)) OR
 					(reg_q556 AND symb_decoder(16#e4#)) OR
 					(reg_q556 AND symb_decoder(16#55#)) OR
 					(reg_q556 AND symb_decoder(16#12#)) OR
 					(reg_q556 AND symb_decoder(16#f6#)) OR
 					(reg_q556 AND symb_decoder(16#af#)) OR
 					(reg_q556 AND symb_decoder(16#91#)) OR
 					(reg_q556 AND symb_decoder(16#25#)) OR
 					(reg_q556 AND symb_decoder(16#e1#)) OR
 					(reg_q556 AND symb_decoder(16#75#)) OR
 					(reg_q556 AND symb_decoder(16#ea#)) OR
 					(reg_q556 AND symb_decoder(16#3f#)) OR
 					(reg_q556 AND symb_decoder(16#0f#)) OR
 					(reg_q556 AND symb_decoder(16#89#)) OR
 					(reg_q556 AND symb_decoder(16#34#)) OR
 					(reg_q556 AND symb_decoder(16#36#)) OR
 					(reg_q556 AND symb_decoder(16#0c#)) OR
 					(reg_q556 AND symb_decoder(16#20#)) OR
 					(reg_q556 AND symb_decoder(16#e5#)) OR
 					(reg_q556 AND symb_decoder(16#f0#)) OR
 					(reg_q556 AND symb_decoder(16#83#)) OR
 					(reg_q556 AND symb_decoder(16#1b#)) OR
 					(reg_q556 AND symb_decoder(16#7e#)) OR
 					(reg_q556 AND symb_decoder(16#dd#)) OR
 					(reg_q556 AND symb_decoder(16#aa#)) OR
 					(reg_q556 AND symb_decoder(16#47#)) OR
 					(reg_q556 AND symb_decoder(16#9a#)) OR
 					(reg_q556 AND symb_decoder(16#68#)) OR
 					(reg_q556 AND symb_decoder(16#63#)) OR
 					(reg_q556 AND symb_decoder(16#69#)) OR
 					(reg_q556 AND symb_decoder(16#ad#)) OR
 					(reg_q556 AND symb_decoder(16#90#)) OR
 					(reg_q556 AND symb_decoder(16#19#)) OR
 					(reg_q556 AND symb_decoder(16#eb#)) OR
 					(reg_q556 AND symb_decoder(16#b7#)) OR
 					(reg_q556 AND symb_decoder(16#b3#)) OR
 					(reg_q556 AND symb_decoder(16#7a#)) OR
 					(reg_q556 AND symb_decoder(16#de#)) OR
 					(reg_q556 AND symb_decoder(16#35#)) OR
 					(reg_q556 AND symb_decoder(16#79#)) OR
 					(reg_q556 AND symb_decoder(16#9c#)) OR
 					(reg_q556 AND symb_decoder(16#fc#)) OR
 					(reg_q556 AND symb_decoder(16#8d#)) OR
 					(reg_q556 AND symb_decoder(16#c1#)) OR
 					(reg_q556 AND symb_decoder(16#6b#)) OR
 					(reg_q556 AND symb_decoder(16#5b#));
reg_q556_init <= '0' ;
	p_reg_q556: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q556 <= reg_q556_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q556 <= reg_q556_init;
        else
          reg_q556 <= reg_q556_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2091_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2091 AND symb_decoder(16#31#)) OR
 					(reg_q2091 AND symb_decoder(16#2d#)) OR
 					(reg_q2091 AND symb_decoder(16#c3#)) OR
 					(reg_q2091 AND symb_decoder(16#32#)) OR
 					(reg_q2091 AND symb_decoder(16#8c#)) OR
 					(reg_q2091 AND symb_decoder(16#bc#)) OR
 					(reg_q2091 AND symb_decoder(16#9c#)) OR
 					(reg_q2091 AND symb_decoder(16#57#)) OR
 					(reg_q2091 AND symb_decoder(16#4f#)) OR
 					(reg_q2091 AND symb_decoder(16#55#)) OR
 					(reg_q2091 AND symb_decoder(16#18#)) OR
 					(reg_q2091 AND symb_decoder(16#7e#)) OR
 					(reg_q2091 AND symb_decoder(16#ef#)) OR
 					(reg_q2091 AND symb_decoder(16#50#)) OR
 					(reg_q2091 AND symb_decoder(16#2e#)) OR
 					(reg_q2091 AND symb_decoder(16#45#)) OR
 					(reg_q2091 AND symb_decoder(16#3f#)) OR
 					(reg_q2091 AND symb_decoder(16#59#)) OR
 					(reg_q2091 AND symb_decoder(16#a4#)) OR
 					(reg_q2091 AND symb_decoder(16#c4#)) OR
 					(reg_q2091 AND symb_decoder(16#34#)) OR
 					(reg_q2091 AND symb_decoder(16#ff#)) OR
 					(reg_q2091 AND symb_decoder(16#3c#)) OR
 					(reg_q2091 AND symb_decoder(16#fc#)) OR
 					(reg_q2091 AND symb_decoder(16#ce#)) OR
 					(reg_q2091 AND symb_decoder(16#72#)) OR
 					(reg_q2091 AND symb_decoder(16#93#)) OR
 					(reg_q2091 AND symb_decoder(16#26#)) OR
 					(reg_q2091 AND symb_decoder(16#23#)) OR
 					(reg_q2091 AND symb_decoder(16#0a#)) OR
 					(reg_q2091 AND symb_decoder(16#19#)) OR
 					(reg_q2091 AND symb_decoder(16#ca#)) OR
 					(reg_q2091 AND symb_decoder(16#73#)) OR
 					(reg_q2091 AND symb_decoder(16#2b#)) OR
 					(reg_q2091 AND symb_decoder(16#b0#)) OR
 					(reg_q2091 AND symb_decoder(16#07#)) OR
 					(reg_q2091 AND symb_decoder(16#96#)) OR
 					(reg_q2091 AND symb_decoder(16#83#)) OR
 					(reg_q2091 AND symb_decoder(16#38#)) OR
 					(reg_q2091 AND symb_decoder(16#0c#)) OR
 					(reg_q2091 AND symb_decoder(16#43#)) OR
 					(reg_q2091 AND symb_decoder(16#89#)) OR
 					(reg_q2091 AND symb_decoder(16#8d#)) OR
 					(reg_q2091 AND symb_decoder(16#7f#)) OR
 					(reg_q2091 AND symb_decoder(16#7c#)) OR
 					(reg_q2091 AND symb_decoder(16#29#)) OR
 					(reg_q2091 AND symb_decoder(16#2a#)) OR
 					(reg_q2091 AND symb_decoder(16#80#)) OR
 					(reg_q2091 AND symb_decoder(16#d3#)) OR
 					(reg_q2091 AND symb_decoder(16#fd#)) OR
 					(reg_q2091 AND symb_decoder(16#cc#)) OR
 					(reg_q2091 AND symb_decoder(16#81#)) OR
 					(reg_q2091 AND symb_decoder(16#84#)) OR
 					(reg_q2091 AND symb_decoder(16#27#)) OR
 					(reg_q2091 AND symb_decoder(16#a8#)) OR
 					(reg_q2091 AND symb_decoder(16#7b#)) OR
 					(reg_q2091 AND symb_decoder(16#60#)) OR
 					(reg_q2091 AND symb_decoder(16#4c#)) OR
 					(reg_q2091 AND symb_decoder(16#04#)) OR
 					(reg_q2091 AND symb_decoder(16#a1#)) OR
 					(reg_q2091 AND symb_decoder(16#de#)) OR
 					(reg_q2091 AND symb_decoder(16#03#)) OR
 					(reg_q2091 AND symb_decoder(16#5a#)) OR
 					(reg_q2091 AND symb_decoder(16#6a#)) OR
 					(reg_q2091 AND symb_decoder(16#fa#)) OR
 					(reg_q2091 AND symb_decoder(16#f1#)) OR
 					(reg_q2091 AND symb_decoder(16#a0#)) OR
 					(reg_q2091 AND symb_decoder(16#1c#)) OR
 					(reg_q2091 AND symb_decoder(16#ab#)) OR
 					(reg_q2091 AND symb_decoder(16#5f#)) OR
 					(reg_q2091 AND symb_decoder(16#cb#)) OR
 					(reg_q2091 AND symb_decoder(16#24#)) OR
 					(reg_q2091 AND symb_decoder(16#6c#)) OR
 					(reg_q2091 AND symb_decoder(16#e9#)) OR
 					(reg_q2091 AND symb_decoder(16#5c#)) OR
 					(reg_q2091 AND symb_decoder(16#90#)) OR
 					(reg_q2091 AND symb_decoder(16#20#)) OR
 					(reg_q2091 AND symb_decoder(16#16#)) OR
 					(reg_q2091 AND symb_decoder(16#c5#)) OR
 					(reg_q2091 AND symb_decoder(16#c1#)) OR
 					(reg_q2091 AND symb_decoder(16#95#)) OR
 					(reg_q2091 AND symb_decoder(16#13#)) OR
 					(reg_q2091 AND symb_decoder(16#4a#)) OR
 					(reg_q2091 AND symb_decoder(16#98#)) OR
 					(reg_q2091 AND symb_decoder(16#c8#)) OR
 					(reg_q2091 AND symb_decoder(16#d1#)) OR
 					(reg_q2091 AND symb_decoder(16#e4#)) OR
 					(reg_q2091 AND symb_decoder(16#11#)) OR
 					(reg_q2091 AND symb_decoder(16#3b#)) OR
 					(reg_q2091 AND symb_decoder(16#25#)) OR
 					(reg_q2091 AND symb_decoder(16#17#)) OR
 					(reg_q2091 AND symb_decoder(16#d5#)) OR
 					(reg_q2091 AND symb_decoder(16#0f#)) OR
 					(reg_q2091 AND symb_decoder(16#f8#)) OR
 					(reg_q2091 AND symb_decoder(16#c7#)) OR
 					(reg_q2091 AND symb_decoder(16#66#)) OR
 					(reg_q2091 AND symb_decoder(16#1d#)) OR
 					(reg_q2091 AND symb_decoder(16#f7#)) OR
 					(reg_q2091 AND symb_decoder(16#d6#)) OR
 					(reg_q2091 AND symb_decoder(16#68#)) OR
 					(reg_q2091 AND symb_decoder(16#ae#)) OR
 					(reg_q2091 AND symb_decoder(16#85#)) OR
 					(reg_q2091 AND symb_decoder(16#6d#)) OR
 					(reg_q2091 AND symb_decoder(16#65#)) OR
 					(reg_q2091 AND symb_decoder(16#b9#)) OR
 					(reg_q2091 AND symb_decoder(16#5b#)) OR
 					(reg_q2091 AND symb_decoder(16#da#)) OR
 					(reg_q2091 AND symb_decoder(16#1f#)) OR
 					(reg_q2091 AND symb_decoder(16#b2#)) OR
 					(reg_q2091 AND symb_decoder(16#dd#)) OR
 					(reg_q2091 AND symb_decoder(16#b1#)) OR
 					(reg_q2091 AND symb_decoder(16#77#)) OR
 					(reg_q2091 AND symb_decoder(16#f6#)) OR
 					(reg_q2091 AND symb_decoder(16#ad#)) OR
 					(reg_q2091 AND symb_decoder(16#e3#)) OR
 					(reg_q2091 AND symb_decoder(16#00#)) OR
 					(reg_q2091 AND symb_decoder(16#bb#)) OR
 					(reg_q2091 AND symb_decoder(16#02#)) OR
 					(reg_q2091 AND symb_decoder(16#bf#)) OR
 					(reg_q2091 AND symb_decoder(16#06#)) OR
 					(reg_q2091 AND symb_decoder(16#a9#)) OR
 					(reg_q2091 AND symb_decoder(16#67#)) OR
 					(reg_q2091 AND symb_decoder(16#e6#)) OR
 					(reg_q2091 AND symb_decoder(16#c9#)) OR
 					(reg_q2091 AND symb_decoder(16#37#)) OR
 					(reg_q2091 AND symb_decoder(16#05#)) OR
 					(reg_q2091 AND symb_decoder(16#9b#)) OR
 					(reg_q2091 AND symb_decoder(16#ea#)) OR
 					(reg_q2091 AND symb_decoder(16#b4#)) OR
 					(reg_q2091 AND symb_decoder(16#d4#)) OR
 					(reg_q2091 AND symb_decoder(16#5d#)) OR
 					(reg_q2091 AND symb_decoder(16#be#)) OR
 					(reg_q2091 AND symb_decoder(16#61#)) OR
 					(reg_q2091 AND symb_decoder(16#1a#)) OR
 					(reg_q2091 AND symb_decoder(16#6b#)) OR
 					(reg_q2091 AND symb_decoder(16#87#)) OR
 					(reg_q2091 AND symb_decoder(16#44#)) OR
 					(reg_q2091 AND symb_decoder(16#12#)) OR
 					(reg_q2091 AND symb_decoder(16#21#)) OR
 					(reg_q2091 AND symb_decoder(16#a5#)) OR
 					(reg_q2091 AND symb_decoder(16#3a#)) OR
 					(reg_q2091 AND symb_decoder(16#91#)) OR
 					(reg_q2091 AND symb_decoder(16#3e#)) OR
 					(reg_q2091 AND symb_decoder(16#ed#)) OR
 					(reg_q2091 AND symb_decoder(16#46#)) OR
 					(reg_q2091 AND symb_decoder(16#f4#)) OR
 					(reg_q2091 AND symb_decoder(16#dc#)) OR
 					(reg_q2091 AND symb_decoder(16#df#)) OR
 					(reg_q2091 AND symb_decoder(16#47#)) OR
 					(reg_q2091 AND symb_decoder(16#eb#)) OR
 					(reg_q2091 AND symb_decoder(16#0b#)) OR
 					(reg_q2091 AND symb_decoder(16#c6#)) OR
 					(reg_q2091 AND symb_decoder(16#99#)) OR
 					(reg_q2091 AND symb_decoder(16#88#)) OR
 					(reg_q2091 AND symb_decoder(16#71#)) OR
 					(reg_q2091 AND symb_decoder(16#9f#)) OR
 					(reg_q2091 AND symb_decoder(16#78#)) OR
 					(reg_q2091 AND symb_decoder(16#d7#)) OR
 					(reg_q2091 AND symb_decoder(16#af#)) OR
 					(reg_q2091 AND symb_decoder(16#15#)) OR
 					(reg_q2091 AND symb_decoder(16#ba#)) OR
 					(reg_q2091 AND symb_decoder(16#42#)) OR
 					(reg_q2091 AND symb_decoder(16#2f#)) OR
 					(reg_q2091 AND symb_decoder(16#94#)) OR
 					(reg_q2091 AND symb_decoder(16#8b#)) OR
 					(reg_q2091 AND symb_decoder(16#39#)) OR
 					(reg_q2091 AND symb_decoder(16#4b#)) OR
 					(reg_q2091 AND symb_decoder(16#63#)) OR
 					(reg_q2091 AND symb_decoder(16#40#)) OR
 					(reg_q2091 AND symb_decoder(16#e7#)) OR
 					(reg_q2091 AND symb_decoder(16#e1#)) OR
 					(reg_q2091 AND symb_decoder(16#4d#)) OR
 					(reg_q2091 AND symb_decoder(16#30#)) OR
 					(reg_q2091 AND symb_decoder(16#1e#)) OR
 					(reg_q2091 AND symb_decoder(16#56#)) OR
 					(reg_q2091 AND symb_decoder(16#01#)) OR
 					(reg_q2091 AND symb_decoder(16#b6#)) OR
 					(reg_q2091 AND symb_decoder(16#cf#)) OR
 					(reg_q2091 AND symb_decoder(16#53#)) OR
 					(reg_q2091 AND symb_decoder(16#14#)) OR
 					(reg_q2091 AND symb_decoder(16#51#)) OR
 					(reg_q2091 AND symb_decoder(16#f2#)) OR
 					(reg_q2091 AND symb_decoder(16#a2#)) OR
 					(reg_q2091 AND symb_decoder(16#48#)) OR
 					(reg_q2091 AND symb_decoder(16#f0#)) OR
 					(reg_q2091 AND symb_decoder(16#ac#)) OR
 					(reg_q2091 AND symb_decoder(16#f5#)) OR
 					(reg_q2091 AND symb_decoder(16#75#)) OR
 					(reg_q2091 AND symb_decoder(16#9e#)) OR
 					(reg_q2091 AND symb_decoder(16#8e#)) OR
 					(reg_q2091 AND symb_decoder(16#d9#)) OR
 					(reg_q2091 AND symb_decoder(16#a3#)) OR
 					(reg_q2091 AND symb_decoder(16#f9#)) OR
 					(reg_q2091 AND symb_decoder(16#74#)) OR
 					(reg_q2091 AND symb_decoder(16#3d#)) OR
 					(reg_q2091 AND symb_decoder(16#1b#)) OR
 					(reg_q2091 AND symb_decoder(16#6e#)) OR
 					(reg_q2091 AND symb_decoder(16#e8#)) OR
 					(reg_q2091 AND symb_decoder(16#69#)) OR
 					(reg_q2091 AND symb_decoder(16#7d#)) OR
 					(reg_q2091 AND symb_decoder(16#22#)) OR
 					(reg_q2091 AND symb_decoder(16#8f#)) OR
 					(reg_q2091 AND symb_decoder(16#9a#)) OR
 					(reg_q2091 AND symb_decoder(16#9d#)) OR
 					(reg_q2091 AND symb_decoder(16#a7#)) OR
 					(reg_q2091 AND symb_decoder(16#49#)) OR
 					(reg_q2091 AND symb_decoder(16#41#)) OR
 					(reg_q2091 AND symb_decoder(16#4e#)) OR
 					(reg_q2091 AND symb_decoder(16#e5#)) OR
 					(reg_q2091 AND symb_decoder(16#08#)) OR
 					(reg_q2091 AND symb_decoder(16#5e#)) OR
 					(reg_q2091 AND symb_decoder(16#97#)) OR
 					(reg_q2091 AND symb_decoder(16#b7#)) OR
 					(reg_q2091 AND symb_decoder(16#92#)) OR
 					(reg_q2091 AND symb_decoder(16#36#)) OR
 					(reg_q2091 AND symb_decoder(16#82#)) OR
 					(reg_q2091 AND symb_decoder(16#70#)) OR
 					(reg_q2091 AND symb_decoder(16#db#)) OR
 					(reg_q2091 AND symb_decoder(16#79#)) OR
 					(reg_q2091 AND symb_decoder(16#d8#)) OR
 					(reg_q2091 AND symb_decoder(16#d0#)) OR
 					(reg_q2091 AND symb_decoder(16#e0#)) OR
 					(reg_q2091 AND symb_decoder(16#28#)) OR
 					(reg_q2091 AND symb_decoder(16#0e#)) OR
 					(reg_q2091 AND symb_decoder(16#54#)) OR
 					(reg_q2091 AND symb_decoder(16#cd#)) OR
 					(reg_q2091 AND symb_decoder(16#6f#)) OR
 					(reg_q2091 AND symb_decoder(16#2c#)) OR
 					(reg_q2091 AND symb_decoder(16#35#)) OR
 					(reg_q2091 AND symb_decoder(16#64#)) OR
 					(reg_q2091 AND symb_decoder(16#aa#)) OR
 					(reg_q2091 AND symb_decoder(16#fb#)) OR
 					(reg_q2091 AND symb_decoder(16#ee#)) OR
 					(reg_q2091 AND symb_decoder(16#0d#)) OR
 					(reg_q2091 AND symb_decoder(16#09#)) OR
 					(reg_q2091 AND symb_decoder(16#a6#)) OR
 					(reg_q2091 AND symb_decoder(16#e2#)) OR
 					(reg_q2091 AND symb_decoder(16#fe#)) OR
 					(reg_q2091 AND symb_decoder(16#86#)) OR
 					(reg_q2091 AND symb_decoder(16#b3#)) OR
 					(reg_q2091 AND symb_decoder(16#b5#)) OR
 					(reg_q2091 AND symb_decoder(16#62#)) OR
 					(reg_q2091 AND symb_decoder(16#d2#)) OR
 					(reg_q2091 AND symb_decoder(16#33#)) OR
 					(reg_q2091 AND symb_decoder(16#c0#)) OR
 					(reg_q2091 AND symb_decoder(16#8a#)) OR
 					(reg_q2091 AND symb_decoder(16#c2#)) OR
 					(reg_q2091 AND symb_decoder(16#7a#)) OR
 					(reg_q2091 AND symb_decoder(16#bd#)) OR
 					(reg_q2091 AND symb_decoder(16#b8#)) OR
 					(reg_q2091 AND symb_decoder(16#ec#)) OR
 					(reg_q2091 AND symb_decoder(16#58#)) OR
 					(reg_q2091 AND symb_decoder(16#52#)) OR
 					(reg_q2091 AND symb_decoder(16#10#)) OR
 					(reg_q2091 AND symb_decoder(16#f3#)) OR
 					(reg_q2091 AND symb_decoder(16#76#));
reg_q2091_init <= '0' ;
	p_reg_q2091: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2091 <= reg_q2091_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2091 <= reg_q2091_init;
        else
          reg_q2091 <= reg_q2091_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q452_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q452 AND symb_decoder(16#60#)) OR
 					(reg_q452 AND symb_decoder(16#21#)) OR
 					(reg_q452 AND symb_decoder(16#ba#)) OR
 					(reg_q452 AND symb_decoder(16#58#)) OR
 					(reg_q452 AND symb_decoder(16#71#)) OR
 					(reg_q452 AND symb_decoder(16#ec#)) OR
 					(reg_q452 AND symb_decoder(16#c2#)) OR
 					(reg_q452 AND symb_decoder(16#b8#)) OR
 					(reg_q452 AND symb_decoder(16#7d#)) OR
 					(reg_q452 AND symb_decoder(16#6f#)) OR
 					(reg_q452 AND symb_decoder(16#56#)) OR
 					(reg_q452 AND symb_decoder(16#34#)) OR
 					(reg_q452 AND symb_decoder(16#39#)) OR
 					(reg_q452 AND symb_decoder(16#ef#)) OR
 					(reg_q452 AND symb_decoder(16#d2#)) OR
 					(reg_q452 AND symb_decoder(16#66#)) OR
 					(reg_q452 AND symb_decoder(16#16#)) OR
 					(reg_q452 AND symb_decoder(16#f0#)) OR
 					(reg_q452 AND symb_decoder(16#0b#)) OR
 					(reg_q452 AND symb_decoder(16#35#)) OR
 					(reg_q452 AND symb_decoder(16#51#)) OR
 					(reg_q452 AND symb_decoder(16#27#)) OR
 					(reg_q452 AND symb_decoder(16#2c#)) OR
 					(reg_q452 AND symb_decoder(16#e3#)) OR
 					(reg_q452 AND symb_decoder(16#25#)) OR
 					(reg_q452 AND symb_decoder(16#40#)) OR
 					(reg_q452 AND symb_decoder(16#ea#)) OR
 					(reg_q452 AND symb_decoder(16#3b#)) OR
 					(reg_q452 AND symb_decoder(16#7b#)) OR
 					(reg_q452 AND symb_decoder(16#e9#)) OR
 					(reg_q452 AND symb_decoder(16#01#)) OR
 					(reg_q452 AND symb_decoder(16#24#)) OR
 					(reg_q452 AND symb_decoder(16#8e#)) OR
 					(reg_q452 AND symb_decoder(16#a6#)) OR
 					(reg_q452 AND symb_decoder(16#5e#)) OR
 					(reg_q452 AND symb_decoder(16#9f#)) OR
 					(reg_q452 AND symb_decoder(16#c4#)) OR
 					(reg_q452 AND symb_decoder(16#da#)) OR
 					(reg_q452 AND symb_decoder(16#73#)) OR
 					(reg_q452 AND symb_decoder(16#81#)) OR
 					(reg_q452 AND symb_decoder(16#c8#)) OR
 					(reg_q452 AND symb_decoder(16#64#)) OR
 					(reg_q452 AND symb_decoder(16#37#)) OR
 					(reg_q452 AND symb_decoder(16#d1#)) OR
 					(reg_q452 AND symb_decoder(16#50#)) OR
 					(reg_q452 AND symb_decoder(16#7f#)) OR
 					(reg_q452 AND symb_decoder(16#d9#)) OR
 					(reg_q452 AND symb_decoder(16#06#)) OR
 					(reg_q452 AND symb_decoder(16#00#)) OR
 					(reg_q452 AND symb_decoder(16#2d#)) OR
 					(reg_q452 AND symb_decoder(16#85#)) OR
 					(reg_q452 AND symb_decoder(16#8f#)) OR
 					(reg_q452 AND symb_decoder(16#95#)) OR
 					(reg_q452 AND symb_decoder(16#18#)) OR
 					(reg_q452 AND symb_decoder(16#70#)) OR
 					(reg_q452 AND symb_decoder(16#48#)) OR
 					(reg_q452 AND symb_decoder(16#e6#)) OR
 					(reg_q452 AND symb_decoder(16#a8#)) OR
 					(reg_q452 AND symb_decoder(16#3d#)) OR
 					(reg_q452 AND symb_decoder(16#78#)) OR
 					(reg_q452 AND symb_decoder(16#91#)) OR
 					(reg_q452 AND symb_decoder(16#bb#)) OR
 					(reg_q452 AND symb_decoder(16#e0#)) OR
 					(reg_q452 AND symb_decoder(16#db#)) OR
 					(reg_q452 AND symb_decoder(16#44#)) OR
 					(reg_q452 AND symb_decoder(16#92#)) OR
 					(reg_q452 AND symb_decoder(16#46#)) OR
 					(reg_q452 AND symb_decoder(16#f1#)) OR
 					(reg_q452 AND symb_decoder(16#43#)) OR
 					(reg_q452 AND symb_decoder(16#3e#)) OR
 					(reg_q452 AND symb_decoder(16#e8#)) OR
 					(reg_q452 AND symb_decoder(16#ca#)) OR
 					(reg_q452 AND symb_decoder(16#ed#)) OR
 					(reg_q452 AND symb_decoder(16#c6#)) OR
 					(reg_q452 AND symb_decoder(16#9c#)) OR
 					(reg_q452 AND symb_decoder(16#e5#)) OR
 					(reg_q452 AND symb_decoder(16#38#)) OR
 					(reg_q452 AND symb_decoder(16#10#)) OR
 					(reg_q452 AND symb_decoder(16#59#)) OR
 					(reg_q452 AND symb_decoder(16#a1#)) OR
 					(reg_q452 AND symb_decoder(16#82#)) OR
 					(reg_q452 AND symb_decoder(16#a4#)) OR
 					(reg_q452 AND symb_decoder(16#dd#)) OR
 					(reg_q452 AND symb_decoder(16#f3#)) OR
 					(reg_q452 AND symb_decoder(16#f9#)) OR
 					(reg_q452 AND symb_decoder(16#6a#)) OR
 					(reg_q452 AND symb_decoder(16#62#)) OR
 					(reg_q452 AND symb_decoder(16#17#)) OR
 					(reg_q452 AND symb_decoder(16#eb#)) OR
 					(reg_q452 AND symb_decoder(16#b3#)) OR
 					(reg_q452 AND symb_decoder(16#dc#)) OR
 					(reg_q452 AND symb_decoder(16#4e#)) OR
 					(reg_q452 AND symb_decoder(16#5f#)) OR
 					(reg_q452 AND symb_decoder(16#b2#)) OR
 					(reg_q452 AND symb_decoder(16#2b#)) OR
 					(reg_q452 AND symb_decoder(16#cb#)) OR
 					(reg_q452 AND symb_decoder(16#a9#)) OR
 					(reg_q452 AND symb_decoder(16#77#)) OR
 					(reg_q452 AND symb_decoder(16#cd#)) OR
 					(reg_q452 AND symb_decoder(16#54#)) OR
 					(reg_q452 AND symb_decoder(16#a0#)) OR
 					(reg_q452 AND symb_decoder(16#67#)) OR
 					(reg_q452 AND symb_decoder(16#03#)) OR
 					(reg_q452 AND symb_decoder(16#5b#)) OR
 					(reg_q452 AND symb_decoder(16#6d#)) OR
 					(reg_q452 AND symb_decoder(16#e2#)) OR
 					(reg_q452 AND symb_decoder(16#4a#)) OR
 					(reg_q452 AND symb_decoder(16#4d#)) OR
 					(reg_q452 AND symb_decoder(16#bf#)) OR
 					(reg_q452 AND symb_decoder(16#d7#)) OR
 					(reg_q452 AND symb_decoder(16#6b#)) OR
 					(reg_q452 AND symb_decoder(16#ce#)) OR
 					(reg_q452 AND symb_decoder(16#88#)) OR
 					(reg_q452 AND symb_decoder(16#5d#)) OR
 					(reg_q452 AND symb_decoder(16#f8#)) OR
 					(reg_q452 AND symb_decoder(16#26#)) OR
 					(reg_q452 AND symb_decoder(16#53#)) OR
 					(reg_q452 AND symb_decoder(16#76#)) OR
 					(reg_q452 AND symb_decoder(16#fc#)) OR
 					(reg_q452 AND symb_decoder(16#0e#)) OR
 					(reg_q452 AND symb_decoder(16#d0#)) OR
 					(reg_q452 AND symb_decoder(16#45#)) OR
 					(reg_q452 AND symb_decoder(16#d6#)) OR
 					(reg_q452 AND symb_decoder(16#47#)) OR
 					(reg_q452 AND symb_decoder(16#1e#)) OR
 					(reg_q452 AND symb_decoder(16#98#)) OR
 					(reg_q452 AND symb_decoder(16#09#)) OR
 					(reg_q452 AND symb_decoder(16#fa#)) OR
 					(reg_q452 AND symb_decoder(16#20#)) OR
 					(reg_q452 AND symb_decoder(16#b1#)) OR
 					(reg_q452 AND symb_decoder(16#89#)) OR
 					(reg_q452 AND symb_decoder(16#79#)) OR
 					(reg_q452 AND symb_decoder(16#74#)) OR
 					(reg_q452 AND symb_decoder(16#7c#)) OR
 					(reg_q452 AND symb_decoder(16#b4#)) OR
 					(reg_q452 AND symb_decoder(16#29#)) OR
 					(reg_q452 AND symb_decoder(16#c9#)) OR
 					(reg_q452 AND symb_decoder(16#63#)) OR
 					(reg_q452 AND symb_decoder(16#7a#)) OR
 					(reg_q452 AND symb_decoder(16#75#)) OR
 					(reg_q452 AND symb_decoder(16#5a#)) OR
 					(reg_q452 AND symb_decoder(16#52#)) OR
 					(reg_q452 AND symb_decoder(16#ac#)) OR
 					(reg_q452 AND symb_decoder(16#97#)) OR
 					(reg_q452 AND symb_decoder(16#c1#)) OR
 					(reg_q452 AND symb_decoder(16#a7#)) OR
 					(reg_q452 AND symb_decoder(16#3a#)) OR
 					(reg_q452 AND symb_decoder(16#8d#)) OR
 					(reg_q452 AND symb_decoder(16#a3#)) OR
 					(reg_q452 AND symb_decoder(16#2f#)) OR
 					(reg_q452 AND symb_decoder(16#14#)) OR
 					(reg_q452 AND symb_decoder(16#96#)) OR
 					(reg_q452 AND symb_decoder(16#cc#)) OR
 					(reg_q452 AND symb_decoder(16#c0#)) OR
 					(reg_q452 AND symb_decoder(16#d5#)) OR
 					(reg_q452 AND symb_decoder(16#19#)) OR
 					(reg_q452 AND symb_decoder(16#32#)) OR
 					(reg_q452 AND symb_decoder(16#6e#)) OR
 					(reg_q452 AND symb_decoder(16#42#)) OR
 					(reg_q452 AND symb_decoder(16#4c#)) OR
 					(reg_q452 AND symb_decoder(16#0c#)) OR
 					(reg_q452 AND symb_decoder(16#be#)) OR
 					(reg_q452 AND symb_decoder(16#ff#)) OR
 					(reg_q452 AND symb_decoder(16#31#)) OR
 					(reg_q452 AND symb_decoder(16#f6#)) OR
 					(reg_q452 AND symb_decoder(16#61#)) OR
 					(reg_q452 AND symb_decoder(16#f4#)) OR
 					(reg_q452 AND symb_decoder(16#b5#)) OR
 					(reg_q452 AND symb_decoder(16#36#)) OR
 					(reg_q452 AND symb_decoder(16#4f#)) OR
 					(reg_q452 AND symb_decoder(16#1c#)) OR
 					(reg_q452 AND symb_decoder(16#0a#)) OR
 					(reg_q452 AND symb_decoder(16#d8#)) OR
 					(reg_q452 AND symb_decoder(16#8c#)) OR
 					(reg_q452 AND symb_decoder(16#3f#)) OR
 					(reg_q452 AND symb_decoder(16#fb#)) OR
 					(reg_q452 AND symb_decoder(16#57#)) OR
 					(reg_q452 AND symb_decoder(16#80#)) OR
 					(reg_q452 AND symb_decoder(16#b0#)) OR
 					(reg_q452 AND symb_decoder(16#1d#)) OR
 					(reg_q452 AND symb_decoder(16#f2#)) OR
 					(reg_q452 AND symb_decoder(16#02#)) OR
 					(reg_q452 AND symb_decoder(16#84#)) OR
 					(reg_q452 AND symb_decoder(16#fe#)) OR
 					(reg_q452 AND symb_decoder(16#83#)) OR
 					(reg_q452 AND symb_decoder(16#e7#)) OR
 					(reg_q452 AND symb_decoder(16#f7#)) OR
 					(reg_q452 AND symb_decoder(16#68#)) OR
 					(reg_q452 AND symb_decoder(16#ab#)) OR
 					(reg_q452 AND symb_decoder(16#93#)) OR
 					(reg_q452 AND symb_decoder(16#2a#)) OR
 					(reg_q452 AND symb_decoder(16#aa#)) OR
 					(reg_q452 AND symb_decoder(16#23#)) OR
 					(reg_q452 AND symb_decoder(16#04#)) OR
 					(reg_q452 AND symb_decoder(16#99#)) OR
 					(reg_q452 AND symb_decoder(16#28#)) OR
 					(reg_q452 AND symb_decoder(16#41#)) OR
 					(reg_q452 AND symb_decoder(16#bd#)) OR
 					(reg_q452 AND symb_decoder(16#9b#)) OR
 					(reg_q452 AND symb_decoder(16#ee#)) OR
 					(reg_q452 AND symb_decoder(16#94#)) OR
 					(reg_q452 AND symb_decoder(16#0f#)) OR
 					(reg_q452 AND symb_decoder(16#a5#)) OR
 					(reg_q452 AND symb_decoder(16#1f#)) OR
 					(reg_q452 AND symb_decoder(16#90#)) OR
 					(reg_q452 AND symb_decoder(16#c7#)) OR
 					(reg_q452 AND symb_decoder(16#72#)) OR
 					(reg_q452 AND symb_decoder(16#8b#)) OR
 					(reg_q452 AND symb_decoder(16#87#)) OR
 					(reg_q452 AND symb_decoder(16#af#)) OR
 					(reg_q452 AND symb_decoder(16#fd#)) OR
 					(reg_q452 AND symb_decoder(16#de#)) OR
 					(reg_q452 AND symb_decoder(16#5c#)) OR
 					(reg_q452 AND symb_decoder(16#2e#)) OR
 					(reg_q452 AND symb_decoder(16#15#)) OR
 					(reg_q452 AND symb_decoder(16#55#)) OR
 					(reg_q452 AND symb_decoder(16#c5#)) OR
 					(reg_q452 AND symb_decoder(16#9a#)) OR
 					(reg_q452 AND symb_decoder(16#df#)) OR
 					(reg_q452 AND symb_decoder(16#13#)) OR
 					(reg_q452 AND symb_decoder(16#0d#)) OR
 					(reg_q452 AND symb_decoder(16#65#)) OR
 					(reg_q452 AND symb_decoder(16#30#)) OR
 					(reg_q452 AND symb_decoder(16#e4#)) OR
 					(reg_q452 AND symb_decoder(16#cf#)) OR
 					(reg_q452 AND symb_decoder(16#e1#)) OR
 					(reg_q452 AND symb_decoder(16#b6#)) OR
 					(reg_q452 AND symb_decoder(16#7e#)) OR
 					(reg_q452 AND symb_decoder(16#1b#)) OR
 					(reg_q452 AND symb_decoder(16#33#)) OR
 					(reg_q452 AND symb_decoder(16#ae#)) OR
 					(reg_q452 AND symb_decoder(16#4b#)) OR
 					(reg_q452 AND symb_decoder(16#49#)) OR
 					(reg_q452 AND symb_decoder(16#b7#)) OR
 					(reg_q452 AND symb_decoder(16#3c#)) OR
 					(reg_q452 AND symb_decoder(16#69#)) OR
 					(reg_q452 AND symb_decoder(16#9d#)) OR
 					(reg_q452 AND symb_decoder(16#8a#)) OR
 					(reg_q452 AND symb_decoder(16#08#)) OR
 					(reg_q452 AND symb_decoder(16#a2#)) OR
 					(reg_q452 AND symb_decoder(16#22#)) OR
 					(reg_q452 AND symb_decoder(16#9e#)) OR
 					(reg_q452 AND symb_decoder(16#ad#)) OR
 					(reg_q452 AND symb_decoder(16#d3#)) OR
 					(reg_q452 AND symb_decoder(16#86#)) OR
 					(reg_q452 AND symb_decoder(16#bc#)) OR
 					(reg_q452 AND symb_decoder(16#6c#)) OR
 					(reg_q452 AND symb_decoder(16#1a#)) OR
 					(reg_q452 AND symb_decoder(16#07#)) OR
 					(reg_q452 AND symb_decoder(16#d4#)) OR
 					(reg_q452 AND symb_decoder(16#b9#)) OR
 					(reg_q452 AND symb_decoder(16#11#)) OR
 					(reg_q452 AND symb_decoder(16#c3#)) OR
 					(reg_q452 AND symb_decoder(16#f5#)) OR
 					(reg_q452 AND symb_decoder(16#12#)) OR
 					(reg_q452 AND symb_decoder(16#05#));
reg_q452_init <= '0' ;
	p_reg_q452: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q452 <= reg_q452_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q452 <= reg_q452_init;
        else
          reg_q452 <= reg_q452_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1195_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1195 AND symb_decoder(16#e8#)) OR
 					(reg_q1195 AND symb_decoder(16#f5#)) OR
 					(reg_q1195 AND symb_decoder(16#2d#)) OR
 					(reg_q1195 AND symb_decoder(16#d6#)) OR
 					(reg_q1195 AND symb_decoder(16#22#)) OR
 					(reg_q1195 AND symb_decoder(16#82#)) OR
 					(reg_q1195 AND symb_decoder(16#cb#)) OR
 					(reg_q1195 AND symb_decoder(16#fb#)) OR
 					(reg_q1195 AND symb_decoder(16#6d#)) OR
 					(reg_q1195 AND symb_decoder(16#ce#)) OR
 					(reg_q1195 AND symb_decoder(16#7a#)) OR
 					(reg_q1195 AND symb_decoder(16#95#)) OR
 					(reg_q1195 AND symb_decoder(16#93#)) OR
 					(reg_q1195 AND symb_decoder(16#42#)) OR
 					(reg_q1195 AND symb_decoder(16#f6#)) OR
 					(reg_q1195 AND symb_decoder(16#9d#)) OR
 					(reg_q1195 AND symb_decoder(16#04#)) OR
 					(reg_q1195 AND symb_decoder(16#96#)) OR
 					(reg_q1195 AND symb_decoder(16#9c#)) OR
 					(reg_q1195 AND symb_decoder(16#74#)) OR
 					(reg_q1195 AND symb_decoder(16#77#)) OR
 					(reg_q1195 AND symb_decoder(16#53#)) OR
 					(reg_q1195 AND symb_decoder(16#41#)) OR
 					(reg_q1195 AND symb_decoder(16#2a#)) OR
 					(reg_q1195 AND symb_decoder(16#12#)) OR
 					(reg_q1195 AND symb_decoder(16#8c#)) OR
 					(reg_q1195 AND symb_decoder(16#3f#)) OR
 					(reg_q1195 AND symb_decoder(16#aa#)) OR
 					(reg_q1195 AND symb_decoder(16#9f#)) OR
 					(reg_q1195 AND symb_decoder(16#0d#)) OR
 					(reg_q1195 AND symb_decoder(16#ae#)) OR
 					(reg_q1195 AND symb_decoder(16#cd#)) OR
 					(reg_q1195 AND symb_decoder(16#54#)) OR
 					(reg_q1195 AND symb_decoder(16#03#)) OR
 					(reg_q1195 AND symb_decoder(16#8b#)) OR
 					(reg_q1195 AND symb_decoder(16#f4#)) OR
 					(reg_q1195 AND symb_decoder(16#e7#)) OR
 					(reg_q1195 AND symb_decoder(16#e9#)) OR
 					(reg_q1195 AND symb_decoder(16#f2#)) OR
 					(reg_q1195 AND symb_decoder(16#b0#)) OR
 					(reg_q1195 AND symb_decoder(16#d8#)) OR
 					(reg_q1195 AND symb_decoder(16#cf#)) OR
 					(reg_q1195 AND symb_decoder(16#bb#)) OR
 					(reg_q1195 AND symb_decoder(16#36#)) OR
 					(reg_q1195 AND symb_decoder(16#16#)) OR
 					(reg_q1195 AND symb_decoder(16#ff#)) OR
 					(reg_q1195 AND symb_decoder(16#5d#)) OR
 					(reg_q1195 AND symb_decoder(16#ca#)) OR
 					(reg_q1195 AND symb_decoder(16#94#)) OR
 					(reg_q1195 AND symb_decoder(16#2f#)) OR
 					(reg_q1195 AND symb_decoder(16#ba#)) OR
 					(reg_q1195 AND symb_decoder(16#f1#)) OR
 					(reg_q1195 AND symb_decoder(16#df#)) OR
 					(reg_q1195 AND symb_decoder(16#e2#)) OR
 					(reg_q1195 AND symb_decoder(16#01#)) OR
 					(reg_q1195 AND symb_decoder(16#1e#)) OR
 					(reg_q1195 AND symb_decoder(16#17#)) OR
 					(reg_q1195 AND symb_decoder(16#ec#)) OR
 					(reg_q1195 AND symb_decoder(16#50#)) OR
 					(reg_q1195 AND symb_decoder(16#6a#)) OR
 					(reg_q1195 AND symb_decoder(16#a3#)) OR
 					(reg_q1195 AND symb_decoder(16#9b#)) OR
 					(reg_q1195 AND symb_decoder(16#a4#)) OR
 					(reg_q1195 AND symb_decoder(16#90#)) OR
 					(reg_q1195 AND symb_decoder(16#26#)) OR
 					(reg_q1195 AND symb_decoder(16#c1#)) OR
 					(reg_q1195 AND symb_decoder(16#b2#)) OR
 					(reg_q1195 AND symb_decoder(16#c7#)) OR
 					(reg_q1195 AND symb_decoder(16#b5#)) OR
 					(reg_q1195 AND symb_decoder(16#b8#)) OR
 					(reg_q1195 AND symb_decoder(16#97#)) OR
 					(reg_q1195 AND symb_decoder(16#40#)) OR
 					(reg_q1195 AND symb_decoder(16#8f#)) OR
 					(reg_q1195 AND symb_decoder(16#92#)) OR
 					(reg_q1195 AND symb_decoder(16#44#)) OR
 					(reg_q1195 AND symb_decoder(16#ea#)) OR
 					(reg_q1195 AND symb_decoder(16#25#)) OR
 					(reg_q1195 AND symb_decoder(16#05#)) OR
 					(reg_q1195 AND symb_decoder(16#43#)) OR
 					(reg_q1195 AND symb_decoder(16#89#)) OR
 					(reg_q1195 AND symb_decoder(16#98#)) OR
 					(reg_q1195 AND symb_decoder(16#f0#)) OR
 					(reg_q1195 AND symb_decoder(16#11#)) OR
 					(reg_q1195 AND symb_decoder(16#d7#)) OR
 					(reg_q1195 AND symb_decoder(16#87#)) OR
 					(reg_q1195 AND symb_decoder(16#08#)) OR
 					(reg_q1195 AND symb_decoder(16#64#)) OR
 					(reg_q1195 AND symb_decoder(16#88#)) OR
 					(reg_q1195 AND symb_decoder(16#73#)) OR
 					(reg_q1195 AND symb_decoder(16#a5#)) OR
 					(reg_q1195 AND symb_decoder(16#7f#)) OR
 					(reg_q1195 AND symb_decoder(16#5c#)) OR
 					(reg_q1195 AND symb_decoder(16#57#)) OR
 					(reg_q1195 AND symb_decoder(16#62#)) OR
 					(reg_q1195 AND symb_decoder(16#a8#)) OR
 					(reg_q1195 AND symb_decoder(16#3a#)) OR
 					(reg_q1195 AND symb_decoder(16#fc#)) OR
 					(reg_q1195 AND symb_decoder(16#ad#)) OR
 					(reg_q1195 AND symb_decoder(16#55#)) OR
 					(reg_q1195 AND symb_decoder(16#fd#)) OR
 					(reg_q1195 AND symb_decoder(16#58#)) OR
 					(reg_q1195 AND symb_decoder(16#de#)) OR
 					(reg_q1195 AND symb_decoder(16#14#)) OR
 					(reg_q1195 AND symb_decoder(16#46#)) OR
 					(reg_q1195 AND symb_decoder(16#3d#)) OR
 					(reg_q1195 AND symb_decoder(16#eb#)) OR
 					(reg_q1195 AND symb_decoder(16#c3#)) OR
 					(reg_q1195 AND symb_decoder(16#59#)) OR
 					(reg_q1195 AND symb_decoder(16#d3#)) OR
 					(reg_q1195 AND symb_decoder(16#33#)) OR
 					(reg_q1195 AND symb_decoder(16#f7#)) OR
 					(reg_q1195 AND symb_decoder(16#0a#)) OR
 					(reg_q1195 AND symb_decoder(16#06#)) OR
 					(reg_q1195 AND symb_decoder(16#d0#)) OR
 					(reg_q1195 AND symb_decoder(16#28#)) OR
 					(reg_q1195 AND symb_decoder(16#d1#)) OR
 					(reg_q1195 AND symb_decoder(16#02#)) OR
 					(reg_q1195 AND symb_decoder(16#24#)) OR
 					(reg_q1195 AND symb_decoder(16#38#)) OR
 					(reg_q1195 AND symb_decoder(16#5f#)) OR
 					(reg_q1195 AND symb_decoder(16#fa#)) OR
 					(reg_q1195 AND symb_decoder(16#af#)) OR
 					(reg_q1195 AND symb_decoder(16#be#)) OR
 					(reg_q1195 AND symb_decoder(16#e0#)) OR
 					(reg_q1195 AND symb_decoder(16#66#)) OR
 					(reg_q1195 AND symb_decoder(16#f8#)) OR
 					(reg_q1195 AND symb_decoder(16#bf#)) OR
 					(reg_q1195 AND symb_decoder(16#d2#)) OR
 					(reg_q1195 AND symb_decoder(16#c4#)) OR
 					(reg_q1195 AND symb_decoder(16#d9#)) OR
 					(reg_q1195 AND symb_decoder(16#1c#)) OR
 					(reg_q1195 AND symb_decoder(16#ef#)) OR
 					(reg_q1195 AND symb_decoder(16#35#)) OR
 					(reg_q1195 AND symb_decoder(16#e4#)) OR
 					(reg_q1195 AND symb_decoder(16#84#)) OR
 					(reg_q1195 AND symb_decoder(16#dd#)) OR
 					(reg_q1195 AND symb_decoder(16#f3#)) OR
 					(reg_q1195 AND symb_decoder(16#9e#)) OR
 					(reg_q1195 AND symb_decoder(16#45#)) OR
 					(reg_q1195 AND symb_decoder(16#65#)) OR
 					(reg_q1195 AND symb_decoder(16#c0#)) OR
 					(reg_q1195 AND symb_decoder(16#6c#)) OR
 					(reg_q1195 AND symb_decoder(16#cc#)) OR
 					(reg_q1195 AND symb_decoder(16#e6#)) OR
 					(reg_q1195 AND symb_decoder(16#4c#)) OR
 					(reg_q1195 AND symb_decoder(16#0e#)) OR
 					(reg_q1195 AND symb_decoder(16#dc#)) OR
 					(reg_q1195 AND symb_decoder(16#6b#)) OR
 					(reg_q1195 AND symb_decoder(16#7e#)) OR
 					(reg_q1195 AND symb_decoder(16#db#)) OR
 					(reg_q1195 AND symb_decoder(16#70#)) OR
 					(reg_q1195 AND symb_decoder(16#0c#)) OR
 					(reg_q1195 AND symb_decoder(16#d5#)) OR
 					(reg_q1195 AND symb_decoder(16#75#)) OR
 					(reg_q1195 AND symb_decoder(16#52#)) OR
 					(reg_q1195 AND symb_decoder(16#b1#)) OR
 					(reg_q1195 AND symb_decoder(16#1d#)) OR
 					(reg_q1195 AND symb_decoder(16#91#)) OR
 					(reg_q1195 AND symb_decoder(16#1b#)) OR
 					(reg_q1195 AND symb_decoder(16#76#)) OR
 					(reg_q1195 AND symb_decoder(16#47#)) OR
 					(reg_q1195 AND symb_decoder(16#68#)) OR
 					(reg_q1195 AND symb_decoder(16#56#)) OR
 					(reg_q1195 AND symb_decoder(16#c2#)) OR
 					(reg_q1195 AND symb_decoder(16#b6#)) OR
 					(reg_q1195 AND symb_decoder(16#10#)) OR
 					(reg_q1195 AND symb_decoder(16#e1#)) OR
 					(reg_q1195 AND symb_decoder(16#8a#)) OR
 					(reg_q1195 AND symb_decoder(16#2c#)) OR
 					(reg_q1195 AND symb_decoder(16#63#)) OR
 					(reg_q1195 AND symb_decoder(16#09#)) OR
 					(reg_q1195 AND symb_decoder(16#5a#)) OR
 					(reg_q1195 AND symb_decoder(16#18#)) OR
 					(reg_q1195 AND symb_decoder(16#23#)) OR
 					(reg_q1195 AND symb_decoder(16#bc#)) OR
 					(reg_q1195 AND symb_decoder(16#7b#)) OR
 					(reg_q1195 AND symb_decoder(16#99#)) OR
 					(reg_q1195 AND symb_decoder(16#a6#)) OR
 					(reg_q1195 AND symb_decoder(16#48#)) OR
 					(reg_q1195 AND symb_decoder(16#a9#)) OR
 					(reg_q1195 AND symb_decoder(16#80#)) OR
 					(reg_q1195 AND symb_decoder(16#72#)) OR
 					(reg_q1195 AND symb_decoder(16#f9#)) OR
 					(reg_q1195 AND symb_decoder(16#ac#)) OR
 					(reg_q1195 AND symb_decoder(16#27#)) OR
 					(reg_q1195 AND symb_decoder(16#e5#)) OR
 					(reg_q1195 AND symb_decoder(16#19#)) OR
 					(reg_q1195 AND symb_decoder(16#0f#)) OR
 					(reg_q1195 AND symb_decoder(16#20#)) OR
 					(reg_q1195 AND symb_decoder(16#5e#)) OR
 					(reg_q1195 AND symb_decoder(16#c9#)) OR
 					(reg_q1195 AND symb_decoder(16#3b#)) OR
 					(reg_q1195 AND symb_decoder(16#30#)) OR
 					(reg_q1195 AND symb_decoder(16#ee#)) OR
 					(reg_q1195 AND symb_decoder(16#4d#)) OR
 					(reg_q1195 AND symb_decoder(16#c5#)) OR
 					(reg_q1195 AND symb_decoder(16#81#)) OR
 					(reg_q1195 AND symb_decoder(16#3c#)) OR
 					(reg_q1195 AND symb_decoder(16#bd#)) OR
 					(reg_q1195 AND symb_decoder(16#b3#)) OR
 					(reg_q1195 AND symb_decoder(16#b7#)) OR
 					(reg_q1195 AND symb_decoder(16#c8#)) OR
 					(reg_q1195 AND symb_decoder(16#1f#)) OR
 					(reg_q1195 AND symb_decoder(16#3e#)) OR
 					(reg_q1195 AND symb_decoder(16#da#)) OR
 					(reg_q1195 AND symb_decoder(16#ed#)) OR
 					(reg_q1195 AND symb_decoder(16#e3#)) OR
 					(reg_q1195 AND symb_decoder(16#1a#)) OR
 					(reg_q1195 AND symb_decoder(16#ab#)) OR
 					(reg_q1195 AND symb_decoder(16#00#)) OR
 					(reg_q1195 AND symb_decoder(16#6e#)) OR
 					(reg_q1195 AND symb_decoder(16#5b#)) OR
 					(reg_q1195 AND symb_decoder(16#0b#)) OR
 					(reg_q1195 AND symb_decoder(16#69#)) OR
 					(reg_q1195 AND symb_decoder(16#67#)) OR
 					(reg_q1195 AND symb_decoder(16#8e#)) OR
 					(reg_q1195 AND symb_decoder(16#7d#)) OR
 					(reg_q1195 AND symb_decoder(16#9a#)) OR
 					(reg_q1195 AND symb_decoder(16#60#)) OR
 					(reg_q1195 AND symb_decoder(16#b9#)) OR
 					(reg_q1195 AND symb_decoder(16#a7#)) OR
 					(reg_q1195 AND symb_decoder(16#fe#)) OR
 					(reg_q1195 AND symb_decoder(16#51#)) OR
 					(reg_q1195 AND symb_decoder(16#21#)) OR
 					(reg_q1195 AND symb_decoder(16#79#)) OR
 					(reg_q1195 AND symb_decoder(16#c6#)) OR
 					(reg_q1195 AND symb_decoder(16#a2#)) OR
 					(reg_q1195 AND symb_decoder(16#d4#)) OR
 					(reg_q1195 AND symb_decoder(16#37#)) OR
 					(reg_q1195 AND symb_decoder(16#85#)) OR
 					(reg_q1195 AND symb_decoder(16#32#)) OR
 					(reg_q1195 AND symb_decoder(16#78#)) OR
 					(reg_q1195 AND symb_decoder(16#86#)) OR
 					(reg_q1195 AND symb_decoder(16#2e#)) OR
 					(reg_q1195 AND symb_decoder(16#31#)) OR
 					(reg_q1195 AND symb_decoder(16#8d#)) OR
 					(reg_q1195 AND symb_decoder(16#4f#)) OR
 					(reg_q1195 AND symb_decoder(16#4b#)) OR
 					(reg_q1195 AND symb_decoder(16#61#)) OR
 					(reg_q1195 AND symb_decoder(16#2b#)) OR
 					(reg_q1195 AND symb_decoder(16#71#)) OR
 					(reg_q1195 AND symb_decoder(16#b4#)) OR
 					(reg_q1195 AND symb_decoder(16#29#)) OR
 					(reg_q1195 AND symb_decoder(16#a1#)) OR
 					(reg_q1195 AND symb_decoder(16#6f#)) OR
 					(reg_q1195 AND symb_decoder(16#7c#)) OR
 					(reg_q1195 AND symb_decoder(16#a0#)) OR
 					(reg_q1195 AND symb_decoder(16#4e#)) OR
 					(reg_q1195 AND symb_decoder(16#34#)) OR
 					(reg_q1195 AND symb_decoder(16#15#)) OR
 					(reg_q1195 AND symb_decoder(16#13#)) OR
 					(reg_q1195 AND symb_decoder(16#39#)) OR
 					(reg_q1195 AND symb_decoder(16#07#)) OR
 					(reg_q1195 AND symb_decoder(16#4a#)) OR
 					(reg_q1195 AND symb_decoder(16#49#)) OR
 					(reg_q1195 AND symb_decoder(16#83#));
reg_q1195_init <= '0' ;
	p_reg_q1195: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1195 <= reg_q1195_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1195 <= reg_q1195_init;
        else
          reg_q1195 <= reg_q1195_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1644_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1644 AND symb_decoder(16#d6#)) OR
 					(reg_q1644 AND symb_decoder(16#bf#)) OR
 					(reg_q1644 AND symb_decoder(16#43#)) OR
 					(reg_q1644 AND symb_decoder(16#21#)) OR
 					(reg_q1644 AND symb_decoder(16#14#)) OR
 					(reg_q1644 AND symb_decoder(16#e7#)) OR
 					(reg_q1644 AND symb_decoder(16#89#)) OR
 					(reg_q1644 AND symb_decoder(16#0a#)) OR
 					(reg_q1644 AND symb_decoder(16#9e#)) OR
 					(reg_q1644 AND symb_decoder(16#59#)) OR
 					(reg_q1644 AND symb_decoder(16#25#)) OR
 					(reg_q1644 AND symb_decoder(16#2e#)) OR
 					(reg_q1644 AND symb_decoder(16#7e#)) OR
 					(reg_q1644 AND symb_decoder(16#a4#)) OR
 					(reg_q1644 AND symb_decoder(16#4f#)) OR
 					(reg_q1644 AND symb_decoder(16#8a#)) OR
 					(reg_q1644 AND symb_decoder(16#32#)) OR
 					(reg_q1644 AND symb_decoder(16#82#)) OR
 					(reg_q1644 AND symb_decoder(16#02#)) OR
 					(reg_q1644 AND symb_decoder(16#11#)) OR
 					(reg_q1644 AND symb_decoder(16#a7#)) OR
 					(reg_q1644 AND symb_decoder(16#60#)) OR
 					(reg_q1644 AND symb_decoder(16#7d#)) OR
 					(reg_q1644 AND symb_decoder(16#f6#)) OR
 					(reg_q1644 AND symb_decoder(16#91#)) OR
 					(reg_q1644 AND symb_decoder(16#81#)) OR
 					(reg_q1644 AND symb_decoder(16#c2#)) OR
 					(reg_q1644 AND symb_decoder(16#f7#)) OR
 					(reg_q1644 AND symb_decoder(16#52#)) OR
 					(reg_q1644 AND symb_decoder(16#99#)) OR
 					(reg_q1644 AND symb_decoder(16#7c#)) OR
 					(reg_q1644 AND symb_decoder(16#df#)) OR
 					(reg_q1644 AND symb_decoder(16#6e#)) OR
 					(reg_q1644 AND symb_decoder(16#d9#)) OR
 					(reg_q1644 AND symb_decoder(16#c3#)) OR
 					(reg_q1644 AND symb_decoder(16#6b#)) OR
 					(reg_q1644 AND symb_decoder(16#10#)) OR
 					(reg_q1644 AND symb_decoder(16#a9#)) OR
 					(reg_q1644 AND symb_decoder(16#51#)) OR
 					(reg_q1644 AND symb_decoder(16#01#)) OR
 					(reg_q1644 AND symb_decoder(16#57#)) OR
 					(reg_q1644 AND symb_decoder(16#de#)) OR
 					(reg_q1644 AND symb_decoder(16#ac#)) OR
 					(reg_q1644 AND symb_decoder(16#b3#)) OR
 					(reg_q1644 AND symb_decoder(16#d5#)) OR
 					(reg_q1644 AND symb_decoder(16#09#)) OR
 					(reg_q1644 AND symb_decoder(16#9a#)) OR
 					(reg_q1644 AND symb_decoder(16#8c#)) OR
 					(reg_q1644 AND symb_decoder(16#13#)) OR
 					(reg_q1644 AND symb_decoder(16#36#)) OR
 					(reg_q1644 AND symb_decoder(16#1c#)) OR
 					(reg_q1644 AND symb_decoder(16#f4#)) OR
 					(reg_q1644 AND symb_decoder(16#72#)) OR
 					(reg_q1644 AND symb_decoder(16#78#)) OR
 					(reg_q1644 AND symb_decoder(16#b0#)) OR
 					(reg_q1644 AND symb_decoder(16#44#)) OR
 					(reg_q1644 AND symb_decoder(16#c9#)) OR
 					(reg_q1644 AND symb_decoder(16#18#)) OR
 					(reg_q1644 AND symb_decoder(16#41#)) OR
 					(reg_q1644 AND symb_decoder(16#c8#)) OR
 					(reg_q1644 AND symb_decoder(16#9b#)) OR
 					(reg_q1644 AND symb_decoder(16#da#)) OR
 					(reg_q1644 AND symb_decoder(16#46#)) OR
 					(reg_q1644 AND symb_decoder(16#2b#)) OR
 					(reg_q1644 AND symb_decoder(16#48#)) OR
 					(reg_q1644 AND symb_decoder(16#42#)) OR
 					(reg_q1644 AND symb_decoder(16#9c#)) OR
 					(reg_q1644 AND symb_decoder(16#69#)) OR
 					(reg_q1644 AND symb_decoder(16#4d#)) OR
 					(reg_q1644 AND symb_decoder(16#15#)) OR
 					(reg_q1644 AND symb_decoder(16#49#)) OR
 					(reg_q1644 AND symb_decoder(16#d1#)) OR
 					(reg_q1644 AND symb_decoder(16#ef#)) OR
 					(reg_q1644 AND symb_decoder(16#45#)) OR
 					(reg_q1644 AND symb_decoder(16#62#)) OR
 					(reg_q1644 AND symb_decoder(16#06#)) OR
 					(reg_q1644 AND symb_decoder(16#8b#)) OR
 					(reg_q1644 AND symb_decoder(16#95#)) OR
 					(reg_q1644 AND symb_decoder(16#dd#)) OR
 					(reg_q1644 AND symb_decoder(16#7f#)) OR
 					(reg_q1644 AND symb_decoder(16#1d#)) OR
 					(reg_q1644 AND symb_decoder(16#61#)) OR
 					(reg_q1644 AND symb_decoder(16#3f#)) OR
 					(reg_q1644 AND symb_decoder(16#cb#)) OR
 					(reg_q1644 AND symb_decoder(16#56#)) OR
 					(reg_q1644 AND symb_decoder(16#9d#)) OR
 					(reg_q1644 AND symb_decoder(16#d2#)) OR
 					(reg_q1644 AND symb_decoder(16#6f#)) OR
 					(reg_q1644 AND symb_decoder(16#e0#)) OR
 					(reg_q1644 AND symb_decoder(16#22#)) OR
 					(reg_q1644 AND symb_decoder(16#6c#)) OR
 					(reg_q1644 AND symb_decoder(16#79#)) OR
 					(reg_q1644 AND symb_decoder(16#2a#)) OR
 					(reg_q1644 AND symb_decoder(16#bd#)) OR
 					(reg_q1644 AND symb_decoder(16#ae#)) OR
 					(reg_q1644 AND symb_decoder(16#07#)) OR
 					(reg_q1644 AND symb_decoder(16#b2#)) OR
 					(reg_q1644 AND symb_decoder(16#b7#)) OR
 					(reg_q1644 AND symb_decoder(16#b8#)) OR
 					(reg_q1644 AND symb_decoder(16#27#)) OR
 					(reg_q1644 AND symb_decoder(16#e1#)) OR
 					(reg_q1644 AND symb_decoder(16#6a#)) OR
 					(reg_q1644 AND symb_decoder(16#83#)) OR
 					(reg_q1644 AND symb_decoder(16#5f#)) OR
 					(reg_q1644 AND symb_decoder(16#dc#)) OR
 					(reg_q1644 AND symb_decoder(16#e8#)) OR
 					(reg_q1644 AND symb_decoder(16#50#)) OR
 					(reg_q1644 AND symb_decoder(16#2f#)) OR
 					(reg_q1644 AND symb_decoder(16#12#)) OR
 					(reg_q1644 AND symb_decoder(16#e3#)) OR
 					(reg_q1644 AND symb_decoder(16#f1#)) OR
 					(reg_q1644 AND symb_decoder(16#ba#)) OR
 					(reg_q1644 AND symb_decoder(16#93#)) OR
 					(reg_q1644 AND symb_decoder(16#20#)) OR
 					(reg_q1644 AND symb_decoder(16#5d#)) OR
 					(reg_q1644 AND symb_decoder(16#3c#)) OR
 					(reg_q1644 AND symb_decoder(16#ad#)) OR
 					(reg_q1644 AND symb_decoder(16#58#)) OR
 					(reg_q1644 AND symb_decoder(16#b4#)) OR
 					(reg_q1644 AND symb_decoder(16#c4#)) OR
 					(reg_q1644 AND symb_decoder(16#1b#)) OR
 					(reg_q1644 AND symb_decoder(16#a0#)) OR
 					(reg_q1644 AND symb_decoder(16#bc#)) OR
 					(reg_q1644 AND symb_decoder(16#c7#)) OR
 					(reg_q1644 AND symb_decoder(16#38#)) OR
 					(reg_q1644 AND symb_decoder(16#4b#)) OR
 					(reg_q1644 AND symb_decoder(16#fc#)) OR
 					(reg_q1644 AND symb_decoder(16#8f#)) OR
 					(reg_q1644 AND symb_decoder(16#5b#)) OR
 					(reg_q1644 AND symb_decoder(16#64#)) OR
 					(reg_q1644 AND symb_decoder(16#f3#)) OR
 					(reg_q1644 AND symb_decoder(16#c6#)) OR
 					(reg_q1644 AND symb_decoder(16#fe#)) OR
 					(reg_q1644 AND symb_decoder(16#55#)) OR
 					(reg_q1644 AND symb_decoder(16#a8#)) OR
 					(reg_q1644 AND symb_decoder(16#68#)) OR
 					(reg_q1644 AND symb_decoder(16#88#)) OR
 					(reg_q1644 AND symb_decoder(16#a1#)) OR
 					(reg_q1644 AND symb_decoder(16#80#)) OR
 					(reg_q1644 AND symb_decoder(16#b9#)) OR
 					(reg_q1644 AND symb_decoder(16#eb#)) OR
 					(reg_q1644 AND symb_decoder(16#ee#)) OR
 					(reg_q1644 AND symb_decoder(16#53#)) OR
 					(reg_q1644 AND symb_decoder(16#b1#)) OR
 					(reg_q1644 AND symb_decoder(16#24#)) OR
 					(reg_q1644 AND symb_decoder(16#03#)) OR
 					(reg_q1644 AND symb_decoder(16#fa#)) OR
 					(reg_q1644 AND symb_decoder(16#85#)) OR
 					(reg_q1644 AND symb_decoder(16#a6#)) OR
 					(reg_q1644 AND symb_decoder(16#2d#)) OR
 					(reg_q1644 AND symb_decoder(16#90#)) OR
 					(reg_q1644 AND symb_decoder(16#98#)) OR
 					(reg_q1644 AND symb_decoder(16#8d#)) OR
 					(reg_q1644 AND symb_decoder(16#19#)) OR
 					(reg_q1644 AND symb_decoder(16#1f#)) OR
 					(reg_q1644 AND symb_decoder(16#3b#)) OR
 					(reg_q1644 AND symb_decoder(16#87#)) OR
 					(reg_q1644 AND symb_decoder(16#a2#)) OR
 					(reg_q1644 AND symb_decoder(16#9f#)) OR
 					(reg_q1644 AND symb_decoder(16#92#)) OR
 					(reg_q1644 AND symb_decoder(16#cf#)) OR
 					(reg_q1644 AND symb_decoder(16#7a#)) OR
 					(reg_q1644 AND symb_decoder(16#d8#)) OR
 					(reg_q1644 AND symb_decoder(16#ce#)) OR
 					(reg_q1644 AND symb_decoder(16#0e#)) OR
 					(reg_q1644 AND symb_decoder(16#5a#)) OR
 					(reg_q1644 AND symb_decoder(16#35#)) OR
 					(reg_q1644 AND symb_decoder(16#0d#)) OR
 					(reg_q1644 AND symb_decoder(16#3e#)) OR
 					(reg_q1644 AND symb_decoder(16#4a#)) OR
 					(reg_q1644 AND symb_decoder(16#77#)) OR
 					(reg_q1644 AND symb_decoder(16#30#)) OR
 					(reg_q1644 AND symb_decoder(16#ca#)) OR
 					(reg_q1644 AND symb_decoder(16#39#)) OR
 					(reg_q1644 AND symb_decoder(16#ea#)) OR
 					(reg_q1644 AND symb_decoder(16#e2#)) OR
 					(reg_q1644 AND symb_decoder(16#1a#)) OR
 					(reg_q1644 AND symb_decoder(16#ed#)) OR
 					(reg_q1644 AND symb_decoder(16#00#)) OR
 					(reg_q1644 AND symb_decoder(16#d4#)) OR
 					(reg_q1644 AND symb_decoder(16#e4#)) OR
 					(reg_q1644 AND symb_decoder(16#5c#)) OR
 					(reg_q1644 AND symb_decoder(16#17#)) OR
 					(reg_q1644 AND symb_decoder(16#76#)) OR
 					(reg_q1644 AND symb_decoder(16#86#)) OR
 					(reg_q1644 AND symb_decoder(16#bb#)) OR
 					(reg_q1644 AND symb_decoder(16#65#)) OR
 					(reg_q1644 AND symb_decoder(16#cd#)) OR
 					(reg_q1644 AND symb_decoder(16#54#)) OR
 					(reg_q1644 AND symb_decoder(16#63#)) OR
 					(reg_q1644 AND symb_decoder(16#aa#)) OR
 					(reg_q1644 AND symb_decoder(16#37#)) OR
 					(reg_q1644 AND symb_decoder(16#29#)) OR
 					(reg_q1644 AND symb_decoder(16#be#)) OR
 					(reg_q1644 AND symb_decoder(16#4e#)) OR
 					(reg_q1644 AND symb_decoder(16#a5#)) OR
 					(reg_q1644 AND symb_decoder(16#7b#)) OR
 					(reg_q1644 AND symb_decoder(16#f0#)) OR
 					(reg_q1644 AND symb_decoder(16#f8#)) OR
 					(reg_q1644 AND symb_decoder(16#16#)) OR
 					(reg_q1644 AND symb_decoder(16#a3#)) OR
 					(reg_q1644 AND symb_decoder(16#71#)) OR
 					(reg_q1644 AND symb_decoder(16#6d#)) OR
 					(reg_q1644 AND symb_decoder(16#ec#)) OR
 					(reg_q1644 AND symb_decoder(16#3a#)) OR
 					(reg_q1644 AND symb_decoder(16#f5#)) OR
 					(reg_q1644 AND symb_decoder(16#33#)) OR
 					(reg_q1644 AND symb_decoder(16#66#)) OR
 					(reg_q1644 AND symb_decoder(16#97#)) OR
 					(reg_q1644 AND symb_decoder(16#0f#)) OR
 					(reg_q1644 AND symb_decoder(16#94#)) OR
 					(reg_q1644 AND symb_decoder(16#fb#)) OR
 					(reg_q1644 AND symb_decoder(16#5e#)) OR
 					(reg_q1644 AND symb_decoder(16#0c#)) OR
 					(reg_q1644 AND symb_decoder(16#1e#)) OR
 					(reg_q1644 AND symb_decoder(16#e5#)) OR
 					(reg_q1644 AND symb_decoder(16#96#)) OR
 					(reg_q1644 AND symb_decoder(16#ff#)) OR
 					(reg_q1644 AND symb_decoder(16#31#)) OR
 					(reg_q1644 AND symb_decoder(16#f9#)) OR
 					(reg_q1644 AND symb_decoder(16#d7#)) OR
 					(reg_q1644 AND symb_decoder(16#d3#)) OR
 					(reg_q1644 AND symb_decoder(16#fd#)) OR
 					(reg_q1644 AND symb_decoder(16#05#)) OR
 					(reg_q1644 AND symb_decoder(16#e6#)) OR
 					(reg_q1644 AND symb_decoder(16#70#)) OR
 					(reg_q1644 AND symb_decoder(16#08#)) OR
 					(reg_q1644 AND symb_decoder(16#ab#)) OR
 					(reg_q1644 AND symb_decoder(16#0b#)) OR
 					(reg_q1644 AND symb_decoder(16#cc#)) OR
 					(reg_q1644 AND symb_decoder(16#2c#)) OR
 					(reg_q1644 AND symb_decoder(16#47#)) OR
 					(reg_q1644 AND symb_decoder(16#04#)) OR
 					(reg_q1644 AND symb_decoder(16#af#)) OR
 					(reg_q1644 AND symb_decoder(16#73#)) OR
 					(reg_q1644 AND symb_decoder(16#4c#)) OR
 					(reg_q1644 AND symb_decoder(16#8e#)) OR
 					(reg_q1644 AND symb_decoder(16#84#)) OR
 					(reg_q1644 AND symb_decoder(16#f2#)) OR
 					(reg_q1644 AND symb_decoder(16#b5#)) OR
 					(reg_q1644 AND symb_decoder(16#b6#)) OR
 					(reg_q1644 AND symb_decoder(16#e9#)) OR
 					(reg_q1644 AND symb_decoder(16#34#)) OR
 					(reg_q1644 AND symb_decoder(16#c0#)) OR
 					(reg_q1644 AND symb_decoder(16#c1#)) OR
 					(reg_q1644 AND symb_decoder(16#28#)) OR
 					(reg_q1644 AND symb_decoder(16#75#)) OR
 					(reg_q1644 AND symb_decoder(16#23#)) OR
 					(reg_q1644 AND symb_decoder(16#26#)) OR
 					(reg_q1644 AND symb_decoder(16#c5#)) OR
 					(reg_q1644 AND symb_decoder(16#67#)) OR
 					(reg_q1644 AND symb_decoder(16#74#)) OR
 					(reg_q1644 AND symb_decoder(16#40#)) OR
 					(reg_q1644 AND symb_decoder(16#3d#)) OR
 					(reg_q1644 AND symb_decoder(16#d0#)) OR
 					(reg_q1644 AND symb_decoder(16#db#));
reg_q1644_init <= '0' ;
	p_reg_q1644: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1644 <= reg_q1644_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1644 <= reg_q1644_init;
        else
          reg_q1644 <= reg_q1644_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1603_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1603 AND symb_decoder(16#21#)) OR
 					(reg_q1603 AND symb_decoder(16#2a#)) OR
 					(reg_q1603 AND symb_decoder(16#40#)) OR
 					(reg_q1603 AND symb_decoder(16#85#)) OR
 					(reg_q1603 AND symb_decoder(16#47#)) OR
 					(reg_q1603 AND symb_decoder(16#e8#)) OR
 					(reg_q1603 AND symb_decoder(16#84#)) OR
 					(reg_q1603 AND symb_decoder(16#c7#)) OR
 					(reg_q1603 AND symb_decoder(16#b7#)) OR
 					(reg_q1603 AND symb_decoder(16#d5#)) OR
 					(reg_q1603 AND symb_decoder(16#a4#)) OR
 					(reg_q1603 AND symb_decoder(16#be#)) OR
 					(reg_q1603 AND symb_decoder(16#ea#)) OR
 					(reg_q1603 AND symb_decoder(16#27#)) OR
 					(reg_q1603 AND symb_decoder(16#dd#)) OR
 					(reg_q1603 AND symb_decoder(16#13#)) OR
 					(reg_q1603 AND symb_decoder(16#04#)) OR
 					(reg_q1603 AND symb_decoder(16#da#)) OR
 					(reg_q1603 AND symb_decoder(16#16#)) OR
 					(reg_q1603 AND symb_decoder(16#20#)) OR
 					(reg_q1603 AND symb_decoder(16#bf#)) OR
 					(reg_q1603 AND symb_decoder(16#57#)) OR
 					(reg_q1603 AND symb_decoder(16#c9#)) OR
 					(reg_q1603 AND symb_decoder(16#7f#)) OR
 					(reg_q1603 AND symb_decoder(16#9e#)) OR
 					(reg_q1603 AND symb_decoder(16#a0#)) OR
 					(reg_q1603 AND symb_decoder(16#e9#)) OR
 					(reg_q1603 AND symb_decoder(16#58#)) OR
 					(reg_q1603 AND symb_decoder(16#7a#)) OR
 					(reg_q1603 AND symb_decoder(16#de#)) OR
 					(reg_q1603 AND symb_decoder(16#14#)) OR
 					(reg_q1603 AND symb_decoder(16#bd#)) OR
 					(reg_q1603 AND symb_decoder(16#e0#)) OR
 					(reg_q1603 AND symb_decoder(16#4b#)) OR
 					(reg_q1603 AND symb_decoder(16#e1#)) OR
 					(reg_q1603 AND symb_decoder(16#a7#)) OR
 					(reg_q1603 AND symb_decoder(16#fb#)) OR
 					(reg_q1603 AND symb_decoder(16#4f#)) OR
 					(reg_q1603 AND symb_decoder(16#0d#)) OR
 					(reg_q1603 AND symb_decoder(16#ac#)) OR
 					(reg_q1603 AND symb_decoder(16#39#)) OR
 					(reg_q1603 AND symb_decoder(16#7b#)) OR
 					(reg_q1603 AND symb_decoder(16#17#)) OR
 					(reg_q1603 AND symb_decoder(16#5f#)) OR
 					(reg_q1603 AND symb_decoder(16#25#)) OR
 					(reg_q1603 AND symb_decoder(16#09#)) OR
 					(reg_q1603 AND symb_decoder(16#f3#)) OR
 					(reg_q1603 AND symb_decoder(16#ad#)) OR
 					(reg_q1603 AND symb_decoder(16#6f#)) OR
 					(reg_q1603 AND symb_decoder(16#b2#)) OR
 					(reg_q1603 AND symb_decoder(16#ce#)) OR
 					(reg_q1603 AND symb_decoder(16#c5#)) OR
 					(reg_q1603 AND symb_decoder(16#ff#)) OR
 					(reg_q1603 AND symb_decoder(16#44#)) OR
 					(reg_q1603 AND symb_decoder(16#30#)) OR
 					(reg_q1603 AND symb_decoder(16#64#)) OR
 					(reg_q1603 AND symb_decoder(16#1f#)) OR
 					(reg_q1603 AND symb_decoder(16#2c#)) OR
 					(reg_q1603 AND symb_decoder(16#6a#)) OR
 					(reg_q1603 AND symb_decoder(16#a5#)) OR
 					(reg_q1603 AND symb_decoder(16#5c#)) OR
 					(reg_q1603 AND symb_decoder(16#c8#)) OR
 					(reg_q1603 AND symb_decoder(16#ef#)) OR
 					(reg_q1603 AND symb_decoder(16#eb#)) OR
 					(reg_q1603 AND symb_decoder(16#f2#)) OR
 					(reg_q1603 AND symb_decoder(16#1b#)) OR
 					(reg_q1603 AND symb_decoder(16#2d#)) OR
 					(reg_q1603 AND symb_decoder(16#0e#)) OR
 					(reg_q1603 AND symb_decoder(16#f0#)) OR
 					(reg_q1603 AND symb_decoder(16#f6#)) OR
 					(reg_q1603 AND symb_decoder(16#23#)) OR
 					(reg_q1603 AND symb_decoder(16#15#)) OR
 					(reg_q1603 AND symb_decoder(16#33#)) OR
 					(reg_q1603 AND symb_decoder(16#49#)) OR
 					(reg_q1603 AND symb_decoder(16#df#)) OR
 					(reg_q1603 AND symb_decoder(16#8d#)) OR
 					(reg_q1603 AND symb_decoder(16#52#)) OR
 					(reg_q1603 AND symb_decoder(16#9f#)) OR
 					(reg_q1603 AND symb_decoder(16#9a#)) OR
 					(reg_q1603 AND symb_decoder(16#e7#)) OR
 					(reg_q1603 AND symb_decoder(16#73#)) OR
 					(reg_q1603 AND symb_decoder(16#06#)) OR
 					(reg_q1603 AND symb_decoder(16#0a#)) OR
 					(reg_q1603 AND symb_decoder(16#61#)) OR
 					(reg_q1603 AND symb_decoder(16#a6#)) OR
 					(reg_q1603 AND symb_decoder(16#1a#)) OR
 					(reg_q1603 AND symb_decoder(16#1e#)) OR
 					(reg_q1603 AND symb_decoder(16#5d#)) OR
 					(reg_q1603 AND symb_decoder(16#ca#)) OR
 					(reg_q1603 AND symb_decoder(16#91#)) OR
 					(reg_q1603 AND symb_decoder(16#4e#)) OR
 					(reg_q1603 AND symb_decoder(16#f1#)) OR
 					(reg_q1603 AND symb_decoder(16#ec#)) OR
 					(reg_q1603 AND symb_decoder(16#31#)) OR
 					(reg_q1603 AND symb_decoder(16#87#)) OR
 					(reg_q1603 AND symb_decoder(16#c3#)) OR
 					(reg_q1603 AND symb_decoder(16#c6#)) OR
 					(reg_q1603 AND symb_decoder(16#d3#)) OR
 					(reg_q1603 AND symb_decoder(16#7d#)) OR
 					(reg_q1603 AND symb_decoder(16#2b#)) OR
 					(reg_q1603 AND symb_decoder(16#9d#)) OR
 					(reg_q1603 AND symb_decoder(16#83#)) OR
 					(reg_q1603 AND symb_decoder(16#34#)) OR
 					(reg_q1603 AND symb_decoder(16#4c#)) OR
 					(reg_q1603 AND symb_decoder(16#9b#)) OR
 					(reg_q1603 AND symb_decoder(16#89#)) OR
 					(reg_q1603 AND symb_decoder(16#4a#)) OR
 					(reg_q1603 AND symb_decoder(16#bc#)) OR
 					(reg_q1603 AND symb_decoder(16#28#)) OR
 					(reg_q1603 AND symb_decoder(16#69#)) OR
 					(reg_q1603 AND symb_decoder(16#b9#)) OR
 					(reg_q1603 AND symb_decoder(16#29#)) OR
 					(reg_q1603 AND symb_decoder(16#99#)) OR
 					(reg_q1603 AND symb_decoder(16#70#)) OR
 					(reg_q1603 AND symb_decoder(16#8f#)) OR
 					(reg_q1603 AND symb_decoder(16#d4#)) OR
 					(reg_q1603 AND symb_decoder(16#5b#)) OR
 					(reg_q1603 AND symb_decoder(16#10#)) OR
 					(reg_q1603 AND symb_decoder(16#56#)) OR
 					(reg_q1603 AND symb_decoder(16#4d#)) OR
 					(reg_q1603 AND symb_decoder(16#8c#)) OR
 					(reg_q1603 AND symb_decoder(16#0c#)) OR
 					(reg_q1603 AND symb_decoder(16#79#)) OR
 					(reg_q1603 AND symb_decoder(16#07#)) OR
 					(reg_q1603 AND symb_decoder(16#3a#)) OR
 					(reg_q1603 AND symb_decoder(16#82#)) OR
 					(reg_q1603 AND symb_decoder(16#08#)) OR
 					(reg_q1603 AND symb_decoder(16#18#)) OR
 					(reg_q1603 AND symb_decoder(16#8a#)) OR
 					(reg_q1603 AND symb_decoder(16#96#)) OR
 					(reg_q1603 AND symb_decoder(16#af#)) OR
 					(reg_q1603 AND symb_decoder(16#05#)) OR
 					(reg_q1603 AND symb_decoder(16#3d#)) OR
 					(reg_q1603 AND symb_decoder(16#41#)) OR
 					(reg_q1603 AND symb_decoder(16#e3#)) OR
 					(reg_q1603 AND symb_decoder(16#cf#)) OR
 					(reg_q1603 AND symb_decoder(16#b6#)) OR
 					(reg_q1603 AND symb_decoder(16#48#)) OR
 					(reg_q1603 AND symb_decoder(16#2e#)) OR
 					(reg_q1603 AND symb_decoder(16#cc#)) OR
 					(reg_q1603 AND symb_decoder(16#0b#)) OR
 					(reg_q1603 AND symb_decoder(16#dc#)) OR
 					(reg_q1603 AND symb_decoder(16#01#)) OR
 					(reg_q1603 AND symb_decoder(16#d1#)) OR
 					(reg_q1603 AND symb_decoder(16#cb#)) OR
 					(reg_q1603 AND symb_decoder(16#45#)) OR
 					(reg_q1603 AND symb_decoder(16#37#)) OR
 					(reg_q1603 AND symb_decoder(16#00#)) OR
 					(reg_q1603 AND symb_decoder(16#80#)) OR
 					(reg_q1603 AND symb_decoder(16#b5#)) OR
 					(reg_q1603 AND symb_decoder(16#94#)) OR
 					(reg_q1603 AND symb_decoder(16#90#)) OR
 					(reg_q1603 AND symb_decoder(16#db#)) OR
 					(reg_q1603 AND symb_decoder(16#03#)) OR
 					(reg_q1603 AND symb_decoder(16#22#)) OR
 					(reg_q1603 AND symb_decoder(16#e4#)) OR
 					(reg_q1603 AND symb_decoder(16#66#)) OR
 					(reg_q1603 AND symb_decoder(16#36#)) OR
 					(reg_q1603 AND symb_decoder(16#7e#)) OR
 					(reg_q1603 AND symb_decoder(16#32#)) OR
 					(reg_q1603 AND symb_decoder(16#d2#)) OR
 					(reg_q1603 AND symb_decoder(16#b4#)) OR
 					(reg_q1603 AND symb_decoder(16#8e#)) OR
 					(reg_q1603 AND symb_decoder(16#7c#)) OR
 					(reg_q1603 AND symb_decoder(16#e6#)) OR
 					(reg_q1603 AND symb_decoder(16#75#)) OR
 					(reg_q1603 AND symb_decoder(16#ab#)) OR
 					(reg_q1603 AND symb_decoder(16#9c#)) OR
 					(reg_q1603 AND symb_decoder(16#02#)) OR
 					(reg_q1603 AND symb_decoder(16#fa#)) OR
 					(reg_q1603 AND symb_decoder(16#43#)) OR
 					(reg_q1603 AND symb_decoder(16#51#)) OR
 					(reg_q1603 AND symb_decoder(16#e5#)) OR
 					(reg_q1603 AND symb_decoder(16#fc#)) OR
 					(reg_q1603 AND symb_decoder(16#d0#)) OR
 					(reg_q1603 AND symb_decoder(16#86#)) OR
 					(reg_q1603 AND symb_decoder(16#6b#)) OR
 					(reg_q1603 AND symb_decoder(16#d8#)) OR
 					(reg_q1603 AND symb_decoder(16#60#)) OR
 					(reg_q1603 AND symb_decoder(16#c0#)) OR
 					(reg_q1603 AND symb_decoder(16#98#)) OR
 					(reg_q1603 AND symb_decoder(16#1d#)) OR
 					(reg_q1603 AND symb_decoder(16#b8#)) OR
 					(reg_q1603 AND symb_decoder(16#bb#)) OR
 					(reg_q1603 AND symb_decoder(16#f9#)) OR
 					(reg_q1603 AND symb_decoder(16#d7#)) OR
 					(reg_q1603 AND symb_decoder(16#ae#)) OR
 					(reg_q1603 AND symb_decoder(16#68#)) OR
 					(reg_q1603 AND symb_decoder(16#b0#)) OR
 					(reg_q1603 AND symb_decoder(16#74#)) OR
 					(reg_q1603 AND symb_decoder(16#f8#)) OR
 					(reg_q1603 AND symb_decoder(16#38#)) OR
 					(reg_q1603 AND symb_decoder(16#54#)) OR
 					(reg_q1603 AND symb_decoder(16#cd#)) OR
 					(reg_q1603 AND symb_decoder(16#5e#)) OR
 					(reg_q1603 AND symb_decoder(16#6d#)) OR
 					(reg_q1603 AND symb_decoder(16#c4#)) OR
 					(reg_q1603 AND symb_decoder(16#42#)) OR
 					(reg_q1603 AND symb_decoder(16#b3#)) OR
 					(reg_q1603 AND symb_decoder(16#76#)) OR
 					(reg_q1603 AND symb_decoder(16#93#)) OR
 					(reg_q1603 AND symb_decoder(16#c2#)) OR
 					(reg_q1603 AND symb_decoder(16#e2#)) OR
 					(reg_q1603 AND symb_decoder(16#77#)) OR
 					(reg_q1603 AND symb_decoder(16#ed#)) OR
 					(reg_q1603 AND symb_decoder(16#1c#)) OR
 					(reg_q1603 AND symb_decoder(16#88#)) OR
 					(reg_q1603 AND symb_decoder(16#2f#)) OR
 					(reg_q1603 AND symb_decoder(16#97#)) OR
 					(reg_q1603 AND symb_decoder(16#35#)) OR
 					(reg_q1603 AND symb_decoder(16#a3#)) OR
 					(reg_q1603 AND symb_decoder(16#a9#)) OR
 					(reg_q1603 AND symb_decoder(16#6e#)) OR
 					(reg_q1603 AND symb_decoder(16#24#)) OR
 					(reg_q1603 AND symb_decoder(16#95#)) OR
 					(reg_q1603 AND symb_decoder(16#78#)) OR
 					(reg_q1603 AND symb_decoder(16#50#)) OR
 					(reg_q1603 AND symb_decoder(16#65#)) OR
 					(reg_q1603 AND symb_decoder(16#fd#)) OR
 					(reg_q1603 AND symb_decoder(16#a8#)) OR
 					(reg_q1603 AND symb_decoder(16#12#)) OR
 					(reg_q1603 AND symb_decoder(16#f5#)) OR
 					(reg_q1603 AND symb_decoder(16#67#)) OR
 					(reg_q1603 AND symb_decoder(16#92#)) OR
 					(reg_q1603 AND symb_decoder(16#59#)) OR
 					(reg_q1603 AND symb_decoder(16#d6#)) OR
 					(reg_q1603 AND symb_decoder(16#fe#)) OR
 					(reg_q1603 AND symb_decoder(16#3e#)) OR
 					(reg_q1603 AND symb_decoder(16#5a#)) OR
 					(reg_q1603 AND symb_decoder(16#8b#)) OR
 					(reg_q1603 AND symb_decoder(16#ee#)) OR
 					(reg_q1603 AND symb_decoder(16#f4#)) OR
 					(reg_q1603 AND symb_decoder(16#71#)) OR
 					(reg_q1603 AND symb_decoder(16#81#)) OR
 					(reg_q1603 AND symb_decoder(16#d9#)) OR
 					(reg_q1603 AND symb_decoder(16#b1#)) OR
 					(reg_q1603 AND symb_decoder(16#46#)) OR
 					(reg_q1603 AND symb_decoder(16#53#)) OR
 					(reg_q1603 AND symb_decoder(16#f7#)) OR
 					(reg_q1603 AND symb_decoder(16#3f#)) OR
 					(reg_q1603 AND symb_decoder(16#3c#)) OR
 					(reg_q1603 AND symb_decoder(16#ba#)) OR
 					(reg_q1603 AND symb_decoder(16#a2#)) OR
 					(reg_q1603 AND symb_decoder(16#3b#)) OR
 					(reg_q1603 AND symb_decoder(16#72#)) OR
 					(reg_q1603 AND symb_decoder(16#62#)) OR
 					(reg_q1603 AND symb_decoder(16#11#)) OR
 					(reg_q1603 AND symb_decoder(16#aa#)) OR
 					(reg_q1603 AND symb_decoder(16#a1#)) OR
 					(reg_q1603 AND symb_decoder(16#19#)) OR
 					(reg_q1603 AND symb_decoder(16#6c#)) OR
 					(reg_q1603 AND symb_decoder(16#26#)) OR
 					(reg_q1603 AND symb_decoder(16#55#)) OR
 					(reg_q1603 AND symb_decoder(16#63#)) OR
 					(reg_q1603 AND symb_decoder(16#0f#)) OR
 					(reg_q1603 AND symb_decoder(16#c1#));
reg_q1603_init <= '0' ;
	p_reg_q1603: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1603 <= reg_q1603_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1603 <= reg_q1603_init;
        else
          reg_q1603 <= reg_q1603_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2323_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2323 AND symb_decoder(16#64#)) OR
 					(reg_q2323 AND symb_decoder(16#42#)) OR
 					(reg_q2323 AND symb_decoder(16#11#)) OR
 					(reg_q2323 AND symb_decoder(16#b3#)) OR
 					(reg_q2323 AND symb_decoder(16#e0#)) OR
 					(reg_q2323 AND symb_decoder(16#1c#)) OR
 					(reg_q2323 AND symb_decoder(16#f9#)) OR
 					(reg_q2323 AND symb_decoder(16#dd#)) OR
 					(reg_q2323 AND symb_decoder(16#c3#)) OR
 					(reg_q2323 AND symb_decoder(16#26#)) OR
 					(reg_q2323 AND symb_decoder(16#85#)) OR
 					(reg_q2323 AND symb_decoder(16#43#)) OR
 					(reg_q2323 AND symb_decoder(16#c8#)) OR
 					(reg_q2323 AND symb_decoder(16#cd#)) OR
 					(reg_q2323 AND symb_decoder(16#54#)) OR
 					(reg_q2323 AND symb_decoder(16#2a#)) OR
 					(reg_q2323 AND symb_decoder(16#0a#)) OR
 					(reg_q2323 AND symb_decoder(16#37#)) OR
 					(reg_q2323 AND symb_decoder(16#1f#)) OR
 					(reg_q2323 AND symb_decoder(16#92#)) OR
 					(reg_q2323 AND symb_decoder(16#6c#)) OR
 					(reg_q2323 AND symb_decoder(16#59#)) OR
 					(reg_q2323 AND symb_decoder(16#14#)) OR
 					(reg_q2323 AND symb_decoder(16#61#)) OR
 					(reg_q2323 AND symb_decoder(16#b8#)) OR
 					(reg_q2323 AND symb_decoder(16#fe#)) OR
 					(reg_q2323 AND symb_decoder(16#9b#)) OR
 					(reg_q2323 AND symb_decoder(16#41#)) OR
 					(reg_q2323 AND symb_decoder(16#5f#)) OR
 					(reg_q2323 AND symb_decoder(16#58#)) OR
 					(reg_q2323 AND symb_decoder(16#8a#)) OR
 					(reg_q2323 AND symb_decoder(16#d4#)) OR
 					(reg_q2323 AND symb_decoder(16#77#)) OR
 					(reg_q2323 AND symb_decoder(16#06#)) OR
 					(reg_q2323 AND symb_decoder(16#c7#)) OR
 					(reg_q2323 AND symb_decoder(16#ce#)) OR
 					(reg_q2323 AND symb_decoder(16#2b#)) OR
 					(reg_q2323 AND symb_decoder(16#d7#)) OR
 					(reg_q2323 AND symb_decoder(16#4a#)) OR
 					(reg_q2323 AND symb_decoder(16#19#)) OR
 					(reg_q2323 AND symb_decoder(16#25#)) OR
 					(reg_q2323 AND symb_decoder(16#46#)) OR
 					(reg_q2323 AND symb_decoder(16#fd#)) OR
 					(reg_q2323 AND symb_decoder(16#a7#)) OR
 					(reg_q2323 AND symb_decoder(16#3d#)) OR
 					(reg_q2323 AND symb_decoder(16#21#)) OR
 					(reg_q2323 AND symb_decoder(16#97#)) OR
 					(reg_q2323 AND symb_decoder(16#7c#)) OR
 					(reg_q2323 AND symb_decoder(16#d2#)) OR
 					(reg_q2323 AND symb_decoder(16#91#)) OR
 					(reg_q2323 AND symb_decoder(16#af#)) OR
 					(reg_q2323 AND symb_decoder(16#3a#)) OR
 					(reg_q2323 AND symb_decoder(16#4e#)) OR
 					(reg_q2323 AND symb_decoder(16#dc#)) OR
 					(reg_q2323 AND symb_decoder(16#8d#)) OR
 					(reg_q2323 AND symb_decoder(16#94#)) OR
 					(reg_q2323 AND symb_decoder(16#ec#)) OR
 					(reg_q2323 AND symb_decoder(16#ff#)) OR
 					(reg_q2323 AND symb_decoder(16#c4#)) OR
 					(reg_q2323 AND symb_decoder(16#df#)) OR
 					(reg_q2323 AND symb_decoder(16#fa#)) OR
 					(reg_q2323 AND symb_decoder(16#b6#)) OR
 					(reg_q2323 AND symb_decoder(16#52#)) OR
 					(reg_q2323 AND symb_decoder(16#08#)) OR
 					(reg_q2323 AND symb_decoder(16#a4#)) OR
 					(reg_q2323 AND symb_decoder(16#57#)) OR
 					(reg_q2323 AND symb_decoder(16#3e#)) OR
 					(reg_q2323 AND symb_decoder(16#29#)) OR
 					(reg_q2323 AND symb_decoder(16#53#)) OR
 					(reg_q2323 AND symb_decoder(16#eb#)) OR
 					(reg_q2323 AND symb_decoder(16#67#)) OR
 					(reg_q2323 AND symb_decoder(16#cb#)) OR
 					(reg_q2323 AND symb_decoder(16#bf#)) OR
 					(reg_q2323 AND symb_decoder(16#b4#)) OR
 					(reg_q2323 AND symb_decoder(16#02#)) OR
 					(reg_q2323 AND symb_decoder(16#5b#)) OR
 					(reg_q2323 AND symb_decoder(16#b5#)) OR
 					(reg_q2323 AND symb_decoder(16#2d#)) OR
 					(reg_q2323 AND symb_decoder(16#a0#)) OR
 					(reg_q2323 AND symb_decoder(16#56#)) OR
 					(reg_q2323 AND symb_decoder(16#32#)) OR
 					(reg_q2323 AND symb_decoder(16#87#)) OR
 					(reg_q2323 AND symb_decoder(16#89#)) OR
 					(reg_q2323 AND symb_decoder(16#b9#)) OR
 					(reg_q2323 AND symb_decoder(16#51#)) OR
 					(reg_q2323 AND symb_decoder(16#b2#)) OR
 					(reg_q2323 AND symb_decoder(16#db#)) OR
 					(reg_q2323 AND symb_decoder(16#3f#)) OR
 					(reg_q2323 AND symb_decoder(16#7d#)) OR
 					(reg_q2323 AND symb_decoder(16#84#)) OR
 					(reg_q2323 AND symb_decoder(16#ed#)) OR
 					(reg_q2323 AND symb_decoder(16#27#)) OR
 					(reg_q2323 AND symb_decoder(16#98#)) OR
 					(reg_q2323 AND symb_decoder(16#0c#)) OR
 					(reg_q2323 AND symb_decoder(16#01#)) OR
 					(reg_q2323 AND symb_decoder(16#4f#)) OR
 					(reg_q2323 AND symb_decoder(16#3c#)) OR
 					(reg_q2323 AND symb_decoder(16#70#)) OR
 					(reg_q2323 AND symb_decoder(16#f3#)) OR
 					(reg_q2323 AND symb_decoder(16#49#)) OR
 					(reg_q2323 AND symb_decoder(16#0b#)) OR
 					(reg_q2323 AND symb_decoder(16#b1#)) OR
 					(reg_q2323 AND symb_decoder(16#d3#)) OR
 					(reg_q2323 AND symb_decoder(16#71#)) OR
 					(reg_q2323 AND symb_decoder(16#13#)) OR
 					(reg_q2323 AND symb_decoder(16#16#)) OR
 					(reg_q2323 AND symb_decoder(16#7a#)) OR
 					(reg_q2323 AND symb_decoder(16#4d#)) OR
 					(reg_q2323 AND symb_decoder(16#6d#)) OR
 					(reg_q2323 AND symb_decoder(16#6f#)) OR
 					(reg_q2323 AND symb_decoder(16#a6#)) OR
 					(reg_q2323 AND symb_decoder(16#31#)) OR
 					(reg_q2323 AND symb_decoder(16#44#)) OR
 					(reg_q2323 AND symb_decoder(16#45#)) OR
 					(reg_q2323 AND symb_decoder(16#cc#)) OR
 					(reg_q2323 AND symb_decoder(16#82#)) OR
 					(reg_q2323 AND symb_decoder(16#e7#)) OR
 					(reg_q2323 AND symb_decoder(16#ef#)) OR
 					(reg_q2323 AND symb_decoder(16#99#)) OR
 					(reg_q2323 AND symb_decoder(16#88#)) OR
 					(reg_q2323 AND symb_decoder(16#9e#)) OR
 					(reg_q2323 AND symb_decoder(16#e2#)) OR
 					(reg_q2323 AND symb_decoder(16#7b#)) OR
 					(reg_q2323 AND symb_decoder(16#8c#)) OR
 					(reg_q2323 AND symb_decoder(16#80#)) OR
 					(reg_q2323 AND symb_decoder(16#5e#)) OR
 					(reg_q2323 AND symb_decoder(16#d0#)) OR
 					(reg_q2323 AND symb_decoder(16#6b#)) OR
 					(reg_q2323 AND symb_decoder(16#39#)) OR
 					(reg_q2323 AND symb_decoder(16#6e#)) OR
 					(reg_q2323 AND symb_decoder(16#e6#)) OR
 					(reg_q2323 AND symb_decoder(16#5c#)) OR
 					(reg_q2323 AND symb_decoder(16#6a#)) OR
 					(reg_q2323 AND symb_decoder(16#18#)) OR
 					(reg_q2323 AND symb_decoder(16#c2#)) OR
 					(reg_q2323 AND symb_decoder(16#8e#)) OR
 					(reg_q2323 AND symb_decoder(16#c5#)) OR
 					(reg_q2323 AND symb_decoder(16#93#)) OR
 					(reg_q2323 AND symb_decoder(16#48#)) OR
 					(reg_q2323 AND symb_decoder(16#78#)) OR
 					(reg_q2323 AND symb_decoder(16#09#)) OR
 					(reg_q2323 AND symb_decoder(16#9c#)) OR
 					(reg_q2323 AND symb_decoder(16#04#)) OR
 					(reg_q2323 AND symb_decoder(16#a2#)) OR
 					(reg_q2323 AND symb_decoder(16#62#)) OR
 					(reg_q2323 AND symb_decoder(16#90#)) OR
 					(reg_q2323 AND symb_decoder(16#b0#)) OR
 					(reg_q2323 AND symb_decoder(16#5a#)) OR
 					(reg_q2323 AND symb_decoder(16#22#)) OR
 					(reg_q2323 AND symb_decoder(16#05#)) OR
 					(reg_q2323 AND symb_decoder(16#24#)) OR
 					(reg_q2323 AND symb_decoder(16#aa#)) OR
 					(reg_q2323 AND symb_decoder(16#1b#)) OR
 					(reg_q2323 AND symb_decoder(16#60#)) OR
 					(reg_q2323 AND symb_decoder(16#79#)) OR
 					(reg_q2323 AND symb_decoder(16#b7#)) OR
 					(reg_q2323 AND symb_decoder(16#d6#)) OR
 					(reg_q2323 AND symb_decoder(16#9d#)) OR
 					(reg_q2323 AND symb_decoder(16#e4#)) OR
 					(reg_q2323 AND symb_decoder(16#ca#)) OR
 					(reg_q2323 AND symb_decoder(16#30#)) OR
 					(reg_q2323 AND symb_decoder(16#1a#)) OR
 					(reg_q2323 AND symb_decoder(16#33#)) OR
 					(reg_q2323 AND symb_decoder(16#2e#)) OR
 					(reg_q2323 AND symb_decoder(16#c6#)) OR
 					(reg_q2323 AND symb_decoder(16#1d#)) OR
 					(reg_q2323 AND symb_decoder(16#d5#)) OR
 					(reg_q2323 AND symb_decoder(16#bd#)) OR
 					(reg_q2323 AND symb_decoder(16#95#)) OR
 					(reg_q2323 AND symb_decoder(16#96#)) OR
 					(reg_q2323 AND symb_decoder(16#d1#)) OR
 					(reg_q2323 AND symb_decoder(16#c1#)) OR
 					(reg_q2323 AND symb_decoder(16#15#)) OR
 					(reg_q2323 AND symb_decoder(16#8b#)) OR
 					(reg_q2323 AND symb_decoder(16#23#)) OR
 					(reg_q2323 AND symb_decoder(16#4c#)) OR
 					(reg_q2323 AND symb_decoder(16#f6#)) OR
 					(reg_q2323 AND symb_decoder(16#50#)) OR
 					(reg_q2323 AND symb_decoder(16#c9#)) OR
 					(reg_q2323 AND symb_decoder(16#ea#)) OR
 					(reg_q2323 AND symb_decoder(16#7f#)) OR
 					(reg_q2323 AND symb_decoder(16#a9#)) OR
 					(reg_q2323 AND symb_decoder(16#68#)) OR
 					(reg_q2323 AND symb_decoder(16#a8#)) OR
 					(reg_q2323 AND symb_decoder(16#63#)) OR
 					(reg_q2323 AND symb_decoder(16#d8#)) OR
 					(reg_q2323 AND symb_decoder(16#0e#)) OR
 					(reg_q2323 AND symb_decoder(16#36#)) OR
 					(reg_q2323 AND symb_decoder(16#47#)) OR
 					(reg_q2323 AND symb_decoder(16#e9#)) OR
 					(reg_q2323 AND symb_decoder(16#72#)) OR
 					(reg_q2323 AND symb_decoder(16#ad#)) OR
 					(reg_q2323 AND symb_decoder(16#bb#)) OR
 					(reg_q2323 AND symb_decoder(16#ae#)) OR
 					(reg_q2323 AND symb_decoder(16#bc#)) OR
 					(reg_q2323 AND symb_decoder(16#73#)) OR
 					(reg_q2323 AND symb_decoder(16#fb#)) OR
 					(reg_q2323 AND symb_decoder(16#ee#)) OR
 					(reg_q2323 AND symb_decoder(16#03#)) OR
 					(reg_q2323 AND symb_decoder(16#40#)) OR
 					(reg_q2323 AND symb_decoder(16#ac#)) OR
 					(reg_q2323 AND symb_decoder(16#10#)) OR
 					(reg_q2323 AND symb_decoder(16#0d#)) OR
 					(reg_q2323 AND symb_decoder(16#1e#)) OR
 					(reg_q2323 AND symb_decoder(16#74#)) OR
 					(reg_q2323 AND symb_decoder(16#ab#)) OR
 					(reg_q2323 AND symb_decoder(16#9a#)) OR
 					(reg_q2323 AND symb_decoder(16#7e#)) OR
 					(reg_q2323 AND symb_decoder(16#4b#)) OR
 					(reg_q2323 AND symb_decoder(16#83#)) OR
 					(reg_q2323 AND symb_decoder(16#f4#)) OR
 					(reg_q2323 AND symb_decoder(16#07#)) OR
 					(reg_q2323 AND symb_decoder(16#2c#)) OR
 					(reg_q2323 AND symb_decoder(16#34#)) OR
 					(reg_q2323 AND symb_decoder(16#55#)) OR
 					(reg_q2323 AND symb_decoder(16#fc#)) OR
 					(reg_q2323 AND symb_decoder(16#35#)) OR
 					(reg_q2323 AND symb_decoder(16#e5#)) OR
 					(reg_q2323 AND symb_decoder(16#f1#)) OR
 					(reg_q2323 AND symb_decoder(16#a3#)) OR
 					(reg_q2323 AND symb_decoder(16#2f#)) OR
 					(reg_q2323 AND symb_decoder(16#00#)) OR
 					(reg_q2323 AND symb_decoder(16#f5#)) OR
 					(reg_q2323 AND symb_decoder(16#c0#)) OR
 					(reg_q2323 AND symb_decoder(16#f8#)) OR
 					(reg_q2323 AND symb_decoder(16#e3#)) OR
 					(reg_q2323 AND symb_decoder(16#f0#)) OR
 					(reg_q2323 AND symb_decoder(16#76#)) OR
 					(reg_q2323 AND symb_decoder(16#3b#)) OR
 					(reg_q2323 AND symb_decoder(16#20#)) OR
 					(reg_q2323 AND symb_decoder(16#28#)) OR
 					(reg_q2323 AND symb_decoder(16#a5#)) OR
 					(reg_q2323 AND symb_decoder(16#be#)) OR
 					(reg_q2323 AND symb_decoder(16#da#)) OR
 					(reg_q2323 AND symb_decoder(16#5d#)) OR
 					(reg_q2323 AND symb_decoder(16#cf#)) OR
 					(reg_q2323 AND symb_decoder(16#75#)) OR
 					(reg_q2323 AND symb_decoder(16#d9#)) OR
 					(reg_q2323 AND symb_decoder(16#de#)) OR
 					(reg_q2323 AND symb_decoder(16#e8#)) OR
 					(reg_q2323 AND symb_decoder(16#ba#)) OR
 					(reg_q2323 AND symb_decoder(16#69#)) OR
 					(reg_q2323 AND symb_decoder(16#9f#)) OR
 					(reg_q2323 AND symb_decoder(16#a1#)) OR
 					(reg_q2323 AND symb_decoder(16#e1#)) OR
 					(reg_q2323 AND symb_decoder(16#12#)) OR
 					(reg_q2323 AND symb_decoder(16#65#)) OR
 					(reg_q2323 AND symb_decoder(16#38#)) OR
 					(reg_q2323 AND symb_decoder(16#86#)) OR
 					(reg_q2323 AND symb_decoder(16#f7#)) OR
 					(reg_q2323 AND symb_decoder(16#81#)) OR
 					(reg_q2323 AND symb_decoder(16#8f#)) OR
 					(reg_q2323 AND symb_decoder(16#66#)) OR
 					(reg_q2323 AND symb_decoder(16#0f#)) OR
 					(reg_q2323 AND symb_decoder(16#17#)) OR
 					(reg_q2323 AND symb_decoder(16#f2#));
reg_q2323_init <= '0' ;
	p_reg_q2323: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2323 <= reg_q2323_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2323 <= reg_q2323_init;
        else
          reg_q2323 <= reg_q2323_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1013_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1013 AND symb_decoder(16#6f#)) OR
 					(reg_q1013 AND symb_decoder(16#eb#)) OR
 					(reg_q1013 AND symb_decoder(16#b4#)) OR
 					(reg_q1013 AND symb_decoder(16#36#)) OR
 					(reg_q1013 AND symb_decoder(16#37#)) OR
 					(reg_q1013 AND symb_decoder(16#7f#)) OR
 					(reg_q1013 AND symb_decoder(16#26#)) OR
 					(reg_q1013 AND symb_decoder(16#53#)) OR
 					(reg_q1013 AND symb_decoder(16#d9#)) OR
 					(reg_q1013 AND symb_decoder(16#e4#)) OR
 					(reg_q1013 AND symb_decoder(16#f8#)) OR
 					(reg_q1013 AND symb_decoder(16#d3#)) OR
 					(reg_q1013 AND symb_decoder(16#1d#)) OR
 					(reg_q1013 AND symb_decoder(16#7d#)) OR
 					(reg_q1013 AND symb_decoder(16#f5#)) OR
 					(reg_q1013 AND symb_decoder(16#1c#)) OR
 					(reg_q1013 AND symb_decoder(16#8b#)) OR
 					(reg_q1013 AND symb_decoder(16#44#)) OR
 					(reg_q1013 AND symb_decoder(16#8a#)) OR
 					(reg_q1013 AND symb_decoder(16#e2#)) OR
 					(reg_q1013 AND symb_decoder(16#f1#)) OR
 					(reg_q1013 AND symb_decoder(16#cb#)) OR
 					(reg_q1013 AND symb_decoder(16#4c#)) OR
 					(reg_q1013 AND symb_decoder(16#14#)) OR
 					(reg_q1013 AND symb_decoder(16#22#)) OR
 					(reg_q1013 AND symb_decoder(16#c6#)) OR
 					(reg_q1013 AND symb_decoder(16#c2#)) OR
 					(reg_q1013 AND symb_decoder(16#c1#)) OR
 					(reg_q1013 AND symb_decoder(16#cd#)) OR
 					(reg_q1013 AND symb_decoder(16#54#)) OR
 					(reg_q1013 AND symb_decoder(16#df#)) OR
 					(reg_q1013 AND symb_decoder(16#35#)) OR
 					(reg_q1013 AND symb_decoder(16#4a#)) OR
 					(reg_q1013 AND symb_decoder(16#3e#)) OR
 					(reg_q1013 AND symb_decoder(16#b2#)) OR
 					(reg_q1013 AND symb_decoder(16#bc#)) OR
 					(reg_q1013 AND symb_decoder(16#63#)) OR
 					(reg_q1013 AND symb_decoder(16#0a#)) OR
 					(reg_q1013 AND symb_decoder(16#e6#)) OR
 					(reg_q1013 AND symb_decoder(16#91#)) OR
 					(reg_q1013 AND symb_decoder(16#0e#)) OR
 					(reg_q1013 AND symb_decoder(16#64#)) OR
 					(reg_q1013 AND symb_decoder(16#05#)) OR
 					(reg_q1013 AND symb_decoder(16#c9#)) OR
 					(reg_q1013 AND symb_decoder(16#5a#)) OR
 					(reg_q1013 AND symb_decoder(16#cf#)) OR
 					(reg_q1013 AND symb_decoder(16#ca#)) OR
 					(reg_q1013 AND symb_decoder(16#ff#)) OR
 					(reg_q1013 AND symb_decoder(16#23#)) OR
 					(reg_q1013 AND symb_decoder(16#4f#)) OR
 					(reg_q1013 AND symb_decoder(16#61#)) OR
 					(reg_q1013 AND symb_decoder(16#81#)) OR
 					(reg_q1013 AND symb_decoder(16#a6#)) OR
 					(reg_q1013 AND symb_decoder(16#6d#)) OR
 					(reg_q1013 AND symb_decoder(16#d2#)) OR
 					(reg_q1013 AND symb_decoder(16#5f#)) OR
 					(reg_q1013 AND symb_decoder(16#d6#)) OR
 					(reg_q1013 AND symb_decoder(16#ef#)) OR
 					(reg_q1013 AND symb_decoder(16#fa#)) OR
 					(reg_q1013 AND symb_decoder(16#2d#)) OR
 					(reg_q1013 AND symb_decoder(16#d4#)) OR
 					(reg_q1013 AND symb_decoder(16#60#)) OR
 					(reg_q1013 AND symb_decoder(16#59#)) OR
 					(reg_q1013 AND symb_decoder(16#57#)) OR
 					(reg_q1013 AND symb_decoder(16#e7#)) OR
 					(reg_q1013 AND symb_decoder(16#97#)) OR
 					(reg_q1013 AND symb_decoder(16#0d#)) OR
 					(reg_q1013 AND symb_decoder(16#c3#)) OR
 					(reg_q1013 AND symb_decoder(16#49#)) OR
 					(reg_q1013 AND symb_decoder(16#c7#)) OR
 					(reg_q1013 AND symb_decoder(16#85#)) OR
 					(reg_q1013 AND symb_decoder(16#48#)) OR
 					(reg_q1013 AND symb_decoder(16#40#)) OR
 					(reg_q1013 AND symb_decoder(16#dc#)) OR
 					(reg_q1013 AND symb_decoder(16#12#)) OR
 					(reg_q1013 AND symb_decoder(16#3a#)) OR
 					(reg_q1013 AND symb_decoder(16#9e#)) OR
 					(reg_q1013 AND symb_decoder(16#c5#)) OR
 					(reg_q1013 AND symb_decoder(16#c4#)) OR
 					(reg_q1013 AND symb_decoder(16#6b#)) OR
 					(reg_q1013 AND symb_decoder(16#e1#)) OR
 					(reg_q1013 AND symb_decoder(16#07#)) OR
 					(reg_q1013 AND symb_decoder(16#db#)) OR
 					(reg_q1013 AND symb_decoder(16#b0#)) OR
 					(reg_q1013 AND symb_decoder(16#27#)) OR
 					(reg_q1013 AND symb_decoder(16#84#)) OR
 					(reg_q1013 AND symb_decoder(16#f9#)) OR
 					(reg_q1013 AND symb_decoder(16#f6#)) OR
 					(reg_q1013 AND symb_decoder(16#82#)) OR
 					(reg_q1013 AND symb_decoder(16#9b#)) OR
 					(reg_q1013 AND symb_decoder(16#9c#)) OR
 					(reg_q1013 AND symb_decoder(16#2a#)) OR
 					(reg_q1013 AND symb_decoder(16#01#)) OR
 					(reg_q1013 AND symb_decoder(16#fc#)) OR
 					(reg_q1013 AND symb_decoder(16#43#)) OR
 					(reg_q1013 AND symb_decoder(16#46#)) OR
 					(reg_q1013 AND symb_decoder(16#70#)) OR
 					(reg_q1013 AND symb_decoder(16#0f#)) OR
 					(reg_q1013 AND symb_decoder(16#98#)) OR
 					(reg_q1013 AND symb_decoder(16#00#)) OR
 					(reg_q1013 AND symb_decoder(16#ab#)) OR
 					(reg_q1013 AND symb_decoder(16#d1#)) OR
 					(reg_q1013 AND symb_decoder(16#c0#)) OR
 					(reg_q1013 AND symb_decoder(16#79#)) OR
 					(reg_q1013 AND symb_decoder(16#2f#)) OR
 					(reg_q1013 AND symb_decoder(16#bf#)) OR
 					(reg_q1013 AND symb_decoder(16#b6#)) OR
 					(reg_q1013 AND symb_decoder(16#a8#)) OR
 					(reg_q1013 AND symb_decoder(16#89#)) OR
 					(reg_q1013 AND symb_decoder(16#95#)) OR
 					(reg_q1013 AND symb_decoder(16#69#)) OR
 					(reg_q1013 AND symb_decoder(16#6e#)) OR
 					(reg_q1013 AND symb_decoder(16#bb#)) OR
 					(reg_q1013 AND symb_decoder(16#ce#)) OR
 					(reg_q1013 AND symb_decoder(16#51#)) OR
 					(reg_q1013 AND symb_decoder(16#8e#)) OR
 					(reg_q1013 AND symb_decoder(16#65#)) OR
 					(reg_q1013 AND symb_decoder(16#02#)) OR
 					(reg_q1013 AND symb_decoder(16#31#)) OR
 					(reg_q1013 AND symb_decoder(16#be#)) OR
 					(reg_q1013 AND symb_decoder(16#af#)) OR
 					(reg_q1013 AND symb_decoder(16#e8#)) OR
 					(reg_q1013 AND symb_decoder(16#fb#)) OR
 					(reg_q1013 AND symb_decoder(16#d7#)) OR
 					(reg_q1013 AND symb_decoder(16#a4#)) OR
 					(reg_q1013 AND symb_decoder(16#45#)) OR
 					(reg_q1013 AND symb_decoder(16#a7#)) OR
 					(reg_q1013 AND symb_decoder(16#1e#)) OR
 					(reg_q1013 AND symb_decoder(16#55#)) OR
 					(reg_q1013 AND symb_decoder(16#4d#)) OR
 					(reg_q1013 AND symb_decoder(16#e0#)) OR
 					(reg_q1013 AND symb_decoder(16#8f#)) OR
 					(reg_q1013 AND symb_decoder(16#4b#)) OR
 					(reg_q1013 AND symb_decoder(16#32#)) OR
 					(reg_q1013 AND symb_decoder(16#7e#)) OR
 					(reg_q1013 AND symb_decoder(16#68#)) OR
 					(reg_q1013 AND symb_decoder(16#6a#)) OR
 					(reg_q1013 AND symb_decoder(16#ed#)) OR
 					(reg_q1013 AND symb_decoder(16#80#)) OR
 					(reg_q1013 AND symb_decoder(16#33#)) OR
 					(reg_q1013 AND symb_decoder(16#29#)) OR
 					(reg_q1013 AND symb_decoder(16#06#)) OR
 					(reg_q1013 AND symb_decoder(16#1a#)) OR
 					(reg_q1013 AND symb_decoder(16#5c#)) OR
 					(reg_q1013 AND symb_decoder(16#87#)) OR
 					(reg_q1013 AND symb_decoder(16#a1#)) OR
 					(reg_q1013 AND symb_decoder(16#74#)) OR
 					(reg_q1013 AND symb_decoder(16#42#)) OR
 					(reg_q1013 AND symb_decoder(16#f4#)) OR
 					(reg_q1013 AND symb_decoder(16#ee#)) OR
 					(reg_q1013 AND symb_decoder(16#73#)) OR
 					(reg_q1013 AND symb_decoder(16#0b#)) OR
 					(reg_q1013 AND symb_decoder(16#7b#)) OR
 					(reg_q1013 AND symb_decoder(16#20#)) OR
 					(reg_q1013 AND symb_decoder(16#76#)) OR
 					(reg_q1013 AND symb_decoder(16#34#)) OR
 					(reg_q1013 AND symb_decoder(16#03#)) OR
 					(reg_q1013 AND symb_decoder(16#30#)) OR
 					(reg_q1013 AND symb_decoder(16#ec#)) OR
 					(reg_q1013 AND symb_decoder(16#28#)) OR
 					(reg_q1013 AND symb_decoder(16#e5#)) OR
 					(reg_q1013 AND symb_decoder(16#5d#)) OR
 					(reg_q1013 AND symb_decoder(16#e3#)) OR
 					(reg_q1013 AND symb_decoder(16#62#)) OR
 					(reg_q1013 AND symb_decoder(16#10#)) OR
 					(reg_q1013 AND symb_decoder(16#88#)) OR
 					(reg_q1013 AND symb_decoder(16#47#)) OR
 					(reg_q1013 AND symb_decoder(16#e9#)) OR
 					(reg_q1013 AND symb_decoder(16#16#)) OR
 					(reg_q1013 AND symb_decoder(16#2e#)) OR
 					(reg_q1013 AND symb_decoder(16#50#)) OR
 					(reg_q1013 AND symb_decoder(16#a0#)) OR
 					(reg_q1013 AND symb_decoder(16#b1#)) OR
 					(reg_q1013 AND symb_decoder(16#96#)) OR
 					(reg_q1013 AND symb_decoder(16#08#)) OR
 					(reg_q1013 AND symb_decoder(16#11#)) OR
 					(reg_q1013 AND symb_decoder(16#1f#)) OR
 					(reg_q1013 AND symb_decoder(16#b5#)) OR
 					(reg_q1013 AND symb_decoder(16#0c#)) OR
 					(reg_q1013 AND symb_decoder(16#83#)) OR
 					(reg_q1013 AND symb_decoder(16#25#)) OR
 					(reg_q1013 AND symb_decoder(16#56#)) OR
 					(reg_q1013 AND symb_decoder(16#86#)) OR
 					(reg_q1013 AND symb_decoder(16#67#)) OR
 					(reg_q1013 AND symb_decoder(16#ac#)) OR
 					(reg_q1013 AND symb_decoder(16#f3#)) OR
 					(reg_q1013 AND symb_decoder(16#3b#)) OR
 					(reg_q1013 AND symb_decoder(16#2b#)) OR
 					(reg_q1013 AND symb_decoder(16#41#)) OR
 					(reg_q1013 AND symb_decoder(16#24#)) OR
 					(reg_q1013 AND symb_decoder(16#9f#)) OR
 					(reg_q1013 AND symb_decoder(16#90#)) OR
 					(reg_q1013 AND symb_decoder(16#15#)) OR
 					(reg_q1013 AND symb_decoder(16#9a#)) OR
 					(reg_q1013 AND symb_decoder(16#3c#)) OR
 					(reg_q1013 AND symb_decoder(16#66#)) OR
 					(reg_q1013 AND symb_decoder(16#13#)) OR
 					(reg_q1013 AND symb_decoder(16#de#)) OR
 					(reg_q1013 AND symb_decoder(16#5b#)) OR
 					(reg_q1013 AND symb_decoder(16#d5#)) OR
 					(reg_q1013 AND symb_decoder(16#93#)) OR
 					(reg_q1013 AND symb_decoder(16#fd#)) OR
 					(reg_q1013 AND symb_decoder(16#bd#)) OR
 					(reg_q1013 AND symb_decoder(16#b7#)) OR
 					(reg_q1013 AND symb_decoder(16#a5#)) OR
 					(reg_q1013 AND symb_decoder(16#92#)) OR
 					(reg_q1013 AND symb_decoder(16#38#)) OR
 					(reg_q1013 AND symb_decoder(16#71#)) OR
 					(reg_q1013 AND symb_decoder(16#04#)) OR
 					(reg_q1013 AND symb_decoder(16#b9#)) OR
 					(reg_q1013 AND symb_decoder(16#58#)) OR
 					(reg_q1013 AND symb_decoder(16#94#)) OR
 					(reg_q1013 AND symb_decoder(16#8d#)) OR
 					(reg_q1013 AND symb_decoder(16#19#)) OR
 					(reg_q1013 AND symb_decoder(16#da#)) OR
 					(reg_q1013 AND symb_decoder(16#fe#)) OR
 					(reg_q1013 AND symb_decoder(16#cc#)) OR
 					(reg_q1013 AND symb_decoder(16#7a#)) OR
 					(reg_q1013 AND symb_decoder(16#f7#)) OR
 					(reg_q1013 AND symb_decoder(16#b8#)) OR
 					(reg_q1013 AND symb_decoder(16#9d#)) OR
 					(reg_q1013 AND symb_decoder(16#d0#)) OR
 					(reg_q1013 AND symb_decoder(16#3d#)) OR
 					(reg_q1013 AND symb_decoder(16#21#)) OR
 					(reg_q1013 AND symb_decoder(16#f0#)) OR
 					(reg_q1013 AND symb_decoder(16#09#)) OR
 					(reg_q1013 AND symb_decoder(16#f2#)) OR
 					(reg_q1013 AND symb_decoder(16#a3#)) OR
 					(reg_q1013 AND symb_decoder(16#aa#)) OR
 					(reg_q1013 AND symb_decoder(16#d8#)) OR
 					(reg_q1013 AND symb_decoder(16#c8#)) OR
 					(reg_q1013 AND symb_decoder(16#5e#)) OR
 					(reg_q1013 AND symb_decoder(16#2c#)) OR
 					(reg_q1013 AND symb_decoder(16#77#)) OR
 					(reg_q1013 AND symb_decoder(16#a2#)) OR
 					(reg_q1013 AND symb_decoder(16#4e#)) OR
 					(reg_q1013 AND symb_decoder(16#52#)) OR
 					(reg_q1013 AND symb_decoder(16#17#)) OR
 					(reg_q1013 AND symb_decoder(16#ae#)) OR
 					(reg_q1013 AND symb_decoder(16#99#)) OR
 					(reg_q1013 AND symb_decoder(16#ba#)) OR
 					(reg_q1013 AND symb_decoder(16#1b#)) OR
 					(reg_q1013 AND symb_decoder(16#3f#)) OR
 					(reg_q1013 AND symb_decoder(16#72#)) OR
 					(reg_q1013 AND symb_decoder(16#78#)) OR
 					(reg_q1013 AND symb_decoder(16#18#)) OR
 					(reg_q1013 AND symb_decoder(16#ea#)) OR
 					(reg_q1013 AND symb_decoder(16#8c#)) OR
 					(reg_q1013 AND symb_decoder(16#39#)) OR
 					(reg_q1013 AND symb_decoder(16#dd#)) OR
 					(reg_q1013 AND symb_decoder(16#ad#)) OR
 					(reg_q1013 AND symb_decoder(16#75#)) OR
 					(reg_q1013 AND symb_decoder(16#6c#)) OR
 					(reg_q1013 AND symb_decoder(16#b3#)) OR
 					(reg_q1013 AND symb_decoder(16#a9#)) OR
 					(reg_q1013 AND symb_decoder(16#7c#));
reg_q1013_init <= '0' ;
	p_reg_q1013: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1013 <= reg_q1013_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1013 <= reg_q1013_init;
        else
          reg_q1013 <= reg_q1013_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q46_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q46 AND symb_decoder(16#5d#)) OR
 					(reg_q46 AND symb_decoder(16#eb#)) OR
 					(reg_q46 AND symb_decoder(16#38#)) OR
 					(reg_q46 AND symb_decoder(16#94#)) OR
 					(reg_q46 AND symb_decoder(16#3a#)) OR
 					(reg_q46 AND symb_decoder(16#50#)) OR
 					(reg_q46 AND symb_decoder(16#60#)) OR
 					(reg_q46 AND symb_decoder(16#37#)) OR
 					(reg_q46 AND symb_decoder(16#ee#)) OR
 					(reg_q46 AND symb_decoder(16#c0#)) OR
 					(reg_q46 AND symb_decoder(16#4b#)) OR
 					(reg_q46 AND symb_decoder(16#b5#)) OR
 					(reg_q46 AND symb_decoder(16#44#)) OR
 					(reg_q46 AND symb_decoder(16#34#)) OR
 					(reg_q46 AND symb_decoder(16#1d#)) OR
 					(reg_q46 AND symb_decoder(16#07#)) OR
 					(reg_q46 AND symb_decoder(16#28#)) OR
 					(reg_q46 AND symb_decoder(16#70#)) OR
 					(reg_q46 AND symb_decoder(16#ed#)) OR
 					(reg_q46 AND symb_decoder(16#bd#)) OR
 					(reg_q46 AND symb_decoder(16#de#)) OR
 					(reg_q46 AND symb_decoder(16#c6#)) OR
 					(reg_q46 AND symb_decoder(16#5e#)) OR
 					(reg_q46 AND symb_decoder(16#74#)) OR
 					(reg_q46 AND symb_decoder(16#55#)) OR
 					(reg_q46 AND symb_decoder(16#ba#)) OR
 					(reg_q46 AND symb_decoder(16#75#)) OR
 					(reg_q46 AND symb_decoder(16#ea#)) OR
 					(reg_q46 AND symb_decoder(16#2d#)) OR
 					(reg_q46 AND symb_decoder(16#81#)) OR
 					(reg_q46 AND symb_decoder(16#2c#)) OR
 					(reg_q46 AND symb_decoder(16#e9#)) OR
 					(reg_q46 AND symb_decoder(16#af#)) OR
 					(reg_q46 AND symb_decoder(16#7c#)) OR
 					(reg_q46 AND symb_decoder(16#d3#)) OR
 					(reg_q46 AND symb_decoder(16#3e#)) OR
 					(reg_q46 AND symb_decoder(16#c5#)) OR
 					(reg_q46 AND symb_decoder(16#b9#)) OR
 					(reg_q46 AND symb_decoder(16#91#)) OR
 					(reg_q46 AND symb_decoder(16#19#)) OR
 					(reg_q46 AND symb_decoder(16#31#)) OR
 					(reg_q46 AND symb_decoder(16#2b#)) OR
 					(reg_q46 AND symb_decoder(16#11#)) OR
 					(reg_q46 AND symb_decoder(16#92#)) OR
 					(reg_q46 AND symb_decoder(16#e3#)) OR
 					(reg_q46 AND symb_decoder(16#9b#)) OR
 					(reg_q46 AND symb_decoder(16#14#)) OR
 					(reg_q46 AND symb_decoder(16#06#)) OR
 					(reg_q46 AND symb_decoder(16#9c#)) OR
 					(reg_q46 AND symb_decoder(16#96#)) OR
 					(reg_q46 AND symb_decoder(16#8e#)) OR
 					(reg_q46 AND symb_decoder(16#e2#)) OR
 					(reg_q46 AND symb_decoder(16#32#)) OR
 					(reg_q46 AND symb_decoder(16#87#)) OR
 					(reg_q46 AND symb_decoder(16#ff#)) OR
 					(reg_q46 AND symb_decoder(16#73#)) OR
 					(reg_q46 AND symb_decoder(16#4f#)) OR
 					(reg_q46 AND symb_decoder(16#76#)) OR
 					(reg_q46 AND symb_decoder(16#39#)) OR
 					(reg_q46 AND symb_decoder(16#7f#)) OR
 					(reg_q46 AND symb_decoder(16#ac#)) OR
 					(reg_q46 AND symb_decoder(16#f7#)) OR
 					(reg_q46 AND symb_decoder(16#f8#)) OR
 					(reg_q46 AND symb_decoder(16#9d#)) OR
 					(reg_q46 AND symb_decoder(16#cb#)) OR
 					(reg_q46 AND symb_decoder(16#86#)) OR
 					(reg_q46 AND symb_decoder(16#d4#)) OR
 					(reg_q46 AND symb_decoder(16#58#)) OR
 					(reg_q46 AND symb_decoder(16#26#)) OR
 					(reg_q46 AND symb_decoder(16#6c#)) OR
 					(reg_q46 AND symb_decoder(16#67#)) OR
 					(reg_q46 AND symb_decoder(16#52#)) OR
 					(reg_q46 AND symb_decoder(16#f3#)) OR
 					(reg_q46 AND symb_decoder(16#22#)) OR
 					(reg_q46 AND symb_decoder(16#c4#)) OR
 					(reg_q46 AND symb_decoder(16#ca#)) OR
 					(reg_q46 AND symb_decoder(16#9f#)) OR
 					(reg_q46 AND symb_decoder(16#db#)) OR
 					(reg_q46 AND symb_decoder(16#98#)) OR
 					(reg_q46 AND symb_decoder(16#0a#)) OR
 					(reg_q46 AND symb_decoder(16#a2#)) OR
 					(reg_q46 AND symb_decoder(16#30#)) OR
 					(reg_q46 AND symb_decoder(16#1b#)) OR
 					(reg_q46 AND symb_decoder(16#88#)) OR
 					(reg_q46 AND symb_decoder(16#8b#)) OR
 					(reg_q46 AND symb_decoder(16#a5#)) OR
 					(reg_q46 AND symb_decoder(16#8d#)) OR
 					(reg_q46 AND symb_decoder(16#dd#)) OR
 					(reg_q46 AND symb_decoder(16#8f#)) OR
 					(reg_q46 AND symb_decoder(16#0b#)) OR
 					(reg_q46 AND symb_decoder(16#4d#)) OR
 					(reg_q46 AND symb_decoder(16#0c#)) OR
 					(reg_q46 AND symb_decoder(16#e8#)) OR
 					(reg_q46 AND symb_decoder(16#84#)) OR
 					(reg_q46 AND symb_decoder(16#79#)) OR
 					(reg_q46 AND symb_decoder(16#53#)) OR
 					(reg_q46 AND symb_decoder(16#64#)) OR
 					(reg_q46 AND symb_decoder(16#2a#)) OR
 					(reg_q46 AND symb_decoder(16#bc#)) OR
 					(reg_q46 AND symb_decoder(16#8a#)) OR
 					(reg_q46 AND symb_decoder(16#fc#)) OR
 					(reg_q46 AND symb_decoder(16#49#)) OR
 					(reg_q46 AND symb_decoder(16#b0#)) OR
 					(reg_q46 AND symb_decoder(16#05#)) OR
 					(reg_q46 AND symb_decoder(16#24#)) OR
 					(reg_q46 AND symb_decoder(16#c7#)) OR
 					(reg_q46 AND symb_decoder(16#3b#)) OR
 					(reg_q46 AND symb_decoder(16#99#)) OR
 					(reg_q46 AND symb_decoder(16#fe#)) OR
 					(reg_q46 AND symb_decoder(16#09#)) OR
 					(reg_q46 AND symb_decoder(16#d2#)) OR
 					(reg_q46 AND symb_decoder(16#b1#)) OR
 					(reg_q46 AND symb_decoder(16#f0#)) OR
 					(reg_q46 AND symb_decoder(16#fb#)) OR
 					(reg_q46 AND symb_decoder(16#42#)) OR
 					(reg_q46 AND symb_decoder(16#be#)) OR
 					(reg_q46 AND symb_decoder(16#59#)) OR
 					(reg_q46 AND symb_decoder(16#1e#)) OR
 					(reg_q46 AND symb_decoder(16#ad#)) OR
 					(reg_q46 AND symb_decoder(16#fa#)) OR
 					(reg_q46 AND symb_decoder(16#56#)) OR
 					(reg_q46 AND symb_decoder(16#18#)) OR
 					(reg_q46 AND symb_decoder(16#aa#)) OR
 					(reg_q46 AND symb_decoder(16#c1#)) OR
 					(reg_q46 AND symb_decoder(16#d6#)) OR
 					(reg_q46 AND symb_decoder(16#43#)) OR
 					(reg_q46 AND symb_decoder(16#9a#)) OR
 					(reg_q46 AND symb_decoder(16#e6#)) OR
 					(reg_q46 AND symb_decoder(16#0e#)) OR
 					(reg_q46 AND symb_decoder(16#e0#)) OR
 					(reg_q46 AND symb_decoder(16#01#)) OR
 					(reg_q46 AND symb_decoder(16#16#)) OR
 					(reg_q46 AND symb_decoder(16#f1#)) OR
 					(reg_q46 AND symb_decoder(16#d8#)) OR
 					(reg_q46 AND symb_decoder(16#4e#)) OR
 					(reg_q46 AND symb_decoder(16#12#)) OR
 					(reg_q46 AND symb_decoder(16#15#)) OR
 					(reg_q46 AND symb_decoder(16#4a#)) OR
 					(reg_q46 AND symb_decoder(16#9e#)) OR
 					(reg_q46 AND symb_decoder(16#ce#)) OR
 					(reg_q46 AND symb_decoder(16#41#)) OR
 					(reg_q46 AND symb_decoder(16#1a#)) OR
 					(reg_q46 AND symb_decoder(16#6b#)) OR
 					(reg_q46 AND symb_decoder(16#c8#)) OR
 					(reg_q46 AND symb_decoder(16#72#)) OR
 					(reg_q46 AND symb_decoder(16#66#)) OR
 					(reg_q46 AND symb_decoder(16#1f#)) OR
 					(reg_q46 AND symb_decoder(16#dc#)) OR
 					(reg_q46 AND symb_decoder(16#e1#)) OR
 					(reg_q46 AND symb_decoder(16#7d#)) OR
 					(reg_q46 AND symb_decoder(16#d9#)) OR
 					(reg_q46 AND symb_decoder(16#ae#)) OR
 					(reg_q46 AND symb_decoder(16#f9#)) OR
 					(reg_q46 AND symb_decoder(16#a9#)) OR
 					(reg_q46 AND symb_decoder(16#48#)) OR
 					(reg_q46 AND symb_decoder(16#02#)) OR
 					(reg_q46 AND symb_decoder(16#b8#)) OR
 					(reg_q46 AND symb_decoder(16#46#)) OR
 					(reg_q46 AND symb_decoder(16#b4#)) OR
 					(reg_q46 AND symb_decoder(16#2e#)) OR
 					(reg_q46 AND symb_decoder(16#8c#)) OR
 					(reg_q46 AND symb_decoder(16#17#)) OR
 					(reg_q46 AND symb_decoder(16#61#)) OR
 					(reg_q46 AND symb_decoder(16#57#)) OR
 					(reg_q46 AND symb_decoder(16#ab#)) OR
 					(reg_q46 AND symb_decoder(16#c2#)) OR
 					(reg_q46 AND symb_decoder(16#5b#)) OR
 					(reg_q46 AND symb_decoder(16#c3#)) OR
 					(reg_q46 AND symb_decoder(16#b6#)) OR
 					(reg_q46 AND symb_decoder(16#5c#)) OR
 					(reg_q46 AND symb_decoder(16#63#)) OR
 					(reg_q46 AND symb_decoder(16#a3#)) OR
 					(reg_q46 AND symb_decoder(16#51#)) OR
 					(reg_q46 AND symb_decoder(16#04#)) OR
 					(reg_q46 AND symb_decoder(16#a6#)) OR
 					(reg_q46 AND symb_decoder(16#78#)) OR
 					(reg_q46 AND symb_decoder(16#4c#)) OR
 					(reg_q46 AND symb_decoder(16#bb#)) OR
 					(reg_q46 AND symb_decoder(16#f2#)) OR
 					(reg_q46 AND symb_decoder(16#95#)) OR
 					(reg_q46 AND symb_decoder(16#d5#)) OR
 					(reg_q46 AND symb_decoder(16#21#)) OR
 					(reg_q46 AND symb_decoder(16#3f#)) OR
 					(reg_q46 AND symb_decoder(16#2f#)) OR
 					(reg_q46 AND symb_decoder(16#cd#)) OR
 					(reg_q46 AND symb_decoder(16#54#)) OR
 					(reg_q46 AND symb_decoder(16#80#)) OR
 					(reg_q46 AND symb_decoder(16#35#)) OR
 					(reg_q46 AND symb_decoder(16#ef#)) OR
 					(reg_q46 AND symb_decoder(16#7b#)) OR
 					(reg_q46 AND symb_decoder(16#25#)) OR
 					(reg_q46 AND symb_decoder(16#85#)) OR
 					(reg_q46 AND symb_decoder(16#68#)) OR
 					(reg_q46 AND symb_decoder(16#13#)) OR
 					(reg_q46 AND symb_decoder(16#33#)) OR
 					(reg_q46 AND symb_decoder(16#62#)) OR
 					(reg_q46 AND symb_decoder(16#a4#)) OR
 					(reg_q46 AND symb_decoder(16#d1#)) OR
 					(reg_q46 AND symb_decoder(16#5f#)) OR
 					(reg_q46 AND symb_decoder(16#7a#)) OR
 					(reg_q46 AND symb_decoder(16#b3#)) OR
 					(reg_q46 AND symb_decoder(16#08#)) OR
 					(reg_q46 AND symb_decoder(16#3c#)) OR
 					(reg_q46 AND symb_decoder(16#e4#)) OR
 					(reg_q46 AND symb_decoder(16#00#)) OR
 					(reg_q46 AND symb_decoder(16#c9#)) OR
 					(reg_q46 AND symb_decoder(16#0d#)) OR
 					(reg_q46 AND symb_decoder(16#7e#)) OR
 					(reg_q46 AND symb_decoder(16#27#)) OR
 					(reg_q46 AND symb_decoder(16#6a#)) OR
 					(reg_q46 AND symb_decoder(16#47#)) OR
 					(reg_q46 AND symb_decoder(16#03#)) OR
 					(reg_q46 AND symb_decoder(16#d0#)) OR
 					(reg_q46 AND symb_decoder(16#69#)) OR
 					(reg_q46 AND symb_decoder(16#e5#)) OR
 					(reg_q46 AND symb_decoder(16#6e#)) OR
 					(reg_q46 AND symb_decoder(16#cf#)) OR
 					(reg_q46 AND symb_decoder(16#83#)) OR
 					(reg_q46 AND symb_decoder(16#5a#)) OR
 					(reg_q46 AND symb_decoder(16#fd#)) OR
 					(reg_q46 AND symb_decoder(16#29#)) OR
 					(reg_q46 AND symb_decoder(16#ec#)) OR
 					(reg_q46 AND symb_decoder(16#f6#)) OR
 					(reg_q46 AND symb_decoder(16#65#)) OR
 					(reg_q46 AND symb_decoder(16#10#)) OR
 					(reg_q46 AND symb_decoder(16#f4#)) OR
 					(reg_q46 AND symb_decoder(16#90#)) OR
 					(reg_q46 AND symb_decoder(16#df#)) OR
 					(reg_q46 AND symb_decoder(16#cc#)) OR
 					(reg_q46 AND symb_decoder(16#89#)) OR
 					(reg_q46 AND symb_decoder(16#82#)) OR
 					(reg_q46 AND symb_decoder(16#b7#)) OR
 					(reg_q46 AND symb_decoder(16#40#)) OR
 					(reg_q46 AND symb_decoder(16#0f#)) OR
 					(reg_q46 AND symb_decoder(16#da#)) OR
 					(reg_q46 AND symb_decoder(16#1c#)) OR
 					(reg_q46 AND symb_decoder(16#d7#)) OR
 					(reg_q46 AND symb_decoder(16#71#)) OR
 					(reg_q46 AND symb_decoder(16#bf#)) OR
 					(reg_q46 AND symb_decoder(16#a1#)) OR
 					(reg_q46 AND symb_decoder(16#93#)) OR
 					(reg_q46 AND symb_decoder(16#36#)) OR
 					(reg_q46 AND symb_decoder(16#6f#)) OR
 					(reg_q46 AND symb_decoder(16#a7#)) OR
 					(reg_q46 AND symb_decoder(16#a0#)) OR
 					(reg_q46 AND symb_decoder(16#3d#)) OR
 					(reg_q46 AND symb_decoder(16#45#)) OR
 					(reg_q46 AND symb_decoder(16#b2#)) OR
 					(reg_q46 AND symb_decoder(16#6d#)) OR
 					(reg_q46 AND symb_decoder(16#e7#)) OR
 					(reg_q46 AND symb_decoder(16#a8#)) OR
 					(reg_q46 AND symb_decoder(16#97#)) OR
 					(reg_q46 AND symb_decoder(16#20#)) OR
 					(reg_q46 AND symb_decoder(16#f5#)) OR
 					(reg_q46 AND symb_decoder(16#77#)) OR
 					(reg_q46 AND symb_decoder(16#23#));
reg_q46_init <= '0' ;
	p_reg_q46: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q46 <= reg_q46_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q46 <= reg_q46_init;
        else
          reg_q46 <= reg_q46_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1050_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1050 AND symb_decoder(16#e7#)) OR
 					(reg_q1050 AND symb_decoder(16#57#)) OR
 					(reg_q1050 AND symb_decoder(16#92#)) OR
 					(reg_q1050 AND symb_decoder(16#c9#)) OR
 					(reg_q1050 AND symb_decoder(16#30#)) OR
 					(reg_q1050 AND symb_decoder(16#d0#)) OR
 					(reg_q1050 AND symb_decoder(16#05#)) OR
 					(reg_q1050 AND symb_decoder(16#61#)) OR
 					(reg_q1050 AND symb_decoder(16#ee#)) OR
 					(reg_q1050 AND symb_decoder(16#4d#)) OR
 					(reg_q1050 AND symb_decoder(16#d8#)) OR
 					(reg_q1050 AND symb_decoder(16#3b#)) OR
 					(reg_q1050 AND symb_decoder(16#0c#)) OR
 					(reg_q1050 AND symb_decoder(16#58#)) OR
 					(reg_q1050 AND symb_decoder(16#12#)) OR
 					(reg_q1050 AND symb_decoder(16#9d#)) OR
 					(reg_q1050 AND symb_decoder(16#45#)) OR
 					(reg_q1050 AND symb_decoder(16#27#)) OR
 					(reg_q1050 AND symb_decoder(16#70#)) OR
 					(reg_q1050 AND symb_decoder(16#6b#)) OR
 					(reg_q1050 AND symb_decoder(16#65#)) OR
 					(reg_q1050 AND symb_decoder(16#9a#)) OR
 					(reg_q1050 AND symb_decoder(16#8b#)) OR
 					(reg_q1050 AND symb_decoder(16#73#)) OR
 					(reg_q1050 AND symb_decoder(16#87#)) OR
 					(reg_q1050 AND symb_decoder(16#f4#)) OR
 					(reg_q1050 AND symb_decoder(16#3f#)) OR
 					(reg_q1050 AND symb_decoder(16#f8#)) OR
 					(reg_q1050 AND symb_decoder(16#a7#)) OR
 					(reg_q1050 AND symb_decoder(16#fe#)) OR
 					(reg_q1050 AND symb_decoder(16#e2#)) OR
 					(reg_q1050 AND symb_decoder(16#dc#)) OR
 					(reg_q1050 AND symb_decoder(16#86#)) OR
 					(reg_q1050 AND symb_decoder(16#a8#)) OR
 					(reg_q1050 AND symb_decoder(16#0e#)) OR
 					(reg_q1050 AND symb_decoder(16#69#)) OR
 					(reg_q1050 AND symb_decoder(16#e4#)) OR
 					(reg_q1050 AND symb_decoder(16#b0#)) OR
 					(reg_q1050 AND symb_decoder(16#8e#)) OR
 					(reg_q1050 AND symb_decoder(16#af#)) OR
 					(reg_q1050 AND symb_decoder(16#0b#)) OR
 					(reg_q1050 AND symb_decoder(16#d3#)) OR
 					(reg_q1050 AND symb_decoder(16#7f#)) OR
 					(reg_q1050 AND symb_decoder(16#34#)) OR
 					(reg_q1050 AND symb_decoder(16#11#)) OR
 					(reg_q1050 AND symb_decoder(16#e6#)) OR
 					(reg_q1050 AND symb_decoder(16#33#)) OR
 					(reg_q1050 AND symb_decoder(16#a0#)) OR
 					(reg_q1050 AND symb_decoder(16#97#)) OR
 					(reg_q1050 AND symb_decoder(16#1c#)) OR
 					(reg_q1050 AND symb_decoder(16#37#)) OR
 					(reg_q1050 AND symb_decoder(16#e3#)) OR
 					(reg_q1050 AND symb_decoder(16#ed#)) OR
 					(reg_q1050 AND symb_decoder(16#ef#)) OR
 					(reg_q1050 AND symb_decoder(16#1a#)) OR
 					(reg_q1050 AND symb_decoder(16#c3#)) OR
 					(reg_q1050 AND symb_decoder(16#b5#)) OR
 					(reg_q1050 AND symb_decoder(16#b3#)) OR
 					(reg_q1050 AND symb_decoder(16#85#)) OR
 					(reg_q1050 AND symb_decoder(16#bd#)) OR
 					(reg_q1050 AND symb_decoder(16#dd#)) OR
 					(reg_q1050 AND symb_decoder(16#40#)) OR
 					(reg_q1050 AND symb_decoder(16#35#)) OR
 					(reg_q1050 AND symb_decoder(16#ac#)) OR
 					(reg_q1050 AND symb_decoder(16#b6#)) OR
 					(reg_q1050 AND symb_decoder(16#ad#)) OR
 					(reg_q1050 AND symb_decoder(16#4f#)) OR
 					(reg_q1050 AND symb_decoder(16#a3#)) OR
 					(reg_q1050 AND symb_decoder(16#39#)) OR
 					(reg_q1050 AND symb_decoder(16#8a#)) OR
 					(reg_q1050 AND symb_decoder(16#0d#)) OR
 					(reg_q1050 AND symb_decoder(16#02#)) OR
 					(reg_q1050 AND symb_decoder(16#20#)) OR
 					(reg_q1050 AND symb_decoder(16#42#)) OR
 					(reg_q1050 AND symb_decoder(16#5f#)) OR
 					(reg_q1050 AND symb_decoder(16#f1#)) OR
 					(reg_q1050 AND symb_decoder(16#53#)) OR
 					(reg_q1050 AND symb_decoder(16#f6#)) OR
 					(reg_q1050 AND symb_decoder(16#e5#)) OR
 					(reg_q1050 AND symb_decoder(16#aa#)) OR
 					(reg_q1050 AND symb_decoder(16#c4#)) OR
 					(reg_q1050 AND symb_decoder(16#cf#)) OR
 					(reg_q1050 AND symb_decoder(16#04#)) OR
 					(reg_q1050 AND symb_decoder(16#de#)) OR
 					(reg_q1050 AND symb_decoder(16#c8#)) OR
 					(reg_q1050 AND symb_decoder(16#8c#)) OR
 					(reg_q1050 AND symb_decoder(16#1b#)) OR
 					(reg_q1050 AND symb_decoder(16#b8#)) OR
 					(reg_q1050 AND symb_decoder(16#6d#)) OR
 					(reg_q1050 AND symb_decoder(16#0f#)) OR
 					(reg_q1050 AND symb_decoder(16#82#)) OR
 					(reg_q1050 AND symb_decoder(16#fb#)) OR
 					(reg_q1050 AND symb_decoder(16#c0#)) OR
 					(reg_q1050 AND symb_decoder(16#75#)) OR
 					(reg_q1050 AND symb_decoder(16#72#)) OR
 					(reg_q1050 AND symb_decoder(16#7d#)) OR
 					(reg_q1050 AND symb_decoder(16#d6#)) OR
 					(reg_q1050 AND symb_decoder(16#eb#)) OR
 					(reg_q1050 AND symb_decoder(16#4c#)) OR
 					(reg_q1050 AND symb_decoder(16#ab#)) OR
 					(reg_q1050 AND symb_decoder(16#b4#)) OR
 					(reg_q1050 AND symb_decoder(16#c7#)) OR
 					(reg_q1050 AND symb_decoder(16#2f#)) OR
 					(reg_q1050 AND symb_decoder(16#c2#)) OR
 					(reg_q1050 AND symb_decoder(16#68#)) OR
 					(reg_q1050 AND symb_decoder(16#a1#)) OR
 					(reg_q1050 AND symb_decoder(16#59#)) OR
 					(reg_q1050 AND symb_decoder(16#b9#)) OR
 					(reg_q1050 AND symb_decoder(16#7a#)) OR
 					(reg_q1050 AND symb_decoder(16#df#)) OR
 					(reg_q1050 AND symb_decoder(16#2d#)) OR
 					(reg_q1050 AND symb_decoder(16#b1#)) OR
 					(reg_q1050 AND symb_decoder(16#0a#)) OR
 					(reg_q1050 AND symb_decoder(16#14#)) OR
 					(reg_q1050 AND symb_decoder(16#b7#)) OR
 					(reg_q1050 AND symb_decoder(16#d9#)) OR
 					(reg_q1050 AND symb_decoder(16#6f#)) OR
 					(reg_q1050 AND symb_decoder(16#19#)) OR
 					(reg_q1050 AND symb_decoder(16#2e#)) OR
 					(reg_q1050 AND symb_decoder(16#6c#)) OR
 					(reg_q1050 AND symb_decoder(16#2b#)) OR
 					(reg_q1050 AND symb_decoder(16#17#)) OR
 					(reg_q1050 AND symb_decoder(16#71#)) OR
 					(reg_q1050 AND symb_decoder(16#7e#)) OR
 					(reg_q1050 AND symb_decoder(16#ce#)) OR
 					(reg_q1050 AND symb_decoder(16#46#)) OR
 					(reg_q1050 AND symb_decoder(16#62#)) OR
 					(reg_q1050 AND symb_decoder(16#18#)) OR
 					(reg_q1050 AND symb_decoder(16#f5#)) OR
 					(reg_q1050 AND symb_decoder(16#ca#)) OR
 					(reg_q1050 AND symb_decoder(16#89#)) OR
 					(reg_q1050 AND symb_decoder(16#15#)) OR
 					(reg_q1050 AND symb_decoder(16#50#)) OR
 					(reg_q1050 AND symb_decoder(16#be#)) OR
 					(reg_q1050 AND symb_decoder(16#29#)) OR
 					(reg_q1050 AND symb_decoder(16#55#)) OR
 					(reg_q1050 AND symb_decoder(16#94#)) OR
 					(reg_q1050 AND symb_decoder(16#21#)) OR
 					(reg_q1050 AND symb_decoder(16#e0#)) OR
 					(reg_q1050 AND symb_decoder(16#1d#)) OR
 					(reg_q1050 AND symb_decoder(16#c6#)) OR
 					(reg_q1050 AND symb_decoder(16#8d#)) OR
 					(reg_q1050 AND symb_decoder(16#cd#)) OR
 					(reg_q1050 AND symb_decoder(16#54#)) OR
 					(reg_q1050 AND symb_decoder(16#36#)) OR
 					(reg_q1050 AND symb_decoder(16#07#)) OR
 					(reg_q1050 AND symb_decoder(16#6e#)) OR
 					(reg_q1050 AND symb_decoder(16#ec#)) OR
 					(reg_q1050 AND symb_decoder(16#6a#)) OR
 					(reg_q1050 AND symb_decoder(16#83#)) OR
 					(reg_q1050 AND symb_decoder(16#d1#)) OR
 					(reg_q1050 AND symb_decoder(16#b2#)) OR
 					(reg_q1050 AND symb_decoder(16#24#)) OR
 					(reg_q1050 AND symb_decoder(16#db#)) OR
 					(reg_q1050 AND symb_decoder(16#fd#)) OR
 					(reg_q1050 AND symb_decoder(16#da#)) OR
 					(reg_q1050 AND symb_decoder(16#64#)) OR
 					(reg_q1050 AND symb_decoder(16#2c#)) OR
 					(reg_q1050 AND symb_decoder(16#ea#)) OR
 					(reg_q1050 AND symb_decoder(16#5b#)) OR
 					(reg_q1050 AND symb_decoder(16#ae#)) OR
 					(reg_q1050 AND symb_decoder(16#25#)) OR
 					(reg_q1050 AND symb_decoder(16#1e#)) OR
 					(reg_q1050 AND symb_decoder(16#fc#)) OR
 					(reg_q1050 AND symb_decoder(16#5e#)) OR
 					(reg_q1050 AND symb_decoder(16#38#)) OR
 					(reg_q1050 AND symb_decoder(16#44#)) OR
 					(reg_q1050 AND symb_decoder(16#63#)) OR
 					(reg_q1050 AND symb_decoder(16#e1#)) OR
 					(reg_q1050 AND symb_decoder(16#5c#)) OR
 					(reg_q1050 AND symb_decoder(16#48#)) OR
 					(reg_q1050 AND symb_decoder(16#ff#)) OR
 					(reg_q1050 AND symb_decoder(16#d7#)) OR
 					(reg_q1050 AND symb_decoder(16#99#)) OR
 					(reg_q1050 AND symb_decoder(16#3c#)) OR
 					(reg_q1050 AND symb_decoder(16#22#)) OR
 					(reg_q1050 AND symb_decoder(16#3e#)) OR
 					(reg_q1050 AND symb_decoder(16#56#)) OR
 					(reg_q1050 AND symb_decoder(16#d4#)) OR
 					(reg_q1050 AND symb_decoder(16#9e#)) OR
 					(reg_q1050 AND symb_decoder(16#23#)) OR
 					(reg_q1050 AND symb_decoder(16#74#)) OR
 					(reg_q1050 AND symb_decoder(16#a9#)) OR
 					(reg_q1050 AND symb_decoder(16#f2#)) OR
 					(reg_q1050 AND symb_decoder(16#28#)) OR
 					(reg_q1050 AND symb_decoder(16#2a#)) OR
 					(reg_q1050 AND symb_decoder(16#96#)) OR
 					(reg_q1050 AND symb_decoder(16#bf#)) OR
 					(reg_q1050 AND symb_decoder(16#08#)) OR
 					(reg_q1050 AND symb_decoder(16#98#)) OR
 					(reg_q1050 AND symb_decoder(16#a5#)) OR
 					(reg_q1050 AND symb_decoder(16#9b#)) OR
 					(reg_q1050 AND symb_decoder(16#43#)) OR
 					(reg_q1050 AND symb_decoder(16#90#)) OR
 					(reg_q1050 AND symb_decoder(16#fa#)) OR
 					(reg_q1050 AND symb_decoder(16#76#)) OR
 					(reg_q1050 AND symb_decoder(16#f0#)) OR
 					(reg_q1050 AND symb_decoder(16#09#)) OR
 					(reg_q1050 AND symb_decoder(16#47#)) OR
 					(reg_q1050 AND symb_decoder(16#10#)) OR
 					(reg_q1050 AND symb_decoder(16#06#)) OR
 					(reg_q1050 AND symb_decoder(16#26#)) OR
 					(reg_q1050 AND symb_decoder(16#a4#)) OR
 					(reg_q1050 AND symb_decoder(16#f7#)) OR
 					(reg_q1050 AND symb_decoder(16#03#)) OR
 					(reg_q1050 AND symb_decoder(16#d5#)) OR
 					(reg_q1050 AND symb_decoder(16#31#)) OR
 					(reg_q1050 AND symb_decoder(16#91#)) OR
 					(reg_q1050 AND symb_decoder(16#8f#)) OR
 					(reg_q1050 AND symb_decoder(16#79#)) OR
 					(reg_q1050 AND symb_decoder(16#52#)) OR
 					(reg_q1050 AND symb_decoder(16#ba#)) OR
 					(reg_q1050 AND symb_decoder(16#1f#)) OR
 					(reg_q1050 AND symb_decoder(16#67#)) OR
 					(reg_q1050 AND symb_decoder(16#f9#)) OR
 					(reg_q1050 AND symb_decoder(16#7b#)) OR
 					(reg_q1050 AND symb_decoder(16#f3#)) OR
 					(reg_q1050 AND symb_decoder(16#32#)) OR
 					(reg_q1050 AND symb_decoder(16#13#)) OR
 					(reg_q1050 AND symb_decoder(16#c5#)) OR
 					(reg_q1050 AND symb_decoder(16#49#)) OR
 					(reg_q1050 AND symb_decoder(16#9c#)) OR
 					(reg_q1050 AND symb_decoder(16#4b#)) OR
 					(reg_q1050 AND symb_decoder(16#bc#)) OR
 					(reg_q1050 AND symb_decoder(16#a6#)) OR
 					(reg_q1050 AND symb_decoder(16#e8#)) OR
 					(reg_q1050 AND symb_decoder(16#81#)) OR
 					(reg_q1050 AND symb_decoder(16#93#)) OR
 					(reg_q1050 AND symb_decoder(16#01#)) OR
 					(reg_q1050 AND symb_decoder(16#88#)) OR
 					(reg_q1050 AND symb_decoder(16#a2#)) OR
 					(reg_q1050 AND symb_decoder(16#51#)) OR
 					(reg_q1050 AND symb_decoder(16#5d#)) OR
 					(reg_q1050 AND symb_decoder(16#bb#)) OR
 					(reg_q1050 AND symb_decoder(16#3a#)) OR
 					(reg_q1050 AND symb_decoder(16#84#)) OR
 					(reg_q1050 AND symb_decoder(16#60#)) OR
 					(reg_q1050 AND symb_decoder(16#16#)) OR
 					(reg_q1050 AND symb_decoder(16#95#)) OR
 					(reg_q1050 AND symb_decoder(16#d2#)) OR
 					(reg_q1050 AND symb_decoder(16#78#)) OR
 					(reg_q1050 AND symb_decoder(16#77#)) OR
 					(reg_q1050 AND symb_decoder(16#00#)) OR
 					(reg_q1050 AND symb_decoder(16#9f#)) OR
 					(reg_q1050 AND symb_decoder(16#41#)) OR
 					(reg_q1050 AND symb_decoder(16#4a#)) OR
 					(reg_q1050 AND symb_decoder(16#cc#)) OR
 					(reg_q1050 AND symb_decoder(16#80#)) OR
 					(reg_q1050 AND symb_decoder(16#5a#)) OR
 					(reg_q1050 AND symb_decoder(16#cb#)) OR
 					(reg_q1050 AND symb_decoder(16#e9#)) OR
 					(reg_q1050 AND symb_decoder(16#c1#)) OR
 					(reg_q1050 AND symb_decoder(16#7c#)) OR
 					(reg_q1050 AND symb_decoder(16#3d#)) OR
 					(reg_q1050 AND symb_decoder(16#4e#)) OR
 					(reg_q1050 AND symb_decoder(16#66#));
reg_q1050_init <= '0' ;
	p_reg_q1050: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1050 <= reg_q1050_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1050 <= reg_q1050_init;
        else
          reg_q1050 <= reg_q1050_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q680_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q680 AND symb_decoder(16#c8#)) OR
 					(reg_q680 AND symb_decoder(16#c4#)) OR
 					(reg_q680 AND symb_decoder(16#27#)) OR
 					(reg_q680 AND symb_decoder(16#33#)) OR
 					(reg_q680 AND symb_decoder(16#98#)) OR
 					(reg_q680 AND symb_decoder(16#bb#)) OR
 					(reg_q680 AND symb_decoder(16#dd#)) OR
 					(reg_q680 AND symb_decoder(16#93#)) OR
 					(reg_q680 AND symb_decoder(16#3b#)) OR
 					(reg_q680 AND symb_decoder(16#6a#)) OR
 					(reg_q680 AND symb_decoder(16#30#)) OR
 					(reg_q680 AND symb_decoder(16#07#)) OR
 					(reg_q680 AND symb_decoder(16#68#)) OR
 					(reg_q680 AND symb_decoder(16#43#)) OR
 					(reg_q680 AND symb_decoder(16#f8#)) OR
 					(reg_q680 AND symb_decoder(16#81#)) OR
 					(reg_q680 AND symb_decoder(16#b3#)) OR
 					(reg_q680 AND symb_decoder(16#be#)) OR
 					(reg_q680 AND symb_decoder(16#24#)) OR
 					(reg_q680 AND symb_decoder(16#7a#)) OR
 					(reg_q680 AND symb_decoder(16#a1#)) OR
 					(reg_q680 AND symb_decoder(16#2d#)) OR
 					(reg_q680 AND symb_decoder(16#ee#)) OR
 					(reg_q680 AND symb_decoder(16#67#)) OR
 					(reg_q680 AND symb_decoder(16#72#)) OR
 					(reg_q680 AND symb_decoder(16#e6#)) OR
 					(reg_q680 AND symb_decoder(16#4b#)) OR
 					(reg_q680 AND symb_decoder(16#02#)) OR
 					(reg_q680 AND symb_decoder(16#70#)) OR
 					(reg_q680 AND symb_decoder(16#ec#)) OR
 					(reg_q680 AND symb_decoder(16#f3#)) OR
 					(reg_q680 AND symb_decoder(16#7b#)) OR
 					(reg_q680 AND symb_decoder(16#56#)) OR
 					(reg_q680 AND symb_decoder(16#73#)) OR
 					(reg_q680 AND symb_decoder(16#d5#)) OR
 					(reg_q680 AND symb_decoder(16#6f#)) OR
 					(reg_q680 AND symb_decoder(16#a9#)) OR
 					(reg_q680 AND symb_decoder(16#6b#)) OR
 					(reg_q680 AND symb_decoder(16#1b#)) OR
 					(reg_q680 AND symb_decoder(16#17#)) OR
 					(reg_q680 AND symb_decoder(16#09#)) OR
 					(reg_q680 AND symb_decoder(16#34#)) OR
 					(reg_q680 AND symb_decoder(16#9e#)) OR
 					(reg_q680 AND symb_decoder(16#60#)) OR
 					(reg_q680 AND symb_decoder(16#2c#)) OR
 					(reg_q680 AND symb_decoder(16#76#)) OR
 					(reg_q680 AND symb_decoder(16#78#)) OR
 					(reg_q680 AND symb_decoder(16#74#)) OR
 					(reg_q680 AND symb_decoder(16#e3#)) OR
 					(reg_q680 AND symb_decoder(16#03#)) OR
 					(reg_q680 AND symb_decoder(16#f7#)) OR
 					(reg_q680 AND symb_decoder(16#9b#)) OR
 					(reg_q680 AND symb_decoder(16#6d#)) OR
 					(reg_q680 AND symb_decoder(16#22#)) OR
 					(reg_q680 AND symb_decoder(16#0e#)) OR
 					(reg_q680 AND symb_decoder(16#cc#)) OR
 					(reg_q680 AND symb_decoder(16#49#)) OR
 					(reg_q680 AND symb_decoder(16#f4#)) OR
 					(reg_q680 AND symb_decoder(16#b8#)) OR
 					(reg_q680 AND symb_decoder(16#80#)) OR
 					(reg_q680 AND symb_decoder(16#57#)) OR
 					(reg_q680 AND symb_decoder(16#d9#)) OR
 					(reg_q680 AND symb_decoder(16#64#)) OR
 					(reg_q680 AND symb_decoder(16#5b#)) OR
 					(reg_q680 AND symb_decoder(16#90#)) OR
 					(reg_q680 AND symb_decoder(16#b9#)) OR
 					(reg_q680 AND symb_decoder(16#79#)) OR
 					(reg_q680 AND symb_decoder(16#bc#)) OR
 					(reg_q680 AND symb_decoder(16#16#)) OR
 					(reg_q680 AND symb_decoder(16#12#)) OR
 					(reg_q680 AND symb_decoder(16#fd#)) OR
 					(reg_q680 AND symb_decoder(16#31#)) OR
 					(reg_q680 AND symb_decoder(16#d0#)) OR
 					(reg_q680 AND symb_decoder(16#aa#)) OR
 					(reg_q680 AND symb_decoder(16#e2#)) OR
 					(reg_q680 AND symb_decoder(16#b2#)) OR
 					(reg_q680 AND symb_decoder(16#45#)) OR
 					(reg_q680 AND symb_decoder(16#c6#)) OR
 					(reg_q680 AND symb_decoder(16#fb#)) OR
 					(reg_q680 AND symb_decoder(16#e4#)) OR
 					(reg_q680 AND symb_decoder(16#fa#)) OR
 					(reg_q680 AND symb_decoder(16#55#)) OR
 					(reg_q680 AND symb_decoder(16#04#)) OR
 					(reg_q680 AND symb_decoder(16#da#)) OR
 					(reg_q680 AND symb_decoder(16#a7#)) OR
 					(reg_q680 AND symb_decoder(16#4f#)) OR
 					(reg_q680 AND symb_decoder(16#b0#)) OR
 					(reg_q680 AND symb_decoder(16#0d#)) OR
 					(reg_q680 AND symb_decoder(16#e8#)) OR
 					(reg_q680 AND symb_decoder(16#96#)) OR
 					(reg_q680 AND symb_decoder(16#db#)) OR
 					(reg_q680 AND symb_decoder(16#7f#)) OR
 					(reg_q680 AND symb_decoder(16#f9#)) OR
 					(reg_q680 AND symb_decoder(16#d6#)) OR
 					(reg_q680 AND symb_decoder(16#37#)) OR
 					(reg_q680 AND symb_decoder(16#2e#)) OR
 					(reg_q680 AND symb_decoder(16#95#)) OR
 					(reg_q680 AND symb_decoder(16#b5#)) OR
 					(reg_q680 AND symb_decoder(16#1a#)) OR
 					(reg_q680 AND symb_decoder(16#32#)) OR
 					(reg_q680 AND symb_decoder(16#21#)) OR
 					(reg_q680 AND symb_decoder(16#cf#)) OR
 					(reg_q680 AND symb_decoder(16#d8#)) OR
 					(reg_q680 AND symb_decoder(16#3e#)) OR
 					(reg_q680 AND symb_decoder(16#f0#)) OR
 					(reg_q680 AND symb_decoder(16#66#)) OR
 					(reg_q680 AND symb_decoder(16#63#)) OR
 					(reg_q680 AND symb_decoder(16#f5#)) OR
 					(reg_q680 AND symb_decoder(16#f6#)) OR
 					(reg_q680 AND symb_decoder(16#47#)) OR
 					(reg_q680 AND symb_decoder(16#51#)) OR
 					(reg_q680 AND symb_decoder(16#15#)) OR
 					(reg_q680 AND symb_decoder(16#5f#)) OR
 					(reg_q680 AND symb_decoder(16#ab#)) OR
 					(reg_q680 AND symb_decoder(16#01#)) OR
 					(reg_q680 AND symb_decoder(16#50#)) OR
 					(reg_q680 AND symb_decoder(16#3f#)) OR
 					(reg_q680 AND symb_decoder(16#25#)) OR
 					(reg_q680 AND symb_decoder(16#69#)) OR
 					(reg_q680 AND symb_decoder(16#a2#)) OR
 					(reg_q680 AND symb_decoder(16#0b#)) OR
 					(reg_q680 AND symb_decoder(16#40#)) OR
 					(reg_q680 AND symb_decoder(16#a6#)) OR
 					(reg_q680 AND symb_decoder(16#7d#)) OR
 					(reg_q680 AND symb_decoder(16#9c#)) OR
 					(reg_q680 AND symb_decoder(16#c9#)) OR
 					(reg_q680 AND symb_decoder(16#f2#)) OR
 					(reg_q680 AND symb_decoder(16#6e#)) OR
 					(reg_q680 AND symb_decoder(16#4e#)) OR
 					(reg_q680 AND symb_decoder(16#10#)) OR
 					(reg_q680 AND symb_decoder(16#5e#)) OR
 					(reg_q680 AND symb_decoder(16#b4#)) OR
 					(reg_q680 AND symb_decoder(16#ce#)) OR
 					(reg_q680 AND symb_decoder(16#05#)) OR
 					(reg_q680 AND symb_decoder(16#06#)) OR
 					(reg_q680 AND symb_decoder(16#a5#)) OR
 					(reg_q680 AND symb_decoder(16#e1#)) OR
 					(reg_q680 AND symb_decoder(16#71#)) OR
 					(reg_q680 AND symb_decoder(16#8c#)) OR
 					(reg_q680 AND symb_decoder(16#b6#)) OR
 					(reg_q680 AND symb_decoder(16#3a#)) OR
 					(reg_q680 AND symb_decoder(16#39#)) OR
 					(reg_q680 AND symb_decoder(16#82#)) OR
 					(reg_q680 AND symb_decoder(16#2a#)) OR
 					(reg_q680 AND symb_decoder(16#88#)) OR
 					(reg_q680 AND symb_decoder(16#de#)) OR
 					(reg_q680 AND symb_decoder(16#5d#)) OR
 					(reg_q680 AND symb_decoder(16#99#)) OR
 					(reg_q680 AND symb_decoder(16#84#)) OR
 					(reg_q680 AND symb_decoder(16#ba#)) OR
 					(reg_q680 AND symb_decoder(16#d1#)) OR
 					(reg_q680 AND symb_decoder(16#9f#)) OR
 					(reg_q680 AND symb_decoder(16#c3#)) OR
 					(reg_q680 AND symb_decoder(16#4d#)) OR
 					(reg_q680 AND symb_decoder(16#42#)) OR
 					(reg_q680 AND symb_decoder(16#df#)) OR
 					(reg_q680 AND symb_decoder(16#26#)) OR
 					(reg_q680 AND symb_decoder(16#1c#)) OR
 					(reg_q680 AND symb_decoder(16#92#)) OR
 					(reg_q680 AND symb_decoder(16#44#)) OR
 					(reg_q680 AND symb_decoder(16#48#)) OR
 					(reg_q680 AND symb_decoder(16#1d#)) OR
 					(reg_q680 AND symb_decoder(16#61#)) OR
 					(reg_q680 AND symb_decoder(16#11#)) OR
 					(reg_q680 AND symb_decoder(16#38#)) OR
 					(reg_q680 AND symb_decoder(16#ae#)) OR
 					(reg_q680 AND symb_decoder(16#13#)) OR
 					(reg_q680 AND symb_decoder(16#65#)) OR
 					(reg_q680 AND symb_decoder(16#bf#)) OR
 					(reg_q680 AND symb_decoder(16#c7#)) OR
 					(reg_q680 AND symb_decoder(16#bd#)) OR
 					(reg_q680 AND symb_decoder(16#7e#)) OR
 					(reg_q680 AND symb_decoder(16#53#)) OR
 					(reg_q680 AND symb_decoder(16#ad#)) OR
 					(reg_q680 AND symb_decoder(16#e0#)) OR
 					(reg_q680 AND symb_decoder(16#ff#)) OR
 					(reg_q680 AND symb_decoder(16#0f#)) OR
 					(reg_q680 AND symb_decoder(16#77#)) OR
 					(reg_q680 AND symb_decoder(16#0c#)) OR
 					(reg_q680 AND symb_decoder(16#14#)) OR
 					(reg_q680 AND symb_decoder(16#5c#)) OR
 					(reg_q680 AND symb_decoder(16#d7#)) OR
 					(reg_q680 AND symb_decoder(16#cb#)) OR
 					(reg_q680 AND symb_decoder(16#91#)) OR
 					(reg_q680 AND symb_decoder(16#62#)) OR
 					(reg_q680 AND symb_decoder(16#19#)) OR
 					(reg_q680 AND symb_decoder(16#ea#)) OR
 					(reg_q680 AND symb_decoder(16#ca#)) OR
 					(reg_q680 AND symb_decoder(16#0a#)) OR
 					(reg_q680 AND symb_decoder(16#97#)) OR
 					(reg_q680 AND symb_decoder(16#af#)) OR
 					(reg_q680 AND symb_decoder(16#3c#)) OR
 					(reg_q680 AND symb_decoder(16#1f#)) OR
 					(reg_q680 AND symb_decoder(16#87#)) OR
 					(reg_q680 AND symb_decoder(16#59#)) OR
 					(reg_q680 AND symb_decoder(16#4a#)) OR
 					(reg_q680 AND symb_decoder(16#6c#)) OR
 					(reg_q680 AND symb_decoder(16#8d#)) OR
 					(reg_q680 AND symb_decoder(16#35#)) OR
 					(reg_q680 AND symb_decoder(16#2b#)) OR
 					(reg_q680 AND symb_decoder(16#20#)) OR
 					(reg_q680 AND symb_decoder(16#ef#)) OR
 					(reg_q680 AND symb_decoder(16#7c#)) OR
 					(reg_q680 AND symb_decoder(16#ac#)) OR
 					(reg_q680 AND symb_decoder(16#c1#)) OR
 					(reg_q680 AND symb_decoder(16#89#)) OR
 					(reg_q680 AND symb_decoder(16#8e#)) OR
 					(reg_q680 AND symb_decoder(16#c5#)) OR
 					(reg_q680 AND symb_decoder(16#94#)) OR
 					(reg_q680 AND symb_decoder(16#83#)) OR
 					(reg_q680 AND symb_decoder(16#a3#)) OR
 					(reg_q680 AND symb_decoder(16#23#)) OR
 					(reg_q680 AND symb_decoder(16#d3#)) OR
 					(reg_q680 AND symb_decoder(16#5a#)) OR
 					(reg_q680 AND symb_decoder(16#75#)) OR
 					(reg_q680 AND symb_decoder(16#2f#)) OR
 					(reg_q680 AND symb_decoder(16#d4#)) OR
 					(reg_q680 AND symb_decoder(16#18#)) OR
 					(reg_q680 AND symb_decoder(16#b7#)) OR
 					(reg_q680 AND symb_decoder(16#41#)) OR
 					(reg_q680 AND symb_decoder(16#00#)) OR
 					(reg_q680 AND symb_decoder(16#8a#)) OR
 					(reg_q680 AND symb_decoder(16#52#)) OR
 					(reg_q680 AND symb_decoder(16#9a#)) OR
 					(reg_q680 AND symb_decoder(16#a4#)) OR
 					(reg_q680 AND symb_decoder(16#28#)) OR
 					(reg_q680 AND symb_decoder(16#fe#)) OR
 					(reg_q680 AND symb_decoder(16#f1#)) OR
 					(reg_q680 AND symb_decoder(16#58#)) OR
 					(reg_q680 AND symb_decoder(16#c0#)) OR
 					(reg_q680 AND symb_decoder(16#a8#)) OR
 					(reg_q680 AND symb_decoder(16#1e#)) OR
 					(reg_q680 AND symb_decoder(16#85#)) OR
 					(reg_q680 AND symb_decoder(16#46#)) OR
 					(reg_q680 AND symb_decoder(16#e5#)) OR
 					(reg_q680 AND symb_decoder(16#3d#)) OR
 					(reg_q680 AND symb_decoder(16#8f#)) OR
 					(reg_q680 AND symb_decoder(16#ed#)) OR
 					(reg_q680 AND symb_decoder(16#d2#)) OR
 					(reg_q680 AND symb_decoder(16#8b#)) OR
 					(reg_q680 AND symb_decoder(16#cd#)) OR
 					(reg_q680 AND symb_decoder(16#54#)) OR
 					(reg_q680 AND symb_decoder(16#9d#)) OR
 					(reg_q680 AND symb_decoder(16#e7#)) OR
 					(reg_q680 AND symb_decoder(16#86#)) OR
 					(reg_q680 AND symb_decoder(16#4c#)) OR
 					(reg_q680 AND symb_decoder(16#e9#)) OR
 					(reg_q680 AND symb_decoder(16#c2#)) OR
 					(reg_q680 AND symb_decoder(16#dc#)) OR
 					(reg_q680 AND symb_decoder(16#36#)) OR
 					(reg_q680 AND symb_decoder(16#b1#)) OR
 					(reg_q680 AND symb_decoder(16#a0#)) OR
 					(reg_q680 AND symb_decoder(16#08#)) OR
 					(reg_q680 AND symb_decoder(16#eb#)) OR
 					(reg_q680 AND symb_decoder(16#29#)) OR
 					(reg_q680 AND symb_decoder(16#fc#));
reg_q680_init <= '0' ;
	p_reg_q680: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q680 <= reg_q680_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q680 <= reg_q680_init;
        else
          reg_q680 <= reg_q680_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1521_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1521 AND symb_decoder(16#56#)) OR
 					(reg_q1521 AND symb_decoder(16#b7#)) OR
 					(reg_q1521 AND symb_decoder(16#6c#)) OR
 					(reg_q1521 AND symb_decoder(16#90#)) OR
 					(reg_q1521 AND symb_decoder(16#39#)) OR
 					(reg_q1521 AND symb_decoder(16#52#)) OR
 					(reg_q1521 AND symb_decoder(16#87#)) OR
 					(reg_q1521 AND symb_decoder(16#35#)) OR
 					(reg_q1521 AND symb_decoder(16#ea#)) OR
 					(reg_q1521 AND symb_decoder(16#b3#)) OR
 					(reg_q1521 AND symb_decoder(16#62#)) OR
 					(reg_q1521 AND symb_decoder(16#a9#)) OR
 					(reg_q1521 AND symb_decoder(16#ed#)) OR
 					(reg_q1521 AND symb_decoder(16#2e#)) OR
 					(reg_q1521 AND symb_decoder(16#e4#)) OR
 					(reg_q1521 AND symb_decoder(16#31#)) OR
 					(reg_q1521 AND symb_decoder(16#8f#)) OR
 					(reg_q1521 AND symb_decoder(16#6b#)) OR
 					(reg_q1521 AND symb_decoder(16#9d#)) OR
 					(reg_q1521 AND symb_decoder(16#1c#)) OR
 					(reg_q1521 AND symb_decoder(16#55#)) OR
 					(reg_q1521 AND symb_decoder(16#f2#)) OR
 					(reg_q1521 AND symb_decoder(16#d7#)) OR
 					(reg_q1521 AND symb_decoder(16#d6#)) OR
 					(reg_q1521 AND symb_decoder(16#cb#)) OR
 					(reg_q1521 AND symb_decoder(16#d2#)) OR
 					(reg_q1521 AND symb_decoder(16#79#)) OR
 					(reg_q1521 AND symb_decoder(16#ee#)) OR
 					(reg_q1521 AND symb_decoder(16#95#)) OR
 					(reg_q1521 AND symb_decoder(16#03#)) OR
 					(reg_q1521 AND symb_decoder(16#0d#)) OR
 					(reg_q1521 AND symb_decoder(16#a3#)) OR
 					(reg_q1521 AND symb_decoder(16#4b#)) OR
 					(reg_q1521 AND symb_decoder(16#dd#)) OR
 					(reg_q1521 AND symb_decoder(16#51#)) OR
 					(reg_q1521 AND symb_decoder(16#1a#)) OR
 					(reg_q1521 AND symb_decoder(16#e9#)) OR
 					(reg_q1521 AND symb_decoder(16#e3#)) OR
 					(reg_q1521 AND symb_decoder(16#71#)) OR
 					(reg_q1521 AND symb_decoder(16#de#)) OR
 					(reg_q1521 AND symb_decoder(16#2a#)) OR
 					(reg_q1521 AND symb_decoder(16#06#)) OR
 					(reg_q1521 AND symb_decoder(16#3f#)) OR
 					(reg_q1521 AND symb_decoder(16#78#)) OR
 					(reg_q1521 AND symb_decoder(16#a1#)) OR
 					(reg_q1521 AND symb_decoder(16#aa#)) OR
 					(reg_q1521 AND symb_decoder(16#a6#)) OR
 					(reg_q1521 AND symb_decoder(16#2c#)) OR
 					(reg_q1521 AND symb_decoder(16#cd#)) OR
 					(reg_q1521 AND symb_decoder(16#54#)) OR
 					(reg_q1521 AND symb_decoder(16#1e#)) OR
 					(reg_q1521 AND symb_decoder(16#63#)) OR
 					(reg_q1521 AND symb_decoder(16#cf#)) OR
 					(reg_q1521 AND symb_decoder(16#db#)) OR
 					(reg_q1521 AND symb_decoder(16#5b#)) OR
 					(reg_q1521 AND symb_decoder(16#3d#)) OR
 					(reg_q1521 AND symb_decoder(16#29#)) OR
 					(reg_q1521 AND symb_decoder(16#11#)) OR
 					(reg_q1521 AND symb_decoder(16#5c#)) OR
 					(reg_q1521 AND symb_decoder(16#cc#)) OR
 					(reg_q1521 AND symb_decoder(16#e8#)) OR
 					(reg_q1521 AND symb_decoder(16#f1#)) OR
 					(reg_q1521 AND symb_decoder(16#e2#)) OR
 					(reg_q1521 AND symb_decoder(16#08#)) OR
 					(reg_q1521 AND symb_decoder(16#27#)) OR
 					(reg_q1521 AND symb_decoder(16#80#)) OR
 					(reg_q1521 AND symb_decoder(16#c5#)) OR
 					(reg_q1521 AND symb_decoder(16#7f#)) OR
 					(reg_q1521 AND symb_decoder(16#09#)) OR
 					(reg_q1521 AND symb_decoder(16#f3#)) OR
 					(reg_q1521 AND symb_decoder(16#a8#)) OR
 					(reg_q1521 AND symb_decoder(16#4f#)) OR
 					(reg_q1521 AND symb_decoder(16#b4#)) OR
 					(reg_q1521 AND symb_decoder(16#f4#)) OR
 					(reg_q1521 AND symb_decoder(16#d4#)) OR
 					(reg_q1521 AND symb_decoder(16#c4#)) OR
 					(reg_q1521 AND symb_decoder(16#2f#)) OR
 					(reg_q1521 AND symb_decoder(16#86#)) OR
 					(reg_q1521 AND symb_decoder(16#eb#)) OR
 					(reg_q1521 AND symb_decoder(16#24#)) OR
 					(reg_q1521 AND symb_decoder(16#58#)) OR
 					(reg_q1521 AND symb_decoder(16#ad#)) OR
 					(reg_q1521 AND symb_decoder(16#da#)) OR
 					(reg_q1521 AND symb_decoder(16#9f#)) OR
 					(reg_q1521 AND symb_decoder(16#43#)) OR
 					(reg_q1521 AND symb_decoder(16#92#)) OR
 					(reg_q1521 AND symb_decoder(16#70#)) OR
 					(reg_q1521 AND symb_decoder(16#a0#)) OR
 					(reg_q1521 AND symb_decoder(16#fc#)) OR
 					(reg_q1521 AND symb_decoder(16#e7#)) OR
 					(reg_q1521 AND symb_decoder(16#ca#)) OR
 					(reg_q1521 AND symb_decoder(16#83#)) OR
 					(reg_q1521 AND symb_decoder(16#85#)) OR
 					(reg_q1521 AND symb_decoder(16#ae#)) OR
 					(reg_q1521 AND symb_decoder(16#19#)) OR
 					(reg_q1521 AND symb_decoder(16#e6#)) OR
 					(reg_q1521 AND symb_decoder(16#c1#)) OR
 					(reg_q1521 AND symb_decoder(16#7e#)) OR
 					(reg_q1521 AND symb_decoder(16#34#)) OR
 					(reg_q1521 AND symb_decoder(16#df#)) OR
 					(reg_q1521 AND symb_decoder(16#4a#)) OR
 					(reg_q1521 AND symb_decoder(16#91#)) OR
 					(reg_q1521 AND symb_decoder(16#16#)) OR
 					(reg_q1521 AND symb_decoder(16#f5#)) OR
 					(reg_q1521 AND symb_decoder(16#ac#)) OR
 					(reg_q1521 AND symb_decoder(16#7b#)) OR
 					(reg_q1521 AND symb_decoder(16#17#)) OR
 					(reg_q1521 AND symb_decoder(16#b5#)) OR
 					(reg_q1521 AND symb_decoder(16#d1#)) OR
 					(reg_q1521 AND symb_decoder(16#b8#)) OR
 					(reg_q1521 AND symb_decoder(16#59#)) OR
 					(reg_q1521 AND symb_decoder(16#e5#)) OR
 					(reg_q1521 AND symb_decoder(16#c0#)) OR
 					(reg_q1521 AND symb_decoder(16#97#)) OR
 					(reg_q1521 AND symb_decoder(16#8c#)) OR
 					(reg_q1521 AND symb_decoder(16#04#)) OR
 					(reg_q1521 AND symb_decoder(16#21#)) OR
 					(reg_q1521 AND symb_decoder(16#25#)) OR
 					(reg_q1521 AND symb_decoder(16#84#)) OR
 					(reg_q1521 AND symb_decoder(16#d5#)) OR
 					(reg_q1521 AND symb_decoder(16#0a#)) OR
 					(reg_q1521 AND symb_decoder(16#00#)) OR
 					(reg_q1521 AND symb_decoder(16#77#)) OR
 					(reg_q1521 AND symb_decoder(16#8a#)) OR
 					(reg_q1521 AND symb_decoder(16#23#)) OR
 					(reg_q1521 AND symb_decoder(16#94#)) OR
 					(reg_q1521 AND symb_decoder(16#68#)) OR
 					(reg_q1521 AND symb_decoder(16#13#)) OR
 					(reg_q1521 AND symb_decoder(16#47#)) OR
 					(reg_q1521 AND symb_decoder(16#d0#)) OR
 					(reg_q1521 AND symb_decoder(16#d9#)) OR
 					(reg_q1521 AND symb_decoder(16#75#)) OR
 					(reg_q1521 AND symb_decoder(16#e1#)) OR
 					(reg_q1521 AND symb_decoder(16#9b#)) OR
 					(reg_q1521 AND symb_decoder(16#89#)) OR
 					(reg_q1521 AND symb_decoder(16#bb#)) OR
 					(reg_q1521 AND symb_decoder(16#d8#)) OR
 					(reg_q1521 AND symb_decoder(16#e0#)) OR
 					(reg_q1521 AND symb_decoder(16#f6#)) OR
 					(reg_q1521 AND symb_decoder(16#f7#)) OR
 					(reg_q1521 AND symb_decoder(16#20#)) OR
 					(reg_q1521 AND symb_decoder(16#41#)) OR
 					(reg_q1521 AND symb_decoder(16#07#)) OR
 					(reg_q1521 AND symb_decoder(16#49#)) OR
 					(reg_q1521 AND symb_decoder(16#ef#)) OR
 					(reg_q1521 AND symb_decoder(16#7c#)) OR
 					(reg_q1521 AND symb_decoder(16#12#)) OR
 					(reg_q1521 AND symb_decoder(16#bd#)) OR
 					(reg_q1521 AND symb_decoder(16#37#)) OR
 					(reg_q1521 AND symb_decoder(16#6f#)) OR
 					(reg_q1521 AND symb_decoder(16#be#)) OR
 					(reg_q1521 AND symb_decoder(16#02#)) OR
 					(reg_q1521 AND symb_decoder(16#c7#)) OR
 					(reg_q1521 AND symb_decoder(16#98#)) OR
 					(reg_q1521 AND symb_decoder(16#96#)) OR
 					(reg_q1521 AND symb_decoder(16#6e#)) OR
 					(reg_q1521 AND symb_decoder(16#99#)) OR
 					(reg_q1521 AND symb_decoder(16#a4#)) OR
 					(reg_q1521 AND symb_decoder(16#28#)) OR
 					(reg_q1521 AND symb_decoder(16#b9#)) OR
 					(reg_q1521 AND symb_decoder(16#c6#)) OR
 					(reg_q1521 AND symb_decoder(16#3c#)) OR
 					(reg_q1521 AND symb_decoder(16#01#)) OR
 					(reg_q1521 AND symb_decoder(16#5f#)) OR
 					(reg_q1521 AND symb_decoder(16#4e#)) OR
 					(reg_q1521 AND symb_decoder(16#b2#)) OR
 					(reg_q1521 AND symb_decoder(16#fd#)) OR
 					(reg_q1521 AND symb_decoder(16#10#)) OR
 					(reg_q1521 AND symb_decoder(16#a2#)) OR
 					(reg_q1521 AND symb_decoder(16#af#)) OR
 					(reg_q1521 AND symb_decoder(16#50#)) OR
 					(reg_q1521 AND symb_decoder(16#4d#)) OR
 					(reg_q1521 AND symb_decoder(16#15#)) OR
 					(reg_q1521 AND symb_decoder(16#65#)) OR
 					(reg_q1521 AND symb_decoder(16#fa#)) OR
 					(reg_q1521 AND symb_decoder(16#82#)) OR
 					(reg_q1521 AND symb_decoder(16#f9#)) OR
 					(reg_q1521 AND symb_decoder(16#33#)) OR
 					(reg_q1521 AND symb_decoder(16#61#)) OR
 					(reg_q1521 AND symb_decoder(16#0c#)) OR
 					(reg_q1521 AND symb_decoder(16#9e#)) OR
 					(reg_q1521 AND symb_decoder(16#b1#)) OR
 					(reg_q1521 AND symb_decoder(16#30#)) OR
 					(reg_q1521 AND symb_decoder(16#f8#)) OR
 					(reg_q1521 AND symb_decoder(16#60#)) OR
 					(reg_q1521 AND symb_decoder(16#c2#)) OR
 					(reg_q1521 AND symb_decoder(16#fe#)) OR
 					(reg_q1521 AND symb_decoder(16#14#)) OR
 					(reg_q1521 AND symb_decoder(16#72#)) OR
 					(reg_q1521 AND symb_decoder(16#66#)) OR
 					(reg_q1521 AND symb_decoder(16#44#)) OR
 					(reg_q1521 AND symb_decoder(16#f0#)) OR
 					(reg_q1521 AND symb_decoder(16#26#)) OR
 					(reg_q1521 AND symb_decoder(16#46#)) OR
 					(reg_q1521 AND symb_decoder(16#6d#)) OR
 					(reg_q1521 AND symb_decoder(16#bc#)) OR
 					(reg_q1521 AND symb_decoder(16#88#)) OR
 					(reg_q1521 AND symb_decoder(16#74#)) OR
 					(reg_q1521 AND symb_decoder(16#64#)) OR
 					(reg_q1521 AND symb_decoder(16#0e#)) OR
 					(reg_q1521 AND symb_decoder(16#a5#)) OR
 					(reg_q1521 AND symb_decoder(16#18#)) OR
 					(reg_q1521 AND symb_decoder(16#fb#)) OR
 					(reg_q1521 AND symb_decoder(16#8d#)) OR
 					(reg_q1521 AND symb_decoder(16#bf#)) OR
 					(reg_q1521 AND symb_decoder(16#57#)) OR
 					(reg_q1521 AND symb_decoder(16#c9#)) OR
 					(reg_q1521 AND symb_decoder(16#67#)) OR
 					(reg_q1521 AND symb_decoder(16#ab#)) OR
 					(reg_q1521 AND symb_decoder(16#ec#)) OR
 					(reg_q1521 AND symb_decoder(16#2d#)) OR
 					(reg_q1521 AND symb_decoder(16#45#)) OR
 					(reg_q1521 AND symb_decoder(16#7d#)) OR
 					(reg_q1521 AND symb_decoder(16#c3#)) OR
 					(reg_q1521 AND symb_decoder(16#b6#)) OR
 					(reg_q1521 AND symb_decoder(16#48#)) OR
 					(reg_q1521 AND symb_decoder(16#3e#)) OR
 					(reg_q1521 AND symb_decoder(16#1b#)) OR
 					(reg_q1521 AND symb_decoder(16#1f#)) OR
 					(reg_q1521 AND symb_decoder(16#22#)) OR
 					(reg_q1521 AND symb_decoder(16#36#)) OR
 					(reg_q1521 AND symb_decoder(16#0f#)) OR
 					(reg_q1521 AND symb_decoder(16#b0#)) OR
 					(reg_q1521 AND symb_decoder(16#5d#)) OR
 					(reg_q1521 AND symb_decoder(16#81#)) OR
 					(reg_q1521 AND symb_decoder(16#3b#)) OR
 					(reg_q1521 AND symb_decoder(16#c8#)) OR
 					(reg_q1521 AND symb_decoder(16#ff#)) OR
 					(reg_q1521 AND symb_decoder(16#8b#)) OR
 					(reg_q1521 AND symb_decoder(16#4c#)) OR
 					(reg_q1521 AND symb_decoder(16#38#)) OR
 					(reg_q1521 AND symb_decoder(16#05#)) OR
 					(reg_q1521 AND symb_decoder(16#2b#)) OR
 					(reg_q1521 AND symb_decoder(16#dc#)) OR
 					(reg_q1521 AND symb_decoder(16#53#)) OR
 					(reg_q1521 AND symb_decoder(16#d3#)) OR
 					(reg_q1521 AND symb_decoder(16#40#)) OR
 					(reg_q1521 AND symb_decoder(16#8e#)) OR
 					(reg_q1521 AND symb_decoder(16#6a#)) OR
 					(reg_q1521 AND symb_decoder(16#3a#)) OR
 					(reg_q1521 AND symb_decoder(16#ba#)) OR
 					(reg_q1521 AND symb_decoder(16#69#)) OR
 					(reg_q1521 AND symb_decoder(16#1d#)) OR
 					(reg_q1521 AND symb_decoder(16#76#)) OR
 					(reg_q1521 AND symb_decoder(16#a7#)) OR
 					(reg_q1521 AND symb_decoder(16#ce#)) OR
 					(reg_q1521 AND symb_decoder(16#42#)) OR
 					(reg_q1521 AND symb_decoder(16#5a#)) OR
 					(reg_q1521 AND symb_decoder(16#9c#)) OR
 					(reg_q1521 AND symb_decoder(16#9a#)) OR
 					(reg_q1521 AND symb_decoder(16#5e#)) OR
 					(reg_q1521 AND symb_decoder(16#73#)) OR
 					(reg_q1521 AND symb_decoder(16#32#)) OR
 					(reg_q1521 AND symb_decoder(16#0b#)) OR
 					(reg_q1521 AND symb_decoder(16#93#)) OR
 					(reg_q1521 AND symb_decoder(16#7a#));
reg_q1521_init <= '0' ;
	p_reg_q1521: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1521 <= reg_q1521_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1521 <= reg_q1521_init;
        else
          reg_q1521 <= reg_q1521_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1884_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1884 AND symb_decoder(16#03#)) OR
 					(reg_q1884 AND symb_decoder(16#f5#)) OR
 					(reg_q1884 AND symb_decoder(16#44#)) OR
 					(reg_q1884 AND symb_decoder(16#9a#)) OR
 					(reg_q1884 AND symb_decoder(16#c7#)) OR
 					(reg_q1884 AND symb_decoder(16#10#)) OR
 					(reg_q1884 AND symb_decoder(16#35#)) OR
 					(reg_q1884 AND symb_decoder(16#cc#)) OR
 					(reg_q1884 AND symb_decoder(16#15#)) OR
 					(reg_q1884 AND symb_decoder(16#0a#)) OR
 					(reg_q1884 AND symb_decoder(16#cb#)) OR
 					(reg_q1884 AND symb_decoder(16#77#)) OR
 					(reg_q1884 AND symb_decoder(16#69#)) OR
 					(reg_q1884 AND symb_decoder(16#9f#)) OR
 					(reg_q1884 AND symb_decoder(16#57#)) OR
 					(reg_q1884 AND symb_decoder(16#c9#)) OR
 					(reg_q1884 AND symb_decoder(16#a7#)) OR
 					(reg_q1884 AND symb_decoder(16#4d#)) OR
 					(reg_q1884 AND symb_decoder(16#f1#)) OR
 					(reg_q1884 AND symb_decoder(16#94#)) OR
 					(reg_q1884 AND symb_decoder(16#fc#)) OR
 					(reg_q1884 AND symb_decoder(16#7d#)) OR
 					(reg_q1884 AND symb_decoder(16#41#)) OR
 					(reg_q1884 AND symb_decoder(16#e1#)) OR
 					(reg_q1884 AND symb_decoder(16#12#)) OR
 					(reg_q1884 AND symb_decoder(16#d4#)) OR
 					(reg_q1884 AND symb_decoder(16#f8#)) OR
 					(reg_q1884 AND symb_decoder(16#91#)) OR
 					(reg_q1884 AND symb_decoder(16#71#)) OR
 					(reg_q1884 AND symb_decoder(16#28#)) OR
 					(reg_q1884 AND symb_decoder(16#7b#)) OR
 					(reg_q1884 AND symb_decoder(16#cf#)) OR
 					(reg_q1884 AND symb_decoder(16#d7#)) OR
 					(reg_q1884 AND symb_decoder(16#b3#)) OR
 					(reg_q1884 AND symb_decoder(16#32#)) OR
 					(reg_q1884 AND symb_decoder(16#7e#)) OR
 					(reg_q1884 AND symb_decoder(16#4a#)) OR
 					(reg_q1884 AND symb_decoder(16#7f#)) OR
 					(reg_q1884 AND symb_decoder(16#ba#)) OR
 					(reg_q1884 AND symb_decoder(16#48#)) OR
 					(reg_q1884 AND symb_decoder(16#53#)) OR
 					(reg_q1884 AND symb_decoder(16#1f#)) OR
 					(reg_q1884 AND symb_decoder(16#d6#)) OR
 					(reg_q1884 AND symb_decoder(16#e3#)) OR
 					(reg_q1884 AND symb_decoder(16#84#)) OR
 					(reg_q1884 AND symb_decoder(16#89#)) OR
 					(reg_q1884 AND symb_decoder(16#55#)) OR
 					(reg_q1884 AND symb_decoder(16#2e#)) OR
 					(reg_q1884 AND symb_decoder(16#a2#)) OR
 					(reg_q1884 AND symb_decoder(16#75#)) OR
 					(reg_q1884 AND symb_decoder(16#63#)) OR
 					(reg_q1884 AND symb_decoder(16#09#)) OR
 					(reg_q1884 AND symb_decoder(16#b5#)) OR
 					(reg_q1884 AND symb_decoder(16#d9#)) OR
 					(reg_q1884 AND symb_decoder(16#78#)) OR
 					(reg_q1884 AND symb_decoder(16#9c#)) OR
 					(reg_q1884 AND symb_decoder(16#11#)) OR
 					(reg_q1884 AND symb_decoder(16#22#)) OR
 					(reg_q1884 AND symb_decoder(16#60#)) OR
 					(reg_q1884 AND symb_decoder(16#14#)) OR
 					(reg_q1884 AND symb_decoder(16#39#)) OR
 					(reg_q1884 AND symb_decoder(16#3d#)) OR
 					(reg_q1884 AND symb_decoder(16#d0#)) OR
 					(reg_q1884 AND symb_decoder(16#9e#)) OR
 					(reg_q1884 AND symb_decoder(16#90#)) OR
 					(reg_q1884 AND symb_decoder(16#46#)) OR
 					(reg_q1884 AND symb_decoder(16#42#)) OR
 					(reg_q1884 AND symb_decoder(16#fa#)) OR
 					(reg_q1884 AND symb_decoder(16#bf#)) OR
 					(reg_q1884 AND symb_decoder(16#70#)) OR
 					(reg_q1884 AND symb_decoder(16#3c#)) OR
 					(reg_q1884 AND symb_decoder(16#82#)) OR
 					(reg_q1884 AND symb_decoder(16#49#)) OR
 					(reg_q1884 AND symb_decoder(16#23#)) OR
 					(reg_q1884 AND symb_decoder(16#73#)) OR
 					(reg_q1884 AND symb_decoder(16#4b#)) OR
 					(reg_q1884 AND symb_decoder(16#e8#)) OR
 					(reg_q1884 AND symb_decoder(16#8c#)) OR
 					(reg_q1884 AND symb_decoder(16#ae#)) OR
 					(reg_q1884 AND symb_decoder(16#5c#)) OR
 					(reg_q1884 AND symb_decoder(16#b2#)) OR
 					(reg_q1884 AND symb_decoder(16#aa#)) OR
 					(reg_q1884 AND symb_decoder(16#8d#)) OR
 					(reg_q1884 AND symb_decoder(16#e2#)) OR
 					(reg_q1884 AND symb_decoder(16#d3#)) OR
 					(reg_q1884 AND symb_decoder(16#61#)) OR
 					(reg_q1884 AND symb_decoder(16#b1#)) OR
 					(reg_q1884 AND symb_decoder(16#f3#)) OR
 					(reg_q1884 AND symb_decoder(16#a6#)) OR
 					(reg_q1884 AND symb_decoder(16#6a#)) OR
 					(reg_q1884 AND symb_decoder(16#be#)) OR
 					(reg_q1884 AND symb_decoder(16#dd#)) OR
 					(reg_q1884 AND symb_decoder(16#f6#)) OR
 					(reg_q1884 AND symb_decoder(16#8b#)) OR
 					(reg_q1884 AND symb_decoder(16#db#)) OR
 					(reg_q1884 AND symb_decoder(16#a8#)) OR
 					(reg_q1884 AND symb_decoder(16#4e#)) OR
 					(reg_q1884 AND symb_decoder(16#c3#)) OR
 					(reg_q1884 AND symb_decoder(16#1e#)) OR
 					(reg_q1884 AND symb_decoder(16#ac#)) OR
 					(reg_q1884 AND symb_decoder(16#1c#)) OR
 					(reg_q1884 AND symb_decoder(16#68#)) OR
 					(reg_q1884 AND symb_decoder(16#3f#)) OR
 					(reg_q1884 AND symb_decoder(16#c2#)) OR
 					(reg_q1884 AND symb_decoder(16#b8#)) OR
 					(reg_q1884 AND symb_decoder(16#2a#)) OR
 					(reg_q1884 AND symb_decoder(16#07#)) OR
 					(reg_q1884 AND symb_decoder(16#b6#)) OR
 					(reg_q1884 AND symb_decoder(16#45#)) OR
 					(reg_q1884 AND symb_decoder(16#2f#)) OR
 					(reg_q1884 AND symb_decoder(16#00#)) OR
 					(reg_q1884 AND symb_decoder(16#05#)) OR
 					(reg_q1884 AND symb_decoder(16#79#)) OR
 					(reg_q1884 AND symb_decoder(16#a9#)) OR
 					(reg_q1884 AND symb_decoder(16#98#)) OR
 					(reg_q1884 AND symb_decoder(16#30#)) OR
 					(reg_q1884 AND symb_decoder(16#0b#)) OR
 					(reg_q1884 AND symb_decoder(16#36#)) OR
 					(reg_q1884 AND symb_decoder(16#37#)) OR
 					(reg_q1884 AND symb_decoder(16#66#)) OR
 					(reg_q1884 AND symb_decoder(16#74#)) OR
 					(reg_q1884 AND symb_decoder(16#27#)) OR
 					(reg_q1884 AND symb_decoder(16#52#)) OR
 					(reg_q1884 AND symb_decoder(16#92#)) OR
 					(reg_q1884 AND symb_decoder(16#16#)) OR
 					(reg_q1884 AND symb_decoder(16#e0#)) OR
 					(reg_q1884 AND symb_decoder(16#bc#)) OR
 					(reg_q1884 AND symb_decoder(16#ed#)) OR
 					(reg_q1884 AND symb_decoder(16#83#)) OR
 					(reg_q1884 AND symb_decoder(16#67#)) OR
 					(reg_q1884 AND symb_decoder(16#02#)) OR
 					(reg_q1884 AND symb_decoder(16#34#)) OR
 					(reg_q1884 AND symb_decoder(16#d8#)) OR
 					(reg_q1884 AND symb_decoder(16#9b#)) OR
 					(reg_q1884 AND symb_decoder(16#01#)) OR
 					(reg_q1884 AND symb_decoder(16#c4#)) OR
 					(reg_q1884 AND symb_decoder(16#95#)) OR
 					(reg_q1884 AND symb_decoder(16#76#)) OR
 					(reg_q1884 AND symb_decoder(16#86#)) OR
 					(reg_q1884 AND symb_decoder(16#f9#)) OR
 					(reg_q1884 AND symb_decoder(16#5b#)) OR
 					(reg_q1884 AND symb_decoder(16#7a#)) OR
 					(reg_q1884 AND symb_decoder(16#f0#)) OR
 					(reg_q1884 AND symb_decoder(16#dc#)) OR
 					(reg_q1884 AND symb_decoder(16#56#)) OR
 					(reg_q1884 AND symb_decoder(16#8a#)) OR
 					(reg_q1884 AND symb_decoder(16#e6#)) OR
 					(reg_q1884 AND symb_decoder(16#ff#)) OR
 					(reg_q1884 AND symb_decoder(16#8f#)) OR
 					(reg_q1884 AND symb_decoder(16#25#)) OR
 					(reg_q1884 AND symb_decoder(16#0d#)) OR
 					(reg_q1884 AND symb_decoder(16#eb#)) OR
 					(reg_q1884 AND symb_decoder(16#51#)) OR
 					(reg_q1884 AND symb_decoder(16#a0#)) OR
 					(reg_q1884 AND symb_decoder(16#80#)) OR
 					(reg_q1884 AND symb_decoder(16#04#)) OR
 					(reg_q1884 AND symb_decoder(16#19#)) OR
 					(reg_q1884 AND symb_decoder(16#97#)) OR
 					(reg_q1884 AND symb_decoder(16#a4#)) OR
 					(reg_q1884 AND symb_decoder(16#29#)) OR
 					(reg_q1884 AND symb_decoder(16#bd#)) OR
 					(reg_q1884 AND symb_decoder(16#e7#)) OR
 					(reg_q1884 AND symb_decoder(16#ce#)) OR
 					(reg_q1884 AND symb_decoder(16#20#)) OR
 					(reg_q1884 AND symb_decoder(16#40#)) OR
 					(reg_q1884 AND symb_decoder(16#da#)) OR
 					(reg_q1884 AND symb_decoder(16#a5#)) OR
 					(reg_q1884 AND symb_decoder(16#47#)) OR
 					(reg_q1884 AND symb_decoder(16#58#)) OR
 					(reg_q1884 AND symb_decoder(16#ea#)) OR
 					(reg_q1884 AND symb_decoder(16#3b#)) OR
 					(reg_q1884 AND symb_decoder(16#65#)) OR
 					(reg_q1884 AND symb_decoder(16#ee#)) OR
 					(reg_q1884 AND symb_decoder(16#3e#)) OR
 					(reg_q1884 AND symb_decoder(16#a3#)) OR
 					(reg_q1884 AND symb_decoder(16#b4#)) OR
 					(reg_q1884 AND symb_decoder(16#17#)) OR
 					(reg_q1884 AND symb_decoder(16#e9#)) OR
 					(reg_q1884 AND symb_decoder(16#43#)) OR
 					(reg_q1884 AND symb_decoder(16#0f#)) OR
 					(reg_q1884 AND symb_decoder(16#24#)) OR
 					(reg_q1884 AND symb_decoder(16#e5#)) OR
 					(reg_q1884 AND symb_decoder(16#6d#)) OR
 					(reg_q1884 AND symb_decoder(16#ab#)) OR
 					(reg_q1884 AND symb_decoder(16#ca#)) OR
 					(reg_q1884 AND symb_decoder(16#b9#)) OR
 					(reg_q1884 AND symb_decoder(16#ad#)) OR
 					(reg_q1884 AND symb_decoder(16#62#)) OR
 					(reg_q1884 AND symb_decoder(16#85#)) OR
 					(reg_q1884 AND symb_decoder(16#b7#)) OR
 					(reg_q1884 AND symb_decoder(16#6e#)) OR
 					(reg_q1884 AND symb_decoder(16#18#)) OR
 					(reg_q1884 AND symb_decoder(16#31#)) OR
 					(reg_q1884 AND symb_decoder(16#81#)) OR
 					(reg_q1884 AND symb_decoder(16#9d#)) OR
 					(reg_q1884 AND symb_decoder(16#5a#)) OR
 					(reg_q1884 AND symb_decoder(16#64#)) OR
 					(reg_q1884 AND symb_decoder(16#c8#)) OR
 					(reg_q1884 AND symb_decoder(16#ec#)) OR
 					(reg_q1884 AND symb_decoder(16#26#)) OR
 					(reg_q1884 AND symb_decoder(16#6f#)) OR
 					(reg_q1884 AND symb_decoder(16#1a#)) OR
 					(reg_q1884 AND symb_decoder(16#2d#)) OR
 					(reg_q1884 AND symb_decoder(16#93#)) OR
 					(reg_q1884 AND symb_decoder(16#2c#)) OR
 					(reg_q1884 AND symb_decoder(16#c5#)) OR
 					(reg_q1884 AND symb_decoder(16#d2#)) OR
 					(reg_q1884 AND symb_decoder(16#59#)) OR
 					(reg_q1884 AND symb_decoder(16#21#)) OR
 					(reg_q1884 AND symb_decoder(16#4c#)) OR
 					(reg_q1884 AND symb_decoder(16#de#)) OR
 					(reg_q1884 AND symb_decoder(16#6c#)) OR
 					(reg_q1884 AND symb_decoder(16#a1#)) OR
 					(reg_q1884 AND symb_decoder(16#e4#)) OR
 					(reg_q1884 AND symb_decoder(16#38#)) OR
 					(reg_q1884 AND symb_decoder(16#87#)) OR
 					(reg_q1884 AND symb_decoder(16#c0#)) OR
 					(reg_q1884 AND symb_decoder(16#1d#)) OR
 					(reg_q1884 AND symb_decoder(16#2b#)) OR
 					(reg_q1884 AND symb_decoder(16#3a#)) OR
 					(reg_q1884 AND symb_decoder(16#08#)) OR
 					(reg_q1884 AND symb_decoder(16#f7#)) OR
 					(reg_q1884 AND symb_decoder(16#72#)) OR
 					(reg_q1884 AND symb_decoder(16#fe#)) OR
 					(reg_q1884 AND symb_decoder(16#88#)) OR
 					(reg_q1884 AND symb_decoder(16#5f#)) OR
 					(reg_q1884 AND symb_decoder(16#4f#)) OR
 					(reg_q1884 AND symb_decoder(16#b0#)) OR
 					(reg_q1884 AND symb_decoder(16#06#)) OR
 					(reg_q1884 AND symb_decoder(16#df#)) OR
 					(reg_q1884 AND symb_decoder(16#bb#)) OR
 					(reg_q1884 AND symb_decoder(16#ef#)) OR
 					(reg_q1884 AND symb_decoder(16#cd#)) OR
 					(reg_q1884 AND symb_decoder(16#54#)) OR
 					(reg_q1884 AND symb_decoder(16#fb#)) OR
 					(reg_q1884 AND symb_decoder(16#1b#)) OR
 					(reg_q1884 AND symb_decoder(16#0e#)) OR
 					(reg_q1884 AND symb_decoder(16#7c#)) OR
 					(reg_q1884 AND symb_decoder(16#f2#)) OR
 					(reg_q1884 AND symb_decoder(16#96#)) OR
 					(reg_q1884 AND symb_decoder(16#d5#)) OR
 					(reg_q1884 AND symb_decoder(16#50#)) OR
 					(reg_q1884 AND symb_decoder(16#f4#)) OR
 					(reg_q1884 AND symb_decoder(16#13#)) OR
 					(reg_q1884 AND symb_decoder(16#33#)) OR
 					(reg_q1884 AND symb_decoder(16#5e#)) OR
 					(reg_q1884 AND symb_decoder(16#6b#)) OR
 					(reg_q1884 AND symb_decoder(16#5d#)) OR
 					(reg_q1884 AND symb_decoder(16#0c#)) OR
 					(reg_q1884 AND symb_decoder(16#99#)) OR
 					(reg_q1884 AND symb_decoder(16#d1#)) OR
 					(reg_q1884 AND symb_decoder(16#c1#)) OR
 					(reg_q1884 AND symb_decoder(16#fd#)) OR
 					(reg_q1884 AND symb_decoder(16#af#)) OR
 					(reg_q1884 AND symb_decoder(16#8e#)) OR
 					(reg_q1884 AND symb_decoder(16#c6#));
reg_q1884_init <= '0' ;
	p_reg_q1884: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1884 <= reg_q1884_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1884 <= reg_q1884_init;
        else
          reg_q1884 <= reg_q1884_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1955_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1955 AND symb_decoder(16#3b#)) OR
 					(reg_q1955 AND symb_decoder(16#c2#)) OR
 					(reg_q1955 AND symb_decoder(16#de#)) OR
 					(reg_q1955 AND symb_decoder(16#23#)) OR
 					(reg_q1955 AND symb_decoder(16#a9#)) OR
 					(reg_q1955 AND symb_decoder(16#e2#)) OR
 					(reg_q1955 AND symb_decoder(16#d0#)) OR
 					(reg_q1955 AND symb_decoder(16#ea#)) OR
 					(reg_q1955 AND symb_decoder(16#d8#)) OR
 					(reg_q1955 AND symb_decoder(16#ba#)) OR
 					(reg_q1955 AND symb_decoder(16#f1#)) OR
 					(reg_q1955 AND symb_decoder(16#0f#)) OR
 					(reg_q1955 AND symb_decoder(16#48#)) OR
 					(reg_q1955 AND symb_decoder(16#d3#)) OR
 					(reg_q1955 AND symb_decoder(16#ed#)) OR
 					(reg_q1955 AND symb_decoder(16#d9#)) OR
 					(reg_q1955 AND symb_decoder(16#e8#)) OR
 					(reg_q1955 AND symb_decoder(16#fb#)) OR
 					(reg_q1955 AND symb_decoder(16#ee#)) OR
 					(reg_q1955 AND symb_decoder(16#e3#)) OR
 					(reg_q1955 AND symb_decoder(16#f8#)) OR
 					(reg_q1955 AND symb_decoder(16#b9#)) OR
 					(reg_q1955 AND symb_decoder(16#ab#)) OR
 					(reg_q1955 AND symb_decoder(16#d4#)) OR
 					(reg_q1955 AND symb_decoder(16#a0#)) OR
 					(reg_q1955 AND symb_decoder(16#1a#)) OR
 					(reg_q1955 AND symb_decoder(16#7d#)) OR
 					(reg_q1955 AND symb_decoder(16#c7#)) OR
 					(reg_q1955 AND symb_decoder(16#d2#)) OR
 					(reg_q1955 AND symb_decoder(16#a6#)) OR
 					(reg_q1955 AND symb_decoder(16#b1#)) OR
 					(reg_q1955 AND symb_decoder(16#78#)) OR
 					(reg_q1955 AND symb_decoder(16#06#)) OR
 					(reg_q1955 AND symb_decoder(16#03#)) OR
 					(reg_q1955 AND symb_decoder(16#08#)) OR
 					(reg_q1955 AND symb_decoder(16#3f#)) OR
 					(reg_q1955 AND symb_decoder(16#b8#)) OR
 					(reg_q1955 AND symb_decoder(16#a3#)) OR
 					(reg_q1955 AND symb_decoder(16#e5#)) OR
 					(reg_q1955 AND symb_decoder(16#d7#)) OR
 					(reg_q1955 AND symb_decoder(16#f3#)) OR
 					(reg_q1955 AND symb_decoder(16#c9#)) OR
 					(reg_q1955 AND symb_decoder(16#39#)) OR
 					(reg_q1955 AND symb_decoder(16#5c#)) OR
 					(reg_q1955 AND symb_decoder(16#79#)) OR
 					(reg_q1955 AND symb_decoder(16#2e#)) OR
 					(reg_q1955 AND symb_decoder(16#74#)) OR
 					(reg_q1955 AND symb_decoder(16#8f#)) OR
 					(reg_q1955 AND symb_decoder(16#86#)) OR
 					(reg_q1955 AND symb_decoder(16#da#)) OR
 					(reg_q1955 AND symb_decoder(16#69#)) OR
 					(reg_q1955 AND symb_decoder(16#b3#)) OR
 					(reg_q1955 AND symb_decoder(16#af#)) OR
 					(reg_q1955 AND symb_decoder(16#77#)) OR
 					(reg_q1955 AND symb_decoder(16#59#)) OR
 					(reg_q1955 AND symb_decoder(16#9f#)) OR
 					(reg_q1955 AND symb_decoder(16#49#)) OR
 					(reg_q1955 AND symb_decoder(16#51#)) OR
 					(reg_q1955 AND symb_decoder(16#63#)) OR
 					(reg_q1955 AND symb_decoder(16#be#)) OR
 					(reg_q1955 AND symb_decoder(16#ac#)) OR
 					(reg_q1955 AND symb_decoder(16#2f#)) OR
 					(reg_q1955 AND symb_decoder(16#ad#)) OR
 					(reg_q1955 AND symb_decoder(16#6a#)) OR
 					(reg_q1955 AND symb_decoder(16#46#)) OR
 					(reg_q1955 AND symb_decoder(16#38#)) OR
 					(reg_q1955 AND symb_decoder(16#52#)) OR
 					(reg_q1955 AND symb_decoder(16#64#)) OR
 					(reg_q1955 AND symb_decoder(16#e6#)) OR
 					(reg_q1955 AND symb_decoder(16#bf#)) OR
 					(reg_q1955 AND symb_decoder(16#a1#)) OR
 					(reg_q1955 AND symb_decoder(16#c0#)) OR
 					(reg_q1955 AND symb_decoder(16#70#)) OR
 					(reg_q1955 AND symb_decoder(16#f5#)) OR
 					(reg_q1955 AND symb_decoder(16#dd#)) OR
 					(reg_q1955 AND symb_decoder(16#41#)) OR
 					(reg_q1955 AND symb_decoder(16#c6#)) OR
 					(reg_q1955 AND symb_decoder(16#45#)) OR
 					(reg_q1955 AND symb_decoder(16#47#)) OR
 					(reg_q1955 AND symb_decoder(16#5a#)) OR
 					(reg_q1955 AND symb_decoder(16#9c#)) OR
 					(reg_q1955 AND symb_decoder(16#cf#)) OR
 					(reg_q1955 AND symb_decoder(16#1b#)) OR
 					(reg_q1955 AND symb_decoder(16#2a#)) OR
 					(reg_q1955 AND symb_decoder(16#84#)) OR
 					(reg_q1955 AND symb_decoder(16#fa#)) OR
 					(reg_q1955 AND symb_decoder(16#a2#)) OR
 					(reg_q1955 AND symb_decoder(16#76#)) OR
 					(reg_q1955 AND symb_decoder(16#9a#)) OR
 					(reg_q1955 AND symb_decoder(16#9e#)) OR
 					(reg_q1955 AND symb_decoder(16#eb#)) OR
 					(reg_q1955 AND symb_decoder(16#8a#)) OR
 					(reg_q1955 AND symb_decoder(16#18#)) OR
 					(reg_q1955 AND symb_decoder(16#99#)) OR
 					(reg_q1955 AND symb_decoder(16#9d#)) OR
 					(reg_q1955 AND symb_decoder(16#7c#)) OR
 					(reg_q1955 AND symb_decoder(16#85#)) OR
 					(reg_q1955 AND symb_decoder(16#ca#)) OR
 					(reg_q1955 AND symb_decoder(16#df#)) OR
 					(reg_q1955 AND symb_decoder(16#07#)) OR
 					(reg_q1955 AND symb_decoder(16#16#)) OR
 					(reg_q1955 AND symb_decoder(16#0a#)) OR
 					(reg_q1955 AND symb_decoder(16#aa#)) OR
 					(reg_q1955 AND symb_decoder(16#15#)) OR
 					(reg_q1955 AND symb_decoder(16#56#)) OR
 					(reg_q1955 AND symb_decoder(16#4d#)) OR
 					(reg_q1955 AND symb_decoder(16#0d#)) OR
 					(reg_q1955 AND symb_decoder(16#e9#)) OR
 					(reg_q1955 AND symb_decoder(16#5f#)) OR
 					(reg_q1955 AND symb_decoder(16#7a#)) OR
 					(reg_q1955 AND symb_decoder(16#7b#)) OR
 					(reg_q1955 AND symb_decoder(16#13#)) OR
 					(reg_q1955 AND symb_decoder(16#c3#)) OR
 					(reg_q1955 AND symb_decoder(16#e0#)) OR
 					(reg_q1955 AND symb_decoder(16#bc#)) OR
 					(reg_q1955 AND symb_decoder(16#f6#)) OR
 					(reg_q1955 AND symb_decoder(16#f4#)) OR
 					(reg_q1955 AND symb_decoder(16#27#)) OR
 					(reg_q1955 AND symb_decoder(16#0c#)) OR
 					(reg_q1955 AND symb_decoder(16#2d#)) OR
 					(reg_q1955 AND symb_decoder(16#db#)) OR
 					(reg_q1955 AND symb_decoder(16#95#)) OR
 					(reg_q1955 AND symb_decoder(16#7e#)) OR
 					(reg_q1955 AND symb_decoder(16#72#)) OR
 					(reg_q1955 AND symb_decoder(16#f7#)) OR
 					(reg_q1955 AND symb_decoder(16#a5#)) OR
 					(reg_q1955 AND symb_decoder(16#50#)) OR
 					(reg_q1955 AND symb_decoder(16#4f#)) OR
 					(reg_q1955 AND symb_decoder(16#a7#)) OR
 					(reg_q1955 AND symb_decoder(16#43#)) OR
 					(reg_q1955 AND symb_decoder(16#f9#)) OR
 					(reg_q1955 AND symb_decoder(16#1c#)) OR
 					(reg_q1955 AND symb_decoder(16#25#)) OR
 					(reg_q1955 AND symb_decoder(16#1e#)) OR
 					(reg_q1955 AND symb_decoder(16#d6#)) OR
 					(reg_q1955 AND symb_decoder(16#73#)) OR
 					(reg_q1955 AND symb_decoder(16#83#)) OR
 					(reg_q1955 AND symb_decoder(16#c4#)) OR
 					(reg_q1955 AND symb_decoder(16#bb#)) OR
 					(reg_q1955 AND symb_decoder(16#40#)) OR
 					(reg_q1955 AND symb_decoder(16#58#)) OR
 					(reg_q1955 AND symb_decoder(16#12#)) OR
 					(reg_q1955 AND symb_decoder(16#5d#)) OR
 					(reg_q1955 AND symb_decoder(16#5e#)) OR
 					(reg_q1955 AND symb_decoder(16#97#)) OR
 					(reg_q1955 AND symb_decoder(16#3d#)) OR
 					(reg_q1955 AND symb_decoder(16#4a#)) OR
 					(reg_q1955 AND symb_decoder(16#2c#)) OR
 					(reg_q1955 AND symb_decoder(16#94#)) OR
 					(reg_q1955 AND symb_decoder(16#02#)) OR
 					(reg_q1955 AND symb_decoder(16#21#)) OR
 					(reg_q1955 AND symb_decoder(16#33#)) OR
 					(reg_q1955 AND symb_decoder(16#82#)) OR
 					(reg_q1955 AND symb_decoder(16#36#)) OR
 					(reg_q1955 AND symb_decoder(16#1d#)) OR
 					(reg_q1955 AND symb_decoder(16#75#)) OR
 					(reg_q1955 AND symb_decoder(16#60#)) OR
 					(reg_q1955 AND symb_decoder(16#80#)) OR
 					(reg_q1955 AND symb_decoder(16#e4#)) OR
 					(reg_q1955 AND symb_decoder(16#04#)) OR
 					(reg_q1955 AND symb_decoder(16#44#)) OR
 					(reg_q1955 AND symb_decoder(16#7f#)) OR
 					(reg_q1955 AND symb_decoder(16#cc#)) OR
 					(reg_q1955 AND symb_decoder(16#0e#)) OR
 					(reg_q1955 AND symb_decoder(16#d1#)) OR
 					(reg_q1955 AND symb_decoder(16#ce#)) OR
 					(reg_q1955 AND symb_decoder(16#b2#)) OR
 					(reg_q1955 AND symb_decoder(16#a4#)) OR
 					(reg_q1955 AND symb_decoder(16#87#)) OR
 					(reg_q1955 AND symb_decoder(16#89#)) OR
 					(reg_q1955 AND symb_decoder(16#81#)) OR
 					(reg_q1955 AND symb_decoder(16#1f#)) OR
 					(reg_q1955 AND symb_decoder(16#19#)) OR
 					(reg_q1955 AND symb_decoder(16#53#)) OR
 					(reg_q1955 AND symb_decoder(16#c1#)) OR
 					(reg_q1955 AND symb_decoder(16#42#)) OR
 					(reg_q1955 AND symb_decoder(16#6f#)) OR
 					(reg_q1955 AND symb_decoder(16#57#)) OR
 					(reg_q1955 AND symb_decoder(16#9b#)) OR
 					(reg_q1955 AND symb_decoder(16#5b#)) OR
 					(reg_q1955 AND symb_decoder(16#91#)) OR
 					(reg_q1955 AND symb_decoder(16#ec#)) OR
 					(reg_q1955 AND symb_decoder(16#34#)) OR
 					(reg_q1955 AND symb_decoder(16#68#)) OR
 					(reg_q1955 AND symb_decoder(16#61#)) OR
 					(reg_q1955 AND symb_decoder(16#00#)) OR
 					(reg_q1955 AND symb_decoder(16#29#)) OR
 					(reg_q1955 AND symb_decoder(16#8e#)) OR
 					(reg_q1955 AND symb_decoder(16#b6#)) OR
 					(reg_q1955 AND symb_decoder(16#cb#)) OR
 					(reg_q1955 AND symb_decoder(16#2b#)) OR
 					(reg_q1955 AND symb_decoder(16#65#)) OR
 					(reg_q1955 AND symb_decoder(16#30#)) OR
 					(reg_q1955 AND symb_decoder(16#55#)) OR
 					(reg_q1955 AND symb_decoder(16#d5#)) OR
 					(reg_q1955 AND symb_decoder(16#28#)) OR
 					(reg_q1955 AND symb_decoder(16#b7#)) OR
 					(reg_q1955 AND symb_decoder(16#b5#)) OR
 					(reg_q1955 AND symb_decoder(16#35#)) OR
 					(reg_q1955 AND symb_decoder(16#c5#)) OR
 					(reg_q1955 AND symb_decoder(16#6c#)) OR
 					(reg_q1955 AND symb_decoder(16#05#)) OR
 					(reg_q1955 AND symb_decoder(16#4b#)) OR
 					(reg_q1955 AND symb_decoder(16#c8#)) OR
 					(reg_q1955 AND symb_decoder(16#bd#)) OR
 					(reg_q1955 AND symb_decoder(16#10#)) OR
 					(reg_q1955 AND symb_decoder(16#ff#)) OR
 					(reg_q1955 AND symb_decoder(16#11#)) OR
 					(reg_q1955 AND symb_decoder(16#0b#)) OR
 					(reg_q1955 AND symb_decoder(16#71#)) OR
 					(reg_q1955 AND symb_decoder(16#e1#)) OR
 					(reg_q1955 AND symb_decoder(16#6b#)) OR
 					(reg_q1955 AND symb_decoder(16#4c#)) OR
 					(reg_q1955 AND symb_decoder(16#3e#)) OR
 					(reg_q1955 AND symb_decoder(16#32#)) OR
 					(reg_q1955 AND symb_decoder(16#93#)) OR
 					(reg_q1955 AND symb_decoder(16#cd#)) OR
 					(reg_q1955 AND symb_decoder(16#54#)) OR
 					(reg_q1955 AND symb_decoder(16#b0#)) OR
 					(reg_q1955 AND symb_decoder(16#96#)) OR
 					(reg_q1955 AND symb_decoder(16#e7#)) OR
 					(reg_q1955 AND symb_decoder(16#6d#)) OR
 					(reg_q1955 AND symb_decoder(16#a8#)) OR
 					(reg_q1955 AND symb_decoder(16#31#)) OR
 					(reg_q1955 AND symb_decoder(16#37#)) OR
 					(reg_q1955 AND symb_decoder(16#6e#)) OR
 					(reg_q1955 AND symb_decoder(16#3c#)) OR
 					(reg_q1955 AND symb_decoder(16#17#)) OR
 					(reg_q1955 AND symb_decoder(16#14#)) OR
 					(reg_q1955 AND symb_decoder(16#8d#)) OR
 					(reg_q1955 AND symb_decoder(16#8b#)) OR
 					(reg_q1955 AND symb_decoder(16#22#)) OR
 					(reg_q1955 AND symb_decoder(16#01#)) OR
 					(reg_q1955 AND symb_decoder(16#fc#)) OR
 					(reg_q1955 AND symb_decoder(16#26#)) OR
 					(reg_q1955 AND symb_decoder(16#fe#)) OR
 					(reg_q1955 AND symb_decoder(16#62#)) OR
 					(reg_q1955 AND symb_decoder(16#f2#)) OR
 					(reg_q1955 AND symb_decoder(16#66#)) OR
 					(reg_q1955 AND symb_decoder(16#3a#)) OR
 					(reg_q1955 AND symb_decoder(16#88#)) OR
 					(reg_q1955 AND symb_decoder(16#09#)) OR
 					(reg_q1955 AND symb_decoder(16#ef#)) OR
 					(reg_q1955 AND symb_decoder(16#24#)) OR
 					(reg_q1955 AND symb_decoder(16#20#)) OR
 					(reg_q1955 AND symb_decoder(16#fd#)) OR
 					(reg_q1955 AND symb_decoder(16#4e#)) OR
 					(reg_q1955 AND symb_decoder(16#92#)) OR
 					(reg_q1955 AND symb_decoder(16#90#)) OR
 					(reg_q1955 AND symb_decoder(16#67#)) OR
 					(reg_q1955 AND symb_decoder(16#8c#)) OR
 					(reg_q1955 AND symb_decoder(16#b4#)) OR
 					(reg_q1955 AND symb_decoder(16#dc#)) OR
 					(reg_q1955 AND symb_decoder(16#ae#)) OR
 					(reg_q1955 AND symb_decoder(16#98#)) OR
 					(reg_q1955 AND symb_decoder(16#f0#));
reg_q1955_init <= '0' ;
	p_reg_q1955: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1955 <= reg_q1955_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1955 <= reg_q1955_init;
        else
          reg_q1955 <= reg_q1955_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q262_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q262 AND symb_decoder(16#89#)) OR
 					(reg_q262 AND symb_decoder(16#fa#)) OR
 					(reg_q262 AND symb_decoder(16#55#)) OR
 					(reg_q262 AND symb_decoder(16#01#)) OR
 					(reg_q262 AND symb_decoder(16#a0#)) OR
 					(reg_q262 AND symb_decoder(16#b4#)) OR
 					(reg_q262 AND symb_decoder(16#08#)) OR
 					(reg_q262 AND symb_decoder(16#ba#)) OR
 					(reg_q262 AND symb_decoder(16#6f#)) OR
 					(reg_q262 AND symb_decoder(16#b1#)) OR
 					(reg_q262 AND symb_decoder(16#70#)) OR
 					(reg_q262 AND symb_decoder(16#db#)) OR
 					(reg_q262 AND symb_decoder(16#64#)) OR
 					(reg_q262 AND symb_decoder(16#b9#)) OR
 					(reg_q262 AND symb_decoder(16#22#)) OR
 					(reg_q262 AND symb_decoder(16#96#)) OR
 					(reg_q262 AND symb_decoder(16#c4#)) OR
 					(reg_q262 AND symb_decoder(16#e2#)) OR
 					(reg_q262 AND symb_decoder(16#27#)) OR
 					(reg_q262 AND symb_decoder(16#3d#)) OR
 					(reg_q262 AND symb_decoder(16#dc#)) OR
 					(reg_q262 AND symb_decoder(16#06#)) OR
 					(reg_q262 AND symb_decoder(16#2b#)) OR
 					(reg_q262 AND symb_decoder(16#da#)) OR
 					(reg_q262 AND symb_decoder(16#78#)) OR
 					(reg_q262 AND symb_decoder(16#49#)) OR
 					(reg_q262 AND symb_decoder(16#04#)) OR
 					(reg_q262 AND symb_decoder(16#88#)) OR
 					(reg_q262 AND symb_decoder(16#30#)) OR
 					(reg_q262 AND symb_decoder(16#2f#)) OR
 					(reg_q262 AND symb_decoder(16#f4#)) OR
 					(reg_q262 AND symb_decoder(16#95#)) OR
 					(reg_q262 AND symb_decoder(16#be#)) OR
 					(reg_q262 AND symb_decoder(16#83#)) OR
 					(reg_q262 AND symb_decoder(16#42#)) OR
 					(reg_q262 AND symb_decoder(16#f9#)) OR
 					(reg_q262 AND symb_decoder(16#35#)) OR
 					(reg_q262 AND symb_decoder(16#f8#)) OR
 					(reg_q262 AND symb_decoder(16#fb#)) OR
 					(reg_q262 AND symb_decoder(16#d9#)) OR
 					(reg_q262 AND symb_decoder(16#a9#)) OR
 					(reg_q262 AND symb_decoder(16#a1#)) OR
 					(reg_q262 AND symb_decoder(16#2d#)) OR
 					(reg_q262 AND symb_decoder(16#69#)) OR
 					(reg_q262 AND symb_decoder(16#36#)) OR
 					(reg_q262 AND symb_decoder(16#a3#)) OR
 					(reg_q262 AND symb_decoder(16#ec#)) OR
 					(reg_q262 AND symb_decoder(16#c6#)) OR
 					(reg_q262 AND symb_decoder(16#13#)) OR
 					(reg_q262 AND symb_decoder(16#c8#)) OR
 					(reg_q262 AND symb_decoder(16#3c#)) OR
 					(reg_q262 AND symb_decoder(16#b0#)) OR
 					(reg_q262 AND symb_decoder(16#71#)) OR
 					(reg_q262 AND symb_decoder(16#7c#)) OR
 					(reg_q262 AND symb_decoder(16#59#)) OR
 					(reg_q262 AND symb_decoder(16#38#)) OR
 					(reg_q262 AND symb_decoder(16#10#)) OR
 					(reg_q262 AND symb_decoder(16#29#)) OR
 					(reg_q262 AND symb_decoder(16#39#)) OR
 					(reg_q262 AND symb_decoder(16#12#)) OR
 					(reg_q262 AND symb_decoder(16#ea#)) OR
 					(reg_q262 AND symb_decoder(16#7e#)) OR
 					(reg_q262 AND symb_decoder(16#8c#)) OR
 					(reg_q262 AND symb_decoder(16#fd#)) OR
 					(reg_q262 AND symb_decoder(16#5c#)) OR
 					(reg_q262 AND symb_decoder(16#3e#)) OR
 					(reg_q262 AND symb_decoder(16#19#)) OR
 					(reg_q262 AND symb_decoder(16#9b#)) OR
 					(reg_q262 AND symb_decoder(16#34#)) OR
 					(reg_q262 AND symb_decoder(16#07#)) OR
 					(reg_q262 AND symb_decoder(16#5d#)) OR
 					(reg_q262 AND symb_decoder(16#9a#)) OR
 					(reg_q262 AND symb_decoder(16#dd#)) OR
 					(reg_q262 AND symb_decoder(16#e9#)) OR
 					(reg_q262 AND symb_decoder(16#76#)) OR
 					(reg_q262 AND symb_decoder(16#ac#)) OR
 					(reg_q262 AND symb_decoder(16#7a#)) OR
 					(reg_q262 AND symb_decoder(16#e4#)) OR
 					(reg_q262 AND symb_decoder(16#41#)) OR
 					(reg_q262 AND symb_decoder(16#eb#)) OR
 					(reg_q262 AND symb_decoder(16#50#)) OR
 					(reg_q262 AND symb_decoder(16#48#)) OR
 					(reg_q262 AND symb_decoder(16#d8#)) OR
 					(reg_q262 AND symb_decoder(16#de#)) OR
 					(reg_q262 AND symb_decoder(16#e3#)) OR
 					(reg_q262 AND symb_decoder(16#0a#)) OR
 					(reg_q262 AND symb_decoder(16#03#)) OR
 					(reg_q262 AND symb_decoder(16#e0#)) OR
 					(reg_q262 AND symb_decoder(16#23#)) OR
 					(reg_q262 AND symb_decoder(16#9d#)) OR
 					(reg_q262 AND symb_decoder(16#09#)) OR
 					(reg_q262 AND symb_decoder(16#e7#)) OR
 					(reg_q262 AND symb_decoder(16#f1#)) OR
 					(reg_q262 AND symb_decoder(16#7f#)) OR
 					(reg_q262 AND symb_decoder(16#9f#)) OR
 					(reg_q262 AND symb_decoder(16#c3#)) OR
 					(reg_q262 AND symb_decoder(16#6e#)) OR
 					(reg_q262 AND symb_decoder(16#65#)) OR
 					(reg_q262 AND symb_decoder(16#3b#)) OR
 					(reg_q262 AND symb_decoder(16#16#)) OR
 					(reg_q262 AND symb_decoder(16#ca#)) OR
 					(reg_q262 AND symb_decoder(16#14#)) OR
 					(reg_q262 AND symb_decoder(16#bc#)) OR
 					(reg_q262 AND symb_decoder(16#ab#)) OR
 					(reg_q262 AND symb_decoder(16#5e#)) OR
 					(reg_q262 AND symb_decoder(16#20#)) OR
 					(reg_q262 AND symb_decoder(16#3f#)) OR
 					(reg_q262 AND symb_decoder(16#1f#)) OR
 					(reg_q262 AND symb_decoder(16#82#)) OR
 					(reg_q262 AND symb_decoder(16#a7#)) OR
 					(reg_q262 AND symb_decoder(16#02#)) OR
 					(reg_q262 AND symb_decoder(16#40#)) OR
 					(reg_q262 AND symb_decoder(16#72#)) OR
 					(reg_q262 AND symb_decoder(16#60#)) OR
 					(reg_q262 AND symb_decoder(16#fe#)) OR
 					(reg_q262 AND symb_decoder(16#ef#)) OR
 					(reg_q262 AND symb_decoder(16#4c#)) OR
 					(reg_q262 AND symb_decoder(16#92#)) OR
 					(reg_q262 AND symb_decoder(16#a6#)) OR
 					(reg_q262 AND symb_decoder(16#6b#)) OR
 					(reg_q262 AND symb_decoder(16#fc#)) OR
 					(reg_q262 AND symb_decoder(16#1b#)) OR
 					(reg_q262 AND symb_decoder(16#94#)) OR
 					(reg_q262 AND symb_decoder(16#8e#)) OR
 					(reg_q262 AND symb_decoder(16#85#)) OR
 					(reg_q262 AND symb_decoder(16#aa#)) OR
 					(reg_q262 AND symb_decoder(16#81#)) OR
 					(reg_q262 AND symb_decoder(16#8f#)) OR
 					(reg_q262 AND symb_decoder(16#24#)) OR
 					(reg_q262 AND symb_decoder(16#8b#)) OR
 					(reg_q262 AND symb_decoder(16#d4#)) OR
 					(reg_q262 AND symb_decoder(16#4d#)) OR
 					(reg_q262 AND symb_decoder(16#bb#)) OR
 					(reg_q262 AND symb_decoder(16#0b#)) OR
 					(reg_q262 AND symb_decoder(16#0d#)) OR
 					(reg_q262 AND symb_decoder(16#e1#)) OR
 					(reg_q262 AND symb_decoder(16#21#)) OR
 					(reg_q262 AND symb_decoder(16#b5#)) OR
 					(reg_q262 AND symb_decoder(16#d5#)) OR
 					(reg_q262 AND symb_decoder(16#d2#)) OR
 					(reg_q262 AND symb_decoder(16#e8#)) OR
 					(reg_q262 AND symb_decoder(16#4e#)) OR
 					(reg_q262 AND symb_decoder(16#1c#)) OR
 					(reg_q262 AND symb_decoder(16#90#)) OR
 					(reg_q262 AND symb_decoder(16#62#)) OR
 					(reg_q262 AND symb_decoder(16#a4#)) OR
 					(reg_q262 AND symb_decoder(16#0f#)) OR
 					(reg_q262 AND symb_decoder(16#c1#)) OR
 					(reg_q262 AND symb_decoder(16#33#)) OR
 					(reg_q262 AND symb_decoder(16#56#)) OR
 					(reg_q262 AND symb_decoder(16#57#)) OR
 					(reg_q262 AND symb_decoder(16#b6#)) OR
 					(reg_q262 AND symb_decoder(16#87#)) OR
 					(reg_q262 AND symb_decoder(16#c7#)) OR
 					(reg_q262 AND symb_decoder(16#8a#)) OR
 					(reg_q262 AND symb_decoder(16#ae#)) OR
 					(reg_q262 AND symb_decoder(16#f2#)) OR
 					(reg_q262 AND symb_decoder(16#15#)) OR
 					(reg_q262 AND symb_decoder(16#ad#)) OR
 					(reg_q262 AND symb_decoder(16#b3#)) OR
 					(reg_q262 AND symb_decoder(16#84#)) OR
 					(reg_q262 AND symb_decoder(16#2c#)) OR
 					(reg_q262 AND symb_decoder(16#ff#)) OR
 					(reg_q262 AND symb_decoder(16#4a#)) OR
 					(reg_q262 AND symb_decoder(16#5a#)) OR
 					(reg_q262 AND symb_decoder(16#ce#)) OR
 					(reg_q262 AND symb_decoder(16#91#)) OR
 					(reg_q262 AND symb_decoder(16#1d#)) OR
 					(reg_q262 AND symb_decoder(16#31#)) OR
 					(reg_q262 AND symb_decoder(16#c0#)) OR
 					(reg_q262 AND symb_decoder(16#f3#)) OR
 					(reg_q262 AND symb_decoder(16#ee#)) OR
 					(reg_q262 AND symb_decoder(16#67#)) OR
 					(reg_q262 AND symb_decoder(16#cd#)) OR
 					(reg_q262 AND symb_decoder(16#54#)) OR
 					(reg_q262 AND symb_decoder(16#b7#)) OR
 					(reg_q262 AND symb_decoder(16#00#)) OR
 					(reg_q262 AND symb_decoder(16#a2#)) OR
 					(reg_q262 AND symb_decoder(16#73#)) OR
 					(reg_q262 AND symb_decoder(16#c5#)) OR
 					(reg_q262 AND symb_decoder(16#99#)) OR
 					(reg_q262 AND symb_decoder(16#cc#)) OR
 					(reg_q262 AND symb_decoder(16#c2#)) OR
 					(reg_q262 AND symb_decoder(16#d6#)) OR
 					(reg_q262 AND symb_decoder(16#ed#)) OR
 					(reg_q262 AND symb_decoder(16#17#)) OR
 					(reg_q262 AND symb_decoder(16#b8#)) OR
 					(reg_q262 AND symb_decoder(16#44#)) OR
 					(reg_q262 AND symb_decoder(16#f0#)) OR
 					(reg_q262 AND symb_decoder(16#37#)) OR
 					(reg_q262 AND symb_decoder(16#df#)) OR
 					(reg_q262 AND symb_decoder(16#93#)) OR
 					(reg_q262 AND symb_decoder(16#9c#)) OR
 					(reg_q262 AND symb_decoder(16#c9#)) OR
 					(reg_q262 AND symb_decoder(16#e6#)) OR
 					(reg_q262 AND symb_decoder(16#58#)) OR
 					(reg_q262 AND symb_decoder(16#86#)) OR
 					(reg_q262 AND symb_decoder(16#0e#)) OR
 					(reg_q262 AND symb_decoder(16#79#)) OR
 					(reg_q262 AND symb_decoder(16#43#)) OR
 					(reg_q262 AND symb_decoder(16#f6#)) OR
 					(reg_q262 AND symb_decoder(16#6c#)) OR
 					(reg_q262 AND symb_decoder(16#11#)) OR
 					(reg_q262 AND symb_decoder(16#97#)) OR
 					(reg_q262 AND symb_decoder(16#05#)) OR
 					(reg_q262 AND symb_decoder(16#7d#)) OR
 					(reg_q262 AND symb_decoder(16#32#)) OR
 					(reg_q262 AND symb_decoder(16#47#)) OR
 					(reg_q262 AND symb_decoder(16#80#)) OR
 					(reg_q262 AND symb_decoder(16#7b#)) OR
 					(reg_q262 AND symb_decoder(16#5b#)) OR
 					(reg_q262 AND symb_decoder(16#4f#)) OR
 					(reg_q262 AND symb_decoder(16#cb#)) OR
 					(reg_q262 AND symb_decoder(16#8d#)) OR
 					(reg_q262 AND symb_decoder(16#25#)) OR
 					(reg_q262 AND symb_decoder(16#45#)) OR
 					(reg_q262 AND symb_decoder(16#a5#)) OR
 					(reg_q262 AND symb_decoder(16#b2#)) OR
 					(reg_q262 AND symb_decoder(16#a8#)) OR
 					(reg_q262 AND symb_decoder(16#f7#)) OR
 					(reg_q262 AND symb_decoder(16#1a#)) OR
 					(reg_q262 AND symb_decoder(16#98#)) OR
 					(reg_q262 AND symb_decoder(16#e5#)) OR
 					(reg_q262 AND symb_decoder(16#4b#)) OR
 					(reg_q262 AND symb_decoder(16#cf#)) OR
 					(reg_q262 AND symb_decoder(16#6a#)) OR
 					(reg_q262 AND symb_decoder(16#66#)) OR
 					(reg_q262 AND symb_decoder(16#d1#)) OR
 					(reg_q262 AND symb_decoder(16#d3#)) OR
 					(reg_q262 AND symb_decoder(16#6d#)) OR
 					(reg_q262 AND symb_decoder(16#28#)) OR
 					(reg_q262 AND symb_decoder(16#46#)) OR
 					(reg_q262 AND symb_decoder(16#1e#)) OR
 					(reg_q262 AND symb_decoder(16#51#)) OR
 					(reg_q262 AND symb_decoder(16#0c#)) OR
 					(reg_q262 AND symb_decoder(16#26#)) OR
 					(reg_q262 AND symb_decoder(16#52#)) OR
 					(reg_q262 AND symb_decoder(16#74#)) OR
 					(reg_q262 AND symb_decoder(16#18#)) OR
 					(reg_q262 AND symb_decoder(16#61#)) OR
 					(reg_q262 AND symb_decoder(16#f5#)) OR
 					(reg_q262 AND symb_decoder(16#bd#)) OR
 					(reg_q262 AND symb_decoder(16#d0#)) OR
 					(reg_q262 AND symb_decoder(16#bf#)) OR
 					(reg_q262 AND symb_decoder(16#5f#)) OR
 					(reg_q262 AND symb_decoder(16#d7#)) OR
 					(reg_q262 AND symb_decoder(16#68#)) OR
 					(reg_q262 AND symb_decoder(16#3a#)) OR
 					(reg_q262 AND symb_decoder(16#2a#)) OR
 					(reg_q262 AND symb_decoder(16#2e#)) OR
 					(reg_q262 AND symb_decoder(16#77#)) OR
 					(reg_q262 AND symb_decoder(16#53#)) OR
 					(reg_q262 AND symb_decoder(16#9e#)) OR
 					(reg_q262 AND symb_decoder(16#af#)) OR
 					(reg_q262 AND symb_decoder(16#75#)) OR
 					(reg_q262 AND symb_decoder(16#63#));
reg_q262_init <= '0' ;
	p_reg_q262: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q262 <= reg_q262_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q262 <= reg_q262_init;
        else
          reg_q262 <= reg_q262_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q958_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q958 AND symb_decoder(16#a4#)) OR
 					(reg_q958 AND symb_decoder(16#4c#)) OR
 					(reg_q958 AND symb_decoder(16#e3#)) OR
 					(reg_q958 AND symb_decoder(16#83#)) OR
 					(reg_q958 AND symb_decoder(16#4e#)) OR
 					(reg_q958 AND symb_decoder(16#26#)) OR
 					(reg_q958 AND symb_decoder(16#39#)) OR
 					(reg_q958 AND symb_decoder(16#04#)) OR
 					(reg_q958 AND symb_decoder(16#70#)) OR
 					(reg_q958 AND symb_decoder(16#20#)) OR
 					(reg_q958 AND symb_decoder(16#8c#)) OR
 					(reg_q958 AND symb_decoder(16#43#)) OR
 					(reg_q958 AND symb_decoder(16#87#)) OR
 					(reg_q958 AND symb_decoder(16#ac#)) OR
 					(reg_q958 AND symb_decoder(16#0a#)) OR
 					(reg_q958 AND symb_decoder(16#ba#)) OR
 					(reg_q958 AND symb_decoder(16#ee#)) OR
 					(reg_q958 AND symb_decoder(16#0e#)) OR
 					(reg_q958 AND symb_decoder(16#01#)) OR
 					(reg_q958 AND symb_decoder(16#d6#)) OR
 					(reg_q958 AND symb_decoder(16#00#)) OR
 					(reg_q958 AND symb_decoder(16#40#)) OR
 					(reg_q958 AND symb_decoder(16#1f#)) OR
 					(reg_q958 AND symb_decoder(16#8f#)) OR
 					(reg_q958 AND symb_decoder(16#af#)) OR
 					(reg_q958 AND symb_decoder(16#a8#)) OR
 					(reg_q958 AND symb_decoder(16#e4#)) OR
 					(reg_q958 AND symb_decoder(16#55#)) OR
 					(reg_q958 AND symb_decoder(16#f4#)) OR
 					(reg_q958 AND symb_decoder(16#34#)) OR
 					(reg_q958 AND symb_decoder(16#54#)) OR
 					(reg_q958 AND symb_decoder(16#cd#)) OR
 					(reg_q958 AND symb_decoder(16#ec#)) OR
 					(reg_q958 AND symb_decoder(16#79#)) OR
 					(reg_q958 AND symb_decoder(16#8a#)) OR
 					(reg_q958 AND symb_decoder(16#80#)) OR
 					(reg_q958 AND symb_decoder(16#6f#)) OR
 					(reg_q958 AND symb_decoder(16#09#)) OR
 					(reg_q958 AND symb_decoder(16#46#)) OR
 					(reg_q958 AND symb_decoder(16#ef#)) OR
 					(reg_q958 AND symb_decoder(16#a5#)) OR
 					(reg_q958 AND symb_decoder(16#31#)) OR
 					(reg_q958 AND symb_decoder(16#42#)) OR
 					(reg_q958 AND symb_decoder(16#fe#)) OR
 					(reg_q958 AND symb_decoder(16#e5#)) OR
 					(reg_q958 AND symb_decoder(16#49#)) OR
 					(reg_q958 AND symb_decoder(16#65#)) OR
 					(reg_q958 AND symb_decoder(16#13#)) OR
 					(reg_q958 AND symb_decoder(16#06#)) OR
 					(reg_q958 AND symb_decoder(16#82#)) OR
 					(reg_q958 AND symb_decoder(16#0b#)) OR
 					(reg_q958 AND symb_decoder(16#ab#)) OR
 					(reg_q958 AND symb_decoder(16#02#)) OR
 					(reg_q958 AND symb_decoder(16#5b#)) OR
 					(reg_q958 AND symb_decoder(16#cf#)) OR
 					(reg_q958 AND symb_decoder(16#3a#)) OR
 					(reg_q958 AND symb_decoder(16#84#)) OR
 					(reg_q958 AND symb_decoder(16#52#)) OR
 					(reg_q958 AND symb_decoder(16#da#)) OR
 					(reg_q958 AND symb_decoder(16#7a#)) OR
 					(reg_q958 AND symb_decoder(16#ce#)) OR
 					(reg_q958 AND symb_decoder(16#a9#)) OR
 					(reg_q958 AND symb_decoder(16#69#)) OR
 					(reg_q958 AND symb_decoder(16#c6#)) OR
 					(reg_q958 AND symb_decoder(16#91#)) OR
 					(reg_q958 AND symb_decoder(16#05#)) OR
 					(reg_q958 AND symb_decoder(16#95#)) OR
 					(reg_q958 AND symb_decoder(16#c7#)) OR
 					(reg_q958 AND symb_decoder(16#6d#)) OR
 					(reg_q958 AND symb_decoder(16#76#)) OR
 					(reg_q958 AND symb_decoder(16#a0#)) OR
 					(reg_q958 AND symb_decoder(16#2c#)) OR
 					(reg_q958 AND symb_decoder(16#72#)) OR
 					(reg_q958 AND symb_decoder(16#60#)) OR
 					(reg_q958 AND symb_decoder(16#74#)) OR
 					(reg_q958 AND symb_decoder(16#fd#)) OR
 					(reg_q958 AND symb_decoder(16#38#)) OR
 					(reg_q958 AND symb_decoder(16#35#)) OR
 					(reg_q958 AND symb_decoder(16#86#)) OR
 					(reg_q958 AND symb_decoder(16#c0#)) OR
 					(reg_q958 AND symb_decoder(16#fc#)) OR
 					(reg_q958 AND symb_decoder(16#29#)) OR
 					(reg_q958 AND symb_decoder(16#4b#)) OR
 					(reg_q958 AND symb_decoder(16#1a#)) OR
 					(reg_q958 AND symb_decoder(16#ea#)) OR
 					(reg_q958 AND symb_decoder(16#b3#)) OR
 					(reg_q958 AND symb_decoder(16#ed#)) OR
 					(reg_q958 AND symb_decoder(16#5a#)) OR
 					(reg_q958 AND symb_decoder(16#1d#)) OR
 					(reg_q958 AND symb_decoder(16#f1#)) OR
 					(reg_q958 AND symb_decoder(16#aa#)) OR
 					(reg_q958 AND symb_decoder(16#b9#)) OR
 					(reg_q958 AND symb_decoder(16#cb#)) OR
 					(reg_q958 AND symb_decoder(16#a1#)) OR
 					(reg_q958 AND symb_decoder(16#3c#)) OR
 					(reg_q958 AND symb_decoder(16#18#)) OR
 					(reg_q958 AND symb_decoder(16#77#)) OR
 					(reg_q958 AND symb_decoder(16#53#)) OR
 					(reg_q958 AND symb_decoder(16#88#)) OR
 					(reg_q958 AND symb_decoder(16#50#)) OR
 					(reg_q958 AND symb_decoder(16#bc#)) OR
 					(reg_q958 AND symb_decoder(16#32#)) OR
 					(reg_q958 AND symb_decoder(16#07#)) OR
 					(reg_q958 AND symb_decoder(16#1e#)) OR
 					(reg_q958 AND symb_decoder(16#81#)) OR
 					(reg_q958 AND symb_decoder(16#7b#)) OR
 					(reg_q958 AND symb_decoder(16#9e#)) OR
 					(reg_q958 AND symb_decoder(16#c8#)) OR
 					(reg_q958 AND symb_decoder(16#92#)) OR
 					(reg_q958 AND symb_decoder(16#b5#)) OR
 					(reg_q958 AND symb_decoder(16#2d#)) OR
 					(reg_q958 AND symb_decoder(16#90#)) OR
 					(reg_q958 AND symb_decoder(16#bd#)) OR
 					(reg_q958 AND symb_decoder(16#85#)) OR
 					(reg_q958 AND symb_decoder(16#44#)) OR
 					(reg_q958 AND symb_decoder(16#15#)) OR
 					(reg_q958 AND symb_decoder(16#23#)) OR
 					(reg_q958 AND symb_decoder(16#d7#)) OR
 					(reg_q958 AND symb_decoder(16#37#)) OR
 					(reg_q958 AND symb_decoder(16#16#)) OR
 					(reg_q958 AND symb_decoder(16#45#)) OR
 					(reg_q958 AND symb_decoder(16#dd#)) OR
 					(reg_q958 AND symb_decoder(16#b1#)) OR
 					(reg_q958 AND symb_decoder(16#c5#)) OR
 					(reg_q958 AND symb_decoder(16#5d#)) OR
 					(reg_q958 AND symb_decoder(16#b7#)) OR
 					(reg_q958 AND symb_decoder(16#03#)) OR
 					(reg_q958 AND symb_decoder(16#f6#)) OR
 					(reg_q958 AND symb_decoder(16#a2#)) OR
 					(reg_q958 AND symb_decoder(16#41#)) OR
 					(reg_q958 AND symb_decoder(16#b4#)) OR
 					(reg_q958 AND symb_decoder(16#bb#)) OR
 					(reg_q958 AND symb_decoder(16#9a#)) OR
 					(reg_q958 AND symb_decoder(16#3d#)) OR
 					(reg_q958 AND symb_decoder(16#96#)) OR
 					(reg_q958 AND symb_decoder(16#66#)) OR
 					(reg_q958 AND symb_decoder(16#59#)) OR
 					(reg_q958 AND symb_decoder(16#e7#)) OR
 					(reg_q958 AND symb_decoder(16#10#)) OR
 					(reg_q958 AND symb_decoder(16#3f#)) OR
 					(reg_q958 AND symb_decoder(16#f0#)) OR
 					(reg_q958 AND symb_decoder(16#0d#)) OR
 					(reg_q958 AND symb_decoder(16#36#)) OR
 					(reg_q958 AND symb_decoder(16#97#)) OR
 					(reg_q958 AND symb_decoder(16#e8#)) OR
 					(reg_q958 AND symb_decoder(16#11#)) OR
 					(reg_q958 AND symb_decoder(16#9c#)) OR
 					(reg_q958 AND symb_decoder(16#8d#)) OR
 					(reg_q958 AND symb_decoder(16#93#)) OR
 					(reg_q958 AND symb_decoder(16#58#)) OR
 					(reg_q958 AND symb_decoder(16#56#)) OR
 					(reg_q958 AND symb_decoder(16#75#)) OR
 					(reg_q958 AND symb_decoder(16#bf#)) OR
 					(reg_q958 AND symb_decoder(16#1b#)) OR
 					(reg_q958 AND symb_decoder(16#99#)) OR
 					(reg_q958 AND symb_decoder(16#4a#)) OR
 					(reg_q958 AND symb_decoder(16#e9#)) OR
 					(reg_q958 AND symb_decoder(16#57#)) OR
 					(reg_q958 AND symb_decoder(16#9d#)) OR
 					(reg_q958 AND symb_decoder(16#14#)) OR
 					(reg_q958 AND symb_decoder(16#6a#)) OR
 					(reg_q958 AND symb_decoder(16#7d#)) OR
 					(reg_q958 AND symb_decoder(16#e0#)) OR
 					(reg_q958 AND symb_decoder(16#c9#)) OR
 					(reg_q958 AND symb_decoder(16#8b#)) OR
 					(reg_q958 AND symb_decoder(16#47#)) OR
 					(reg_q958 AND symb_decoder(16#0c#)) OR
 					(reg_q958 AND symb_decoder(16#89#)) OR
 					(reg_q958 AND symb_decoder(16#d2#)) OR
 					(reg_q958 AND symb_decoder(16#a3#)) OR
 					(reg_q958 AND symb_decoder(16#d5#)) OR
 					(reg_q958 AND symb_decoder(16#fa#)) OR
 					(reg_q958 AND symb_decoder(16#d3#)) OR
 					(reg_q958 AND symb_decoder(16#8e#)) OR
 					(reg_q958 AND symb_decoder(16#f9#)) OR
 					(reg_q958 AND symb_decoder(16#21#)) OR
 					(reg_q958 AND symb_decoder(16#4d#)) OR
 					(reg_q958 AND symb_decoder(16#df#)) OR
 					(reg_q958 AND symb_decoder(16#68#)) OR
 					(reg_q958 AND symb_decoder(16#b0#)) OR
 					(reg_q958 AND symb_decoder(16#eb#)) OR
 					(reg_q958 AND symb_decoder(16#3b#)) OR
 					(reg_q958 AND symb_decoder(16#7e#)) OR
 					(reg_q958 AND symb_decoder(16#c2#)) OR
 					(reg_q958 AND symb_decoder(16#d1#)) OR
 					(reg_q958 AND symb_decoder(16#17#)) OR
 					(reg_q958 AND symb_decoder(16#f8#)) OR
 					(reg_q958 AND symb_decoder(16#e1#)) OR
 					(reg_q958 AND symb_decoder(16#67#)) OR
 					(reg_q958 AND symb_decoder(16#6b#)) OR
 					(reg_q958 AND symb_decoder(16#ff#)) OR
 					(reg_q958 AND symb_decoder(16#12#)) OR
 					(reg_q958 AND symb_decoder(16#61#)) OR
 					(reg_q958 AND symb_decoder(16#a7#)) OR
 					(reg_q958 AND symb_decoder(16#19#)) OR
 					(reg_q958 AND symb_decoder(16#be#)) OR
 					(reg_q958 AND symb_decoder(16#28#)) OR
 					(reg_q958 AND symb_decoder(16#71#)) OR
 					(reg_q958 AND symb_decoder(16#e6#)) OR
 					(reg_q958 AND symb_decoder(16#5f#)) OR
 					(reg_q958 AND symb_decoder(16#64#)) OR
 					(reg_q958 AND symb_decoder(16#b6#)) OR
 					(reg_q958 AND symb_decoder(16#f2#)) OR
 					(reg_q958 AND symb_decoder(16#63#)) OR
 					(reg_q958 AND symb_decoder(16#73#)) OR
 					(reg_q958 AND symb_decoder(16#ae#)) OR
 					(reg_q958 AND symb_decoder(16#ca#)) OR
 					(reg_q958 AND symb_decoder(16#48#)) OR
 					(reg_q958 AND symb_decoder(16#d0#)) OR
 					(reg_q958 AND symb_decoder(16#ad#)) OR
 					(reg_q958 AND symb_decoder(16#f7#)) OR
 					(reg_q958 AND symb_decoder(16#c4#)) OR
 					(reg_q958 AND symb_decoder(16#dc#)) OR
 					(reg_q958 AND symb_decoder(16#24#)) OR
 					(reg_q958 AND symb_decoder(16#5c#)) OR
 					(reg_q958 AND symb_decoder(16#f5#)) OR
 					(reg_q958 AND symb_decoder(16#27#)) OR
 					(reg_q958 AND symb_decoder(16#c1#)) OR
 					(reg_q958 AND symb_decoder(16#08#)) OR
 					(reg_q958 AND symb_decoder(16#1c#)) OR
 					(reg_q958 AND symb_decoder(16#5e#)) OR
 					(reg_q958 AND symb_decoder(16#3e#)) OR
 					(reg_q958 AND symb_decoder(16#2e#)) OR
 					(reg_q958 AND symb_decoder(16#6e#)) OR
 					(reg_q958 AND symb_decoder(16#0f#)) OR
 					(reg_q958 AND symb_decoder(16#22#)) OR
 					(reg_q958 AND symb_decoder(16#7f#)) OR
 					(reg_q958 AND symb_decoder(16#2b#)) OR
 					(reg_q958 AND symb_decoder(16#94#)) OR
 					(reg_q958 AND symb_decoder(16#cc#)) OR
 					(reg_q958 AND symb_decoder(16#c3#)) OR
 					(reg_q958 AND symb_decoder(16#de#)) OR
 					(reg_q958 AND symb_decoder(16#b8#)) OR
 					(reg_q958 AND symb_decoder(16#d8#)) OR
 					(reg_q958 AND symb_decoder(16#9f#)) OR
 					(reg_q958 AND symb_decoder(16#98#)) OR
 					(reg_q958 AND symb_decoder(16#fb#)) OR
 					(reg_q958 AND symb_decoder(16#30#)) OR
 					(reg_q958 AND symb_decoder(16#78#)) OR
 					(reg_q958 AND symb_decoder(16#9b#)) OR
 					(reg_q958 AND symb_decoder(16#2f#)) OR
 					(reg_q958 AND symb_decoder(16#d9#)) OR
 					(reg_q958 AND symb_decoder(16#2a#)) OR
 					(reg_q958 AND symb_decoder(16#b2#)) OR
 					(reg_q958 AND symb_decoder(16#e2#)) OR
 					(reg_q958 AND symb_decoder(16#f3#)) OR
 					(reg_q958 AND symb_decoder(16#4f#)) OR
 					(reg_q958 AND symb_decoder(16#25#)) OR
 					(reg_q958 AND symb_decoder(16#62#)) OR
 					(reg_q958 AND symb_decoder(16#33#)) OR
 					(reg_q958 AND symb_decoder(16#a6#)) OR
 					(reg_q958 AND symb_decoder(16#d4#)) OR
 					(reg_q958 AND symb_decoder(16#51#)) OR
 					(reg_q958 AND symb_decoder(16#6c#)) OR
 					(reg_q958 AND symb_decoder(16#db#)) OR
 					(reg_q958 AND symb_decoder(16#7c#));
reg_q958_init <= '0' ;
	p_reg_q958: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q958 <= reg_q958_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q958 <= reg_q958_init;
        else
          reg_q958 <= reg_q958_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q816_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q816 AND symb_decoder(16#4c#)) OR
 					(reg_q816 AND symb_decoder(16#cb#)) OR
 					(reg_q816 AND symb_decoder(16#dd#)) OR
 					(reg_q816 AND symb_decoder(16#3a#)) OR
 					(reg_q816 AND symb_decoder(16#16#)) OR
 					(reg_q816 AND symb_decoder(16#77#)) OR
 					(reg_q816 AND symb_decoder(16#04#)) OR
 					(reg_q816 AND symb_decoder(16#39#)) OR
 					(reg_q816 AND symb_decoder(16#aa#)) OR
 					(reg_q816 AND symb_decoder(16#8e#)) OR
 					(reg_q816 AND symb_decoder(16#93#)) OR
 					(reg_q816 AND symb_decoder(16#05#)) OR
 					(reg_q816 AND symb_decoder(16#0b#)) OR
 					(reg_q816 AND symb_decoder(16#6d#)) OR
 					(reg_q816 AND symb_decoder(16#68#)) OR
 					(reg_q816 AND symb_decoder(16#d4#)) OR
 					(reg_q816 AND symb_decoder(16#9f#)) OR
 					(reg_q816 AND symb_decoder(16#14#)) OR
 					(reg_q816 AND symb_decoder(16#75#)) OR
 					(reg_q816 AND symb_decoder(16#2d#)) OR
 					(reg_q816 AND symb_decoder(16#8f#)) OR
 					(reg_q816 AND symb_decoder(16#42#)) OR
 					(reg_q816 AND symb_decoder(16#60#)) OR
 					(reg_q816 AND symb_decoder(16#ef#)) OR
 					(reg_q816 AND symb_decoder(16#1d#)) OR
 					(reg_q816 AND symb_decoder(16#7d#)) OR
 					(reg_q816 AND symb_decoder(16#8b#)) OR
 					(reg_q816 AND symb_decoder(16#e3#)) OR
 					(reg_q816 AND symb_decoder(16#d8#)) OR
 					(reg_q816 AND symb_decoder(16#6c#)) OR
 					(reg_q816 AND symb_decoder(16#c2#)) OR
 					(reg_q816 AND symb_decoder(16#7a#)) OR
 					(reg_q816 AND symb_decoder(16#9e#)) OR
 					(reg_q816 AND symb_decoder(16#7e#)) OR
 					(reg_q816 AND symb_decoder(16#32#)) OR
 					(reg_q816 AND symb_decoder(16#03#)) OR
 					(reg_q816 AND symb_decoder(16#57#)) OR
 					(reg_q816 AND symb_decoder(16#59#)) OR
 					(reg_q816 AND symb_decoder(16#ce#)) OR
 					(reg_q816 AND symb_decoder(16#c0#)) OR
 					(reg_q816 AND symb_decoder(16#3e#)) OR
 					(reg_q816 AND symb_decoder(16#a9#)) OR
 					(reg_q816 AND symb_decoder(16#82#)) OR
 					(reg_q816 AND symb_decoder(16#6b#)) OR
 					(reg_q816 AND symb_decoder(16#af#)) OR
 					(reg_q816 AND symb_decoder(16#6a#)) OR
 					(reg_q816 AND symb_decoder(16#2f#)) OR
 					(reg_q816 AND symb_decoder(16#b7#)) OR
 					(reg_q816 AND symb_decoder(16#54#)) OR
 					(reg_q816 AND symb_decoder(16#cd#)) OR
 					(reg_q816 AND symb_decoder(16#e7#)) OR
 					(reg_q816 AND symb_decoder(16#dc#)) OR
 					(reg_q816 AND symb_decoder(16#ad#)) OR
 					(reg_q816 AND symb_decoder(16#6e#)) OR
 					(reg_q816 AND symb_decoder(16#a7#)) OR
 					(reg_q816 AND symb_decoder(16#db#)) OR
 					(reg_q816 AND symb_decoder(16#7b#)) OR
 					(reg_q816 AND symb_decoder(16#f2#)) OR
 					(reg_q816 AND symb_decoder(16#17#)) OR
 					(reg_q816 AND symb_decoder(16#cc#)) OR
 					(reg_q816 AND symb_decoder(16#61#)) OR
 					(reg_q816 AND symb_decoder(16#d0#)) OR
 					(reg_q816 AND symb_decoder(16#43#)) OR
 					(reg_q816 AND symb_decoder(16#76#)) OR
 					(reg_q816 AND symb_decoder(16#87#)) OR
 					(reg_q816 AND symb_decoder(16#f9#)) OR
 					(reg_q816 AND symb_decoder(16#66#)) OR
 					(reg_q816 AND symb_decoder(16#e0#)) OR
 					(reg_q816 AND symb_decoder(16#40#)) OR
 					(reg_q816 AND symb_decoder(16#9d#)) OR
 					(reg_q816 AND symb_decoder(16#3b#)) OR
 					(reg_q816 AND symb_decoder(16#80#)) OR
 					(reg_q816 AND symb_decoder(16#bd#)) OR
 					(reg_q816 AND symb_decoder(16#a5#)) OR
 					(reg_q816 AND symb_decoder(16#2a#)) OR
 					(reg_q816 AND symb_decoder(16#33#)) OR
 					(reg_q816 AND symb_decoder(16#a8#)) OR
 					(reg_q816 AND symb_decoder(16#41#)) OR
 					(reg_q816 AND symb_decoder(16#5a#)) OR
 					(reg_q816 AND symb_decoder(16#0f#)) OR
 					(reg_q816 AND symb_decoder(16#11#)) OR
 					(reg_q816 AND symb_decoder(16#47#)) OR
 					(reg_q816 AND symb_decoder(16#29#)) OR
 					(reg_q816 AND symb_decoder(16#50#)) OR
 					(reg_q816 AND symb_decoder(16#53#)) OR
 					(reg_q816 AND symb_decoder(16#de#)) OR
 					(reg_q816 AND symb_decoder(16#fb#)) OR
 					(reg_q816 AND symb_decoder(16#30#)) OR
 					(reg_q816 AND symb_decoder(16#4e#)) OR
 					(reg_q816 AND symb_decoder(16#ac#)) OR
 					(reg_q816 AND symb_decoder(16#98#)) OR
 					(reg_q816 AND symb_decoder(16#91#)) OR
 					(reg_q816 AND symb_decoder(16#63#)) OR
 					(reg_q816 AND symb_decoder(16#28#)) OR
 					(reg_q816 AND symb_decoder(16#09#)) OR
 					(reg_q816 AND symb_decoder(16#88#)) OR
 					(reg_q816 AND symb_decoder(16#00#)) OR
 					(reg_q816 AND symb_decoder(16#b2#)) OR
 					(reg_q816 AND symb_decoder(16#f4#)) OR
 					(reg_q816 AND symb_decoder(16#67#)) OR
 					(reg_q816 AND symb_decoder(16#ee#)) OR
 					(reg_q816 AND symb_decoder(16#b6#)) OR
 					(reg_q816 AND symb_decoder(16#9b#)) OR
 					(reg_q816 AND symb_decoder(16#ff#)) OR
 					(reg_q816 AND symb_decoder(16#ba#)) OR
 					(reg_q816 AND symb_decoder(16#ea#)) OR
 					(reg_q816 AND symb_decoder(16#0e#)) OR
 					(reg_q816 AND symb_decoder(16#18#)) OR
 					(reg_q816 AND symb_decoder(16#5f#)) OR
 					(reg_q816 AND symb_decoder(16#84#)) OR
 					(reg_q816 AND symb_decoder(16#35#)) OR
 					(reg_q816 AND symb_decoder(16#ca#)) OR
 					(reg_q816 AND symb_decoder(16#fe#)) OR
 					(reg_q816 AND symb_decoder(16#bf#)) OR
 					(reg_q816 AND symb_decoder(16#b0#)) OR
 					(reg_q816 AND symb_decoder(16#c5#)) OR
 					(reg_q816 AND symb_decoder(16#f8#)) OR
 					(reg_q816 AND symb_decoder(16#1b#)) OR
 					(reg_q816 AND symb_decoder(16#ab#)) OR
 					(reg_q816 AND symb_decoder(16#c1#)) OR
 					(reg_q816 AND symb_decoder(16#0a#)) OR
 					(reg_q816 AND symb_decoder(16#9a#)) OR
 					(reg_q816 AND symb_decoder(16#f5#)) OR
 					(reg_q816 AND symb_decoder(16#78#)) OR
 					(reg_q816 AND symb_decoder(16#31#)) OR
 					(reg_q816 AND symb_decoder(16#da#)) OR
 					(reg_q816 AND symb_decoder(16#73#)) OR
 					(reg_q816 AND symb_decoder(16#d1#)) OR
 					(reg_q816 AND symb_decoder(16#12#)) OR
 					(reg_q816 AND symb_decoder(16#3d#)) OR
 					(reg_q816 AND symb_decoder(16#38#)) OR
 					(reg_q816 AND symb_decoder(16#ec#)) OR
 					(reg_q816 AND symb_decoder(16#4b#)) OR
 					(reg_q816 AND symb_decoder(16#e2#)) OR
 					(reg_q816 AND symb_decoder(16#a1#)) OR
 					(reg_q816 AND symb_decoder(16#bb#)) OR
 					(reg_q816 AND symb_decoder(16#08#)) OR
 					(reg_q816 AND symb_decoder(16#48#)) OR
 					(reg_q816 AND symb_decoder(16#70#)) OR
 					(reg_q816 AND symb_decoder(16#ed#)) OR
 					(reg_q816 AND symb_decoder(16#b3#)) OR
 					(reg_q816 AND symb_decoder(16#3c#)) OR
 					(reg_q816 AND symb_decoder(16#94#)) OR
 					(reg_q816 AND symb_decoder(16#86#)) OR
 					(reg_q816 AND symb_decoder(16#cf#)) OR
 					(reg_q816 AND symb_decoder(16#fa#)) OR
 					(reg_q816 AND symb_decoder(16#0c#)) OR
 					(reg_q816 AND symb_decoder(16#46#)) OR
 					(reg_q816 AND symb_decoder(16#7c#)) OR
 					(reg_q816 AND symb_decoder(16#37#)) OR
 					(reg_q816 AND symb_decoder(16#20#)) OR
 					(reg_q816 AND symb_decoder(16#c6#)) OR
 					(reg_q816 AND symb_decoder(16#4f#)) OR
 					(reg_q816 AND symb_decoder(16#b4#)) OR
 					(reg_q816 AND symb_decoder(16#07#)) OR
 					(reg_q816 AND symb_decoder(16#52#)) OR
 					(reg_q816 AND symb_decoder(16#c3#)) OR
 					(reg_q816 AND symb_decoder(16#fd#)) OR
 					(reg_q816 AND symb_decoder(16#e9#)) OR
 					(reg_q816 AND symb_decoder(16#45#)) OR
 					(reg_q816 AND symb_decoder(16#22#)) OR
 					(reg_q816 AND symb_decoder(16#27#)) OR
 					(reg_q816 AND symb_decoder(16#e5#)) OR
 					(reg_q816 AND symb_decoder(16#c4#)) OR
 					(reg_q816 AND symb_decoder(16#10#)) OR
 					(reg_q816 AND symb_decoder(16#8d#)) OR
 					(reg_q816 AND symb_decoder(16#0d#)) OR
 					(reg_q816 AND symb_decoder(16#eb#)) OR
 					(reg_q816 AND symb_decoder(16#c9#)) OR
 					(reg_q816 AND symb_decoder(16#3f#)) OR
 					(reg_q816 AND symb_decoder(16#34#)) OR
 					(reg_q816 AND symb_decoder(16#d6#)) OR
 					(reg_q816 AND symb_decoder(16#6f#)) OR
 					(reg_q816 AND symb_decoder(16#55#)) OR
 					(reg_q816 AND symb_decoder(16#d9#)) OR
 					(reg_q816 AND symb_decoder(16#92#)) OR
 					(reg_q816 AND symb_decoder(16#8a#)) OR
 					(reg_q816 AND symb_decoder(16#d2#)) OR
 					(reg_q816 AND symb_decoder(16#15#)) OR
 					(reg_q816 AND symb_decoder(16#be#)) OR
 					(reg_q816 AND symb_decoder(16#79#)) OR
 					(reg_q816 AND symb_decoder(16#4d#)) OR
 					(reg_q816 AND symb_decoder(16#99#)) OR
 					(reg_q816 AND symb_decoder(16#a4#)) OR
 					(reg_q816 AND symb_decoder(16#06#)) OR
 					(reg_q816 AND symb_decoder(16#e6#)) OR
 					(reg_q816 AND symb_decoder(16#4a#)) OR
 					(reg_q816 AND symb_decoder(16#d7#)) OR
 					(reg_q816 AND symb_decoder(16#97#)) OR
 					(reg_q816 AND symb_decoder(16#95#)) OR
 					(reg_q816 AND symb_decoder(16#f6#)) OR
 					(reg_q816 AND symb_decoder(16#13#)) OR
 					(reg_q816 AND symb_decoder(16#a0#)) OR
 					(reg_q816 AND symb_decoder(16#36#)) OR
 					(reg_q816 AND symb_decoder(16#1e#)) OR
 					(reg_q816 AND symb_decoder(16#ae#)) OR
 					(reg_q816 AND symb_decoder(16#df#)) OR
 					(reg_q816 AND symb_decoder(16#e8#)) OR
 					(reg_q816 AND symb_decoder(16#89#)) OR
 					(reg_q816 AND symb_decoder(16#a3#)) OR
 					(reg_q816 AND symb_decoder(16#25#)) OR
 					(reg_q816 AND symb_decoder(16#74#)) OR
 					(reg_q816 AND symb_decoder(16#49#)) OR
 					(reg_q816 AND symb_decoder(16#1f#)) OR
 					(reg_q816 AND symb_decoder(16#56#)) OR
 					(reg_q816 AND symb_decoder(16#69#)) OR
 					(reg_q816 AND symb_decoder(16#e4#)) OR
 					(reg_q816 AND symb_decoder(16#51#)) OR
 					(reg_q816 AND symb_decoder(16#b9#)) OR
 					(reg_q816 AND symb_decoder(16#e1#)) OR
 					(reg_q816 AND symb_decoder(16#58#)) OR
 					(reg_q816 AND symb_decoder(16#62#)) OR
 					(reg_q816 AND symb_decoder(16#f3#)) OR
 					(reg_q816 AND symb_decoder(16#f1#)) OR
 					(reg_q816 AND symb_decoder(16#8c#)) OR
 					(reg_q816 AND symb_decoder(16#2c#)) OR
 					(reg_q816 AND symb_decoder(16#b1#)) OR
 					(reg_q816 AND symb_decoder(16#24#)) OR
 					(reg_q816 AND symb_decoder(16#85#)) OR
 					(reg_q816 AND symb_decoder(16#7f#)) OR
 					(reg_q816 AND symb_decoder(16#1a#)) OR
 					(reg_q816 AND symb_decoder(16#d5#)) OR
 					(reg_q816 AND symb_decoder(16#83#)) OR
 					(reg_q816 AND symb_decoder(16#71#)) OR
 					(reg_q816 AND symb_decoder(16#96#)) OR
 					(reg_q816 AND symb_decoder(16#a2#)) OR
 					(reg_q816 AND symb_decoder(16#44#)) OR
 					(reg_q816 AND symb_decoder(16#5b#)) OR
 					(reg_q816 AND symb_decoder(16#5c#)) OR
 					(reg_q816 AND symb_decoder(16#23#)) OR
 					(reg_q816 AND symb_decoder(16#02#)) OR
 					(reg_q816 AND symb_decoder(16#2e#)) OR
 					(reg_q816 AND symb_decoder(16#01#)) OR
 					(reg_q816 AND symb_decoder(16#1c#)) OR
 					(reg_q816 AND symb_decoder(16#2b#)) OR
 					(reg_q816 AND symb_decoder(16#9c#)) OR
 					(reg_q816 AND symb_decoder(16#19#)) OR
 					(reg_q816 AND symb_decoder(16#64#)) OR
 					(reg_q816 AND symb_decoder(16#a6#)) OR
 					(reg_q816 AND symb_decoder(16#fc#)) OR
 					(reg_q816 AND symb_decoder(16#72#)) OR
 					(reg_q816 AND symb_decoder(16#c8#)) OR
 					(reg_q816 AND symb_decoder(16#5e#)) OR
 					(reg_q816 AND symb_decoder(16#b5#)) OR
 					(reg_q816 AND symb_decoder(16#81#)) OR
 					(reg_q816 AND symb_decoder(16#b8#)) OR
 					(reg_q816 AND symb_decoder(16#f7#)) OR
 					(reg_q816 AND symb_decoder(16#d3#)) OR
 					(reg_q816 AND symb_decoder(16#f0#)) OR
 					(reg_q816 AND symb_decoder(16#26#)) OR
 					(reg_q816 AND symb_decoder(16#90#)) OR
 					(reg_q816 AND symb_decoder(16#c7#)) OR
 					(reg_q816 AND symb_decoder(16#21#)) OR
 					(reg_q816 AND symb_decoder(16#bc#)) OR
 					(reg_q816 AND symb_decoder(16#5d#)) OR
 					(reg_q816 AND symb_decoder(16#65#));
reg_q816_init <= '0' ;
	p_reg_q816: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q816 <= reg_q816_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q816 <= reg_q816_init;
        else
          reg_q816 <= reg_q816_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1224_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1224 AND symb_decoder(16#4f#)) OR
 					(reg_q1224 AND symb_decoder(16#19#)) OR
 					(reg_q1224 AND symb_decoder(16#ba#)) OR
 					(reg_q1224 AND symb_decoder(16#51#)) OR
 					(reg_q1224 AND symb_decoder(16#bc#)) OR
 					(reg_q1224 AND symb_decoder(16#9d#)) OR
 					(reg_q1224 AND symb_decoder(16#88#)) OR
 					(reg_q1224 AND symb_decoder(16#d3#)) OR
 					(reg_q1224 AND symb_decoder(16#a8#)) OR
 					(reg_q1224 AND symb_decoder(16#6a#)) OR
 					(reg_q1224 AND symb_decoder(16#46#)) OR
 					(reg_q1224 AND symb_decoder(16#42#)) OR
 					(reg_q1224 AND symb_decoder(16#3d#)) OR
 					(reg_q1224 AND symb_decoder(16#9a#)) OR
 					(reg_q1224 AND symb_decoder(16#b2#)) OR
 					(reg_q1224 AND symb_decoder(16#00#)) OR
 					(reg_q1224 AND symb_decoder(16#33#)) OR
 					(reg_q1224 AND symb_decoder(16#3e#)) OR
 					(reg_q1224 AND symb_decoder(16#aa#)) OR
 					(reg_q1224 AND symb_decoder(16#58#)) OR
 					(reg_q1224 AND symb_decoder(16#bd#)) OR
 					(reg_q1224 AND symb_decoder(16#3b#)) OR
 					(reg_q1224 AND symb_decoder(16#b9#)) OR
 					(reg_q1224 AND symb_decoder(16#5d#)) OR
 					(reg_q1224 AND symb_decoder(16#af#)) OR
 					(reg_q1224 AND symb_decoder(16#84#)) OR
 					(reg_q1224 AND symb_decoder(16#d1#)) OR
 					(reg_q1224 AND symb_decoder(16#dc#)) OR
 					(reg_q1224 AND symb_decoder(16#e3#)) OR
 					(reg_q1224 AND symb_decoder(16#2d#)) OR
 					(reg_q1224 AND symb_decoder(16#d5#)) OR
 					(reg_q1224 AND symb_decoder(16#fa#)) OR
 					(reg_q1224 AND symb_decoder(16#90#)) OR
 					(reg_q1224 AND symb_decoder(16#7f#)) OR
 					(reg_q1224 AND symb_decoder(16#9e#)) OR
 					(reg_q1224 AND symb_decoder(16#0c#)) OR
 					(reg_q1224 AND symb_decoder(16#d7#)) OR
 					(reg_q1224 AND symb_decoder(16#f0#)) OR
 					(reg_q1224 AND symb_decoder(16#20#)) OR
 					(reg_q1224 AND symb_decoder(16#ff#)) OR
 					(reg_q1224 AND symb_decoder(16#4b#)) OR
 					(reg_q1224 AND symb_decoder(16#4e#)) OR
 					(reg_q1224 AND symb_decoder(16#1c#)) OR
 					(reg_q1224 AND symb_decoder(16#87#)) OR
 					(reg_q1224 AND symb_decoder(16#c4#)) OR
 					(reg_q1224 AND symb_decoder(16#ec#)) OR
 					(reg_q1224 AND symb_decoder(16#c8#)) OR
 					(reg_q1224 AND symb_decoder(16#c9#)) OR
 					(reg_q1224 AND symb_decoder(16#03#)) OR
 					(reg_q1224 AND symb_decoder(16#8c#)) OR
 					(reg_q1224 AND symb_decoder(16#21#)) OR
 					(reg_q1224 AND symb_decoder(16#3f#)) OR
 					(reg_q1224 AND symb_decoder(16#24#)) OR
 					(reg_q1224 AND symb_decoder(16#fb#)) OR
 					(reg_q1224 AND symb_decoder(16#f9#)) OR
 					(reg_q1224 AND symb_decoder(16#67#)) OR
 					(reg_q1224 AND symb_decoder(16#35#)) OR
 					(reg_q1224 AND symb_decoder(16#9c#)) OR
 					(reg_q1224 AND symb_decoder(16#e4#)) OR
 					(reg_q1224 AND symb_decoder(16#29#)) OR
 					(reg_q1224 AND symb_decoder(16#b3#)) OR
 					(reg_q1224 AND symb_decoder(16#50#)) OR
 					(reg_q1224 AND symb_decoder(16#02#)) OR
 					(reg_q1224 AND symb_decoder(16#8b#)) OR
 					(reg_q1224 AND symb_decoder(16#48#)) OR
 					(reg_q1224 AND symb_decoder(16#0b#)) OR
 					(reg_q1224 AND symb_decoder(16#57#)) OR
 					(reg_q1224 AND symb_decoder(16#66#)) OR
 					(reg_q1224 AND symb_decoder(16#60#)) OR
 					(reg_q1224 AND symb_decoder(16#6d#)) OR
 					(reg_q1224 AND symb_decoder(16#b1#)) OR
 					(reg_q1224 AND symb_decoder(16#c7#)) OR
 					(reg_q1224 AND symb_decoder(16#64#)) OR
 					(reg_q1224 AND symb_decoder(16#b4#)) OR
 					(reg_q1224 AND symb_decoder(16#f7#)) OR
 					(reg_q1224 AND symb_decoder(16#06#)) OR
 					(reg_q1224 AND symb_decoder(16#45#)) OR
 					(reg_q1224 AND symb_decoder(16#91#)) OR
 					(reg_q1224 AND symb_decoder(16#77#)) OR
 					(reg_q1224 AND symb_decoder(16#56#)) OR
 					(reg_q1224 AND symb_decoder(16#6b#)) OR
 					(reg_q1224 AND symb_decoder(16#47#)) OR
 					(reg_q1224 AND symb_decoder(16#ab#)) OR
 					(reg_q1224 AND symb_decoder(16#08#)) OR
 					(reg_q1224 AND symb_decoder(16#94#)) OR
 					(reg_q1224 AND symb_decoder(16#17#)) OR
 					(reg_q1224 AND symb_decoder(16#cf#)) OR
 					(reg_q1224 AND symb_decoder(16#bb#)) OR
 					(reg_q1224 AND symb_decoder(16#44#)) OR
 					(reg_q1224 AND symb_decoder(16#1d#)) OR
 					(reg_q1224 AND symb_decoder(16#41#)) OR
 					(reg_q1224 AND symb_decoder(16#e5#)) OR
 					(reg_q1224 AND symb_decoder(16#65#)) OR
 					(reg_q1224 AND symb_decoder(16#82#)) OR
 					(reg_q1224 AND symb_decoder(16#d9#)) OR
 					(reg_q1224 AND symb_decoder(16#92#)) OR
 					(reg_q1224 AND symb_decoder(16#d8#)) OR
 					(reg_q1224 AND symb_decoder(16#f4#)) OR
 					(reg_q1224 AND symb_decoder(16#ed#)) OR
 					(reg_q1224 AND symb_decoder(16#a5#)) OR
 					(reg_q1224 AND symb_decoder(16#c6#)) OR
 					(reg_q1224 AND symb_decoder(16#c3#)) OR
 					(reg_q1224 AND symb_decoder(16#dd#)) OR
 					(reg_q1224 AND symb_decoder(16#83#)) OR
 					(reg_q1224 AND symb_decoder(16#8f#)) OR
 					(reg_q1224 AND symb_decoder(16#4a#)) OR
 					(reg_q1224 AND symb_decoder(16#96#)) OR
 					(reg_q1224 AND symb_decoder(16#14#)) OR
 					(reg_q1224 AND symb_decoder(16#a2#)) OR
 					(reg_q1224 AND symb_decoder(16#a9#)) OR
 					(reg_q1224 AND symb_decoder(16#2c#)) OR
 					(reg_q1224 AND symb_decoder(16#c2#)) OR
 					(reg_q1224 AND symb_decoder(16#fe#)) OR
 					(reg_q1224 AND symb_decoder(16#f3#)) OR
 					(reg_q1224 AND symb_decoder(16#07#)) OR
 					(reg_q1224 AND symb_decoder(16#ca#)) OR
 					(reg_q1224 AND symb_decoder(16#a3#)) OR
 					(reg_q1224 AND symb_decoder(16#38#)) OR
 					(reg_q1224 AND symb_decoder(16#c5#)) OR
 					(reg_q1224 AND symb_decoder(16#5c#)) OR
 					(reg_q1224 AND symb_decoder(16#39#)) OR
 					(reg_q1224 AND symb_decoder(16#8e#)) OR
 					(reg_q1224 AND symb_decoder(16#7c#)) OR
 					(reg_q1224 AND symb_decoder(16#c0#)) OR
 					(reg_q1224 AND symb_decoder(16#1f#)) OR
 					(reg_q1224 AND symb_decoder(16#0a#)) OR
 					(reg_q1224 AND symb_decoder(16#53#)) OR
 					(reg_q1224 AND symb_decoder(16#93#)) OR
 					(reg_q1224 AND symb_decoder(16#cb#)) OR
 					(reg_q1224 AND symb_decoder(16#01#)) OR
 					(reg_q1224 AND symb_decoder(16#85#)) OR
 					(reg_q1224 AND symb_decoder(16#2a#)) OR
 					(reg_q1224 AND symb_decoder(16#70#)) OR
 					(reg_q1224 AND symb_decoder(16#d2#)) OR
 					(reg_q1224 AND symb_decoder(16#db#)) OR
 					(reg_q1224 AND symb_decoder(16#37#)) OR
 					(reg_q1224 AND symb_decoder(16#ee#)) OR
 					(reg_q1224 AND symb_decoder(16#26#)) OR
 					(reg_q1224 AND symb_decoder(16#5b#)) OR
 					(reg_q1224 AND symb_decoder(16#0e#)) OR
 					(reg_q1224 AND symb_decoder(16#7e#)) OR
 					(reg_q1224 AND symb_decoder(16#28#)) OR
 					(reg_q1224 AND symb_decoder(16#ef#)) OR
 					(reg_q1224 AND symb_decoder(16#e1#)) OR
 					(reg_q1224 AND symb_decoder(16#e9#)) OR
 					(reg_q1224 AND symb_decoder(16#0d#)) OR
 					(reg_q1224 AND symb_decoder(16#d6#)) OR
 					(reg_q1224 AND symb_decoder(16#be#)) OR
 					(reg_q1224 AND symb_decoder(16#16#)) OR
 					(reg_q1224 AND symb_decoder(16#05#)) OR
 					(reg_q1224 AND symb_decoder(16#10#)) OR
 					(reg_q1224 AND symb_decoder(16#3c#)) OR
 					(reg_q1224 AND symb_decoder(16#98#)) OR
 					(reg_q1224 AND symb_decoder(16#5f#)) OR
 					(reg_q1224 AND symb_decoder(16#5a#)) OR
 					(reg_q1224 AND symb_decoder(16#34#)) OR
 					(reg_q1224 AND symb_decoder(16#2e#)) OR
 					(reg_q1224 AND symb_decoder(16#7d#)) OR
 					(reg_q1224 AND symb_decoder(16#99#)) OR
 					(reg_q1224 AND symb_decoder(16#e7#)) OR
 					(reg_q1224 AND symb_decoder(16#95#)) OR
 					(reg_q1224 AND symb_decoder(16#25#)) OR
 					(reg_q1224 AND symb_decoder(16#d0#)) OR
 					(reg_q1224 AND symb_decoder(16#6e#)) OR
 					(reg_q1224 AND symb_decoder(16#ae#)) OR
 					(reg_q1224 AND symb_decoder(16#73#)) OR
 					(reg_q1224 AND symb_decoder(16#23#)) OR
 					(reg_q1224 AND symb_decoder(16#89#)) OR
 					(reg_q1224 AND symb_decoder(16#fc#)) OR
 					(reg_q1224 AND symb_decoder(16#61#)) OR
 					(reg_q1224 AND symb_decoder(16#6c#)) OR
 					(reg_q1224 AND symb_decoder(16#a0#)) OR
 					(reg_q1224 AND symb_decoder(16#52#)) OR
 					(reg_q1224 AND symb_decoder(16#e8#)) OR
 					(reg_q1224 AND symb_decoder(16#71#)) OR
 					(reg_q1224 AND symb_decoder(16#15#)) OR
 					(reg_q1224 AND symb_decoder(16#4c#)) OR
 					(reg_q1224 AND symb_decoder(16#43#)) OR
 					(reg_q1224 AND symb_decoder(16#f6#)) OR
 					(reg_q1224 AND symb_decoder(16#bf#)) OR
 					(reg_q1224 AND symb_decoder(16#c1#)) OR
 					(reg_q1224 AND symb_decoder(16#eb#)) OR
 					(reg_q1224 AND symb_decoder(16#ce#)) OR
 					(reg_q1224 AND symb_decoder(16#49#)) OR
 					(reg_q1224 AND symb_decoder(16#8d#)) OR
 					(reg_q1224 AND symb_decoder(16#f2#)) OR
 					(reg_q1224 AND symb_decoder(16#11#)) OR
 					(reg_q1224 AND symb_decoder(16#a7#)) OR
 					(reg_q1224 AND symb_decoder(16#4d#)) OR
 					(reg_q1224 AND symb_decoder(16#3a#)) OR
 					(reg_q1224 AND symb_decoder(16#63#)) OR
 					(reg_q1224 AND symb_decoder(16#da#)) OR
 					(reg_q1224 AND symb_decoder(16#80#)) OR
 					(reg_q1224 AND symb_decoder(16#97#)) OR
 					(reg_q1224 AND symb_decoder(16#76#)) OR
 					(reg_q1224 AND symb_decoder(16#a1#)) OR
 					(reg_q1224 AND symb_decoder(16#0f#)) OR
 					(reg_q1224 AND symb_decoder(16#1e#)) OR
 					(reg_q1224 AND symb_decoder(16#7a#)) OR
 					(reg_q1224 AND symb_decoder(16#1a#)) OR
 					(reg_q1224 AND symb_decoder(16#2f#)) OR
 					(reg_q1224 AND symb_decoder(16#04#)) OR
 					(reg_q1224 AND symb_decoder(16#df#)) OR
 					(reg_q1224 AND symb_decoder(16#8a#)) OR
 					(reg_q1224 AND symb_decoder(16#f1#)) OR
 					(reg_q1224 AND symb_decoder(16#ad#)) OR
 					(reg_q1224 AND symb_decoder(16#b6#)) OR
 					(reg_q1224 AND symb_decoder(16#32#)) OR
 					(reg_q1224 AND symb_decoder(16#7b#)) OR
 					(reg_q1224 AND symb_decoder(16#68#)) OR
 					(reg_q1224 AND symb_decoder(16#36#)) OR
 					(reg_q1224 AND symb_decoder(16#62#)) OR
 					(reg_q1224 AND symb_decoder(16#a4#)) OR
 					(reg_q1224 AND symb_decoder(16#2b#)) OR
 					(reg_q1224 AND symb_decoder(16#9f#)) OR
 					(reg_q1224 AND symb_decoder(16#e2#)) OR
 					(reg_q1224 AND symb_decoder(16#b5#)) OR
 					(reg_q1224 AND symb_decoder(16#ea#)) OR
 					(reg_q1224 AND symb_decoder(16#54#)) OR
 					(reg_q1224 AND symb_decoder(16#cd#)) OR
 					(reg_q1224 AND symb_decoder(16#78#)) OR
 					(reg_q1224 AND symb_decoder(16#a6#)) OR
 					(reg_q1224 AND symb_decoder(16#74#)) OR
 					(reg_q1224 AND symb_decoder(16#1b#)) OR
 					(reg_q1224 AND symb_decoder(16#13#)) OR
 					(reg_q1224 AND symb_decoder(16#79#)) OR
 					(reg_q1224 AND symb_decoder(16#40#)) OR
 					(reg_q1224 AND symb_decoder(16#12#)) OR
 					(reg_q1224 AND symb_decoder(16#75#)) OR
 					(reg_q1224 AND symb_decoder(16#cc#)) OR
 					(reg_q1224 AND symb_decoder(16#30#)) OR
 					(reg_q1224 AND symb_decoder(16#ac#)) OR
 					(reg_q1224 AND symb_decoder(16#09#)) OR
 					(reg_q1224 AND symb_decoder(16#b0#)) OR
 					(reg_q1224 AND symb_decoder(16#f5#)) OR
 					(reg_q1224 AND symb_decoder(16#9b#)) OR
 					(reg_q1224 AND symb_decoder(16#69#)) OR
 					(reg_q1224 AND symb_decoder(16#fd#)) OR
 					(reg_q1224 AND symb_decoder(16#59#)) OR
 					(reg_q1224 AND symb_decoder(16#e0#)) OR
 					(reg_q1224 AND symb_decoder(16#18#)) OR
 					(reg_q1224 AND symb_decoder(16#81#)) OR
 					(reg_q1224 AND symb_decoder(16#b8#)) OR
 					(reg_q1224 AND symb_decoder(16#72#)) OR
 					(reg_q1224 AND symb_decoder(16#d4#)) OR
 					(reg_q1224 AND symb_decoder(16#e6#)) OR
 					(reg_q1224 AND symb_decoder(16#55#)) OR
 					(reg_q1224 AND symb_decoder(16#86#)) OR
 					(reg_q1224 AND symb_decoder(16#f8#)) OR
 					(reg_q1224 AND symb_decoder(16#b7#)) OR
 					(reg_q1224 AND symb_decoder(16#5e#)) OR
 					(reg_q1224 AND symb_decoder(16#22#)) OR
 					(reg_q1224 AND symb_decoder(16#de#)) OR
 					(reg_q1224 AND symb_decoder(16#31#)) OR
 					(reg_q1224 AND symb_decoder(16#6f#)) OR
 					(reg_q1224 AND symb_decoder(16#27#));
reg_q1224_init <= '0' ;
	p_reg_q1224: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1224 <= reg_q1224_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1224 <= reg_q1224_init;
        else
          reg_q1224 <= reg_q1224_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q896_in <= (reg_q889 AND symb_decoder(16#29#)) OR
 					(reg_q889 AND symb_decoder(16#94#)) OR
 					(reg_q889 AND symb_decoder(16#e2#)) OR
 					(reg_q889 AND symb_decoder(16#a0#)) OR
 					(reg_q889 AND symb_decoder(16#bc#)) OR
 					(reg_q889 AND symb_decoder(16#67#)) OR
 					(reg_q889 AND symb_decoder(16#6e#)) OR
 					(reg_q889 AND symb_decoder(16#a7#)) OR
 					(reg_q889 AND symb_decoder(16#e4#)) OR
 					(reg_q889 AND symb_decoder(16#14#)) OR
 					(reg_q889 AND symb_decoder(16#78#)) OR
 					(reg_q889 AND symb_decoder(16#27#)) OR
 					(reg_q889 AND symb_decoder(16#4e#)) OR
 					(reg_q889 AND symb_decoder(16#8b#)) OR
 					(reg_q889 AND symb_decoder(16#aa#)) OR
 					(reg_q889 AND symb_decoder(16#7e#)) OR
 					(reg_q889 AND symb_decoder(16#c2#)) OR
 					(reg_q889 AND symb_decoder(16#98#)) OR
 					(reg_q889 AND symb_decoder(16#31#)) OR
 					(reg_q889 AND symb_decoder(16#33#)) OR
 					(reg_q889 AND symb_decoder(16#5a#)) OR
 					(reg_q889 AND symb_decoder(16#f7#)) OR
 					(reg_q889 AND symb_decoder(16#72#)) OR
 					(reg_q889 AND symb_decoder(16#3b#)) OR
 					(reg_q889 AND symb_decoder(16#4c#)) OR
 					(reg_q889 AND symb_decoder(16#99#)) OR
 					(reg_q889 AND symb_decoder(16#ac#)) OR
 					(reg_q889 AND symb_decoder(16#ec#)) OR
 					(reg_q889 AND symb_decoder(16#b2#)) OR
 					(reg_q889 AND symb_decoder(16#d5#)) OR
 					(reg_q889 AND symb_decoder(16#bf#)) OR
 					(reg_q889 AND symb_decoder(16#fd#)) OR
 					(reg_q889 AND symb_decoder(16#07#)) OR
 					(reg_q889 AND symb_decoder(16#62#)) OR
 					(reg_q889 AND symb_decoder(16#09#)) OR
 					(reg_q889 AND symb_decoder(16#0e#)) OR
 					(reg_q889 AND symb_decoder(16#c1#)) OR
 					(reg_q889 AND symb_decoder(16#a4#)) OR
 					(reg_q889 AND symb_decoder(16#9a#)) OR
 					(reg_q889 AND symb_decoder(16#15#)) OR
 					(reg_q889 AND symb_decoder(16#06#)) OR
 					(reg_q889 AND symb_decoder(16#69#)) OR
 					(reg_q889 AND symb_decoder(16#ce#)) OR
 					(reg_q889 AND symb_decoder(16#76#)) OR
 					(reg_q889 AND symb_decoder(16#61#)) OR
 					(reg_q889 AND symb_decoder(16#e9#)) OR
 					(reg_q889 AND symb_decoder(16#d1#)) OR
 					(reg_q889 AND symb_decoder(16#9e#)) OR
 					(reg_q889 AND symb_decoder(16#85#)) OR
 					(reg_q889 AND symb_decoder(16#ef#)) OR
 					(reg_q889 AND symb_decoder(16#3f#)) OR
 					(reg_q889 AND symb_decoder(16#c5#)) OR
 					(reg_q889 AND symb_decoder(16#7c#)) OR
 					(reg_q889 AND symb_decoder(16#dd#)) OR
 					(reg_q889 AND symb_decoder(16#64#)) OR
 					(reg_q889 AND symb_decoder(16#36#)) OR
 					(reg_q889 AND symb_decoder(16#60#)) OR
 					(reg_q889 AND symb_decoder(16#96#)) OR
 					(reg_q889 AND symb_decoder(16#3a#)) OR
 					(reg_q889 AND symb_decoder(16#d3#)) OR
 					(reg_q889 AND symb_decoder(16#ba#)) OR
 					(reg_q889 AND symb_decoder(16#23#)) OR
 					(reg_q889 AND symb_decoder(16#e1#)) OR
 					(reg_q889 AND symb_decoder(16#32#)) OR
 					(reg_q889 AND symb_decoder(16#04#)) OR
 					(reg_q889 AND symb_decoder(16#03#)) OR
 					(reg_q889 AND symb_decoder(16#c0#)) OR
 					(reg_q889 AND symb_decoder(16#b8#)) OR
 					(reg_q889 AND symb_decoder(16#f5#)) OR
 					(reg_q889 AND symb_decoder(16#2f#)) OR
 					(reg_q889 AND symb_decoder(16#b7#)) OR
 					(reg_q889 AND symb_decoder(16#02#)) OR
 					(reg_q889 AND symb_decoder(16#c9#)) OR
 					(reg_q889 AND symb_decoder(16#f9#)) OR
 					(reg_q889 AND symb_decoder(16#b3#)) OR
 					(reg_q889 AND symb_decoder(16#d4#)) OR
 					(reg_q889 AND symb_decoder(16#d8#)) OR
 					(reg_q889 AND symb_decoder(16#5f#)) OR
 					(reg_q889 AND symb_decoder(16#6c#)) OR
 					(reg_q889 AND symb_decoder(16#95#)) OR
 					(reg_q889 AND symb_decoder(16#6a#)) OR
 					(reg_q889 AND symb_decoder(16#77#)) OR
 					(reg_q889 AND symb_decoder(16#65#)) OR
 					(reg_q889 AND symb_decoder(16#e8#)) OR
 					(reg_q889 AND symb_decoder(16#25#)) OR
 					(reg_q889 AND symb_decoder(16#7d#)) OR
 					(reg_q889 AND symb_decoder(16#9d#)) OR
 					(reg_q889 AND symb_decoder(16#ee#)) OR
 					(reg_q889 AND symb_decoder(16#5e#)) OR
 					(reg_q889 AND symb_decoder(16#1b#)) OR
 					(reg_q889 AND symb_decoder(16#19#)) OR
 					(reg_q889 AND symb_decoder(16#1c#)) OR
 					(reg_q889 AND symb_decoder(16#a1#)) OR
 					(reg_q889 AND symb_decoder(16#83#)) OR
 					(reg_q889 AND symb_decoder(16#45#)) OR
 					(reg_q889 AND symb_decoder(16#c7#)) OR
 					(reg_q889 AND symb_decoder(16#5b#)) OR
 					(reg_q889 AND symb_decoder(16#12#)) OR
 					(reg_q889 AND symb_decoder(16#42#)) OR
 					(reg_q889 AND symb_decoder(16#30#)) OR
 					(reg_q889 AND symb_decoder(16#a8#)) OR
 					(reg_q889 AND symb_decoder(16#fa#)) OR
 					(reg_q889 AND symb_decoder(16#a5#)) OR
 					(reg_q889 AND symb_decoder(16#18#)) OR
 					(reg_q889 AND symb_decoder(16#dc#)) OR
 					(reg_q889 AND symb_decoder(16#00#)) OR
 					(reg_q889 AND symb_decoder(16#6b#)) OR
 					(reg_q889 AND symb_decoder(16#56#)) OR
 					(reg_q889 AND symb_decoder(16#0d#)) OR
 					(reg_q889 AND symb_decoder(16#be#)) OR
 					(reg_q889 AND symb_decoder(16#35#)) OR
 					(reg_q889 AND symb_decoder(16#4a#)) OR
 					(reg_q889 AND symb_decoder(16#7b#)) OR
 					(reg_q889 AND symb_decoder(16#5c#)) OR
 					(reg_q889 AND symb_decoder(16#86#)) OR
 					(reg_q889 AND symb_decoder(16#3d#)) OR
 					(reg_q889 AND symb_decoder(16#2a#)) OR
 					(reg_q889 AND symb_decoder(16#40#)) OR
 					(reg_q889 AND symb_decoder(16#92#)) OR
 					(reg_q889 AND symb_decoder(16#ae#)) OR
 					(reg_q889 AND symb_decoder(16#05#)) OR
 					(reg_q889 AND symb_decoder(16#eb#)) OR
 					(reg_q889 AND symb_decoder(16#4d#)) OR
 					(reg_q889 AND symb_decoder(16#ed#)) OR
 					(reg_q889 AND symb_decoder(16#af#)) OR
 					(reg_q889 AND symb_decoder(16#2b#)) OR
 					(reg_q889 AND symb_decoder(16#9b#)) OR
 					(reg_q889 AND symb_decoder(16#0c#)) OR
 					(reg_q889 AND symb_decoder(16#ca#)) OR
 					(reg_q889 AND symb_decoder(16#39#)) OR
 					(reg_q889 AND symb_decoder(16#b1#)) OR
 					(reg_q889 AND symb_decoder(16#c4#)) OR
 					(reg_q889 AND symb_decoder(16#f1#)) OR
 					(reg_q889 AND symb_decoder(16#d7#)) OR
 					(reg_q889 AND symb_decoder(16#38#)) OR
 					(reg_q889 AND symb_decoder(16#87#)) OR
 					(reg_q889 AND symb_decoder(16#2d#)) OR
 					(reg_q889 AND symb_decoder(16#47#)) OR
 					(reg_q889 AND symb_decoder(16#c3#)) OR
 					(reg_q889 AND symb_decoder(16#13#)) OR
 					(reg_q889 AND symb_decoder(16#3c#)) OR
 					(reg_q889 AND symb_decoder(16#a2#)) OR
 					(reg_q889 AND symb_decoder(16#3e#)) OR
 					(reg_q889 AND symb_decoder(16#cd#)) OR
 					(reg_q889 AND symb_decoder(16#54#)) OR
 					(reg_q889 AND symb_decoder(16#1e#)) OR
 					(reg_q889 AND symb_decoder(16#55#)) OR
 					(reg_q889 AND symb_decoder(16#80#)) OR
 					(reg_q889 AND symb_decoder(16#db#)) OR
 					(reg_q889 AND symb_decoder(16#de#)) OR
 					(reg_q889 AND symb_decoder(16#71#)) OR
 					(reg_q889 AND symb_decoder(16#81#)) OR
 					(reg_q889 AND symb_decoder(16#51#)) OR
 					(reg_q889 AND symb_decoder(16#c8#)) OR
 					(reg_q889 AND symb_decoder(16#ea#)) OR
 					(reg_q889 AND symb_decoder(16#fe#)) OR
 					(reg_q889 AND symb_decoder(16#41#)) OR
 					(reg_q889 AND symb_decoder(16#cf#)) OR
 					(reg_q889 AND symb_decoder(16#1f#)) OR
 					(reg_q889 AND symb_decoder(16#fb#)) OR
 					(reg_q889 AND symb_decoder(16#e6#)) OR
 					(reg_q889 AND symb_decoder(16#17#)) OR
 					(reg_q889 AND symb_decoder(16#6f#)) OR
 					(reg_q889 AND symb_decoder(16#d0#)) OR
 					(reg_q889 AND symb_decoder(16#fc#)) OR
 					(reg_q889 AND symb_decoder(16#53#)) OR
 					(reg_q889 AND symb_decoder(16#5d#)) OR
 					(reg_q889 AND symb_decoder(16#01#)) OR
 					(reg_q889 AND symb_decoder(16#cc#)) OR
 					(reg_q889 AND symb_decoder(16#1d#)) OR
 					(reg_q889 AND symb_decoder(16#0a#)) OR
 					(reg_q889 AND symb_decoder(16#9f#)) OR
 					(reg_q889 AND symb_decoder(16#73#)) OR
 					(reg_q889 AND symb_decoder(16#a9#)) OR
 					(reg_q889 AND symb_decoder(16#a3#)) OR
 					(reg_q889 AND symb_decoder(16#b9#)) OR
 					(reg_q889 AND symb_decoder(16#c6#)) OR
 					(reg_q889 AND symb_decoder(16#b5#)) OR
 					(reg_q889 AND symb_decoder(16#a6#)) OR
 					(reg_q889 AND symb_decoder(16#93#)) OR
 					(reg_q889 AND symb_decoder(16#52#)) OR
 					(reg_q889 AND symb_decoder(16#34#)) OR
 					(reg_q889 AND symb_decoder(16#66#)) OR
 					(reg_q889 AND symb_decoder(16#90#)) OR
 					(reg_q889 AND symb_decoder(16#82#)) OR
 					(reg_q889 AND symb_decoder(16#10#)) OR
 					(reg_q889 AND symb_decoder(16#f8#)) OR
 					(reg_q889 AND symb_decoder(16#58#)) OR
 					(reg_q889 AND symb_decoder(16#22#)) OR
 					(reg_q889 AND symb_decoder(16#21#)) OR
 					(reg_q889 AND symb_decoder(16#2e#)) OR
 					(reg_q889 AND symb_decoder(16#20#)) OR
 					(reg_q889 AND symb_decoder(16#f6#)) OR
 					(reg_q889 AND symb_decoder(16#ad#)) OR
 					(reg_q889 AND symb_decoder(16#4f#)) OR
 					(reg_q889 AND symb_decoder(16#43#)) OR
 					(reg_q889 AND symb_decoder(16#26#)) OR
 					(reg_q889 AND symb_decoder(16#37#)) OR
 					(reg_q889 AND symb_decoder(16#b6#)) OR
 					(reg_q889 AND symb_decoder(16#24#)) OR
 					(reg_q889 AND symb_decoder(16#0b#)) OR
 					(reg_q889 AND symb_decoder(16#44#)) OR
 					(reg_q889 AND symb_decoder(16#b4#)) OR
 					(reg_q889 AND symb_decoder(16#16#)) OR
 					(reg_q889 AND symb_decoder(16#f2#)) OR
 					(reg_q889 AND symb_decoder(16#bb#)) OR
 					(reg_q889 AND symb_decoder(16#d9#)) OR
 					(reg_q889 AND symb_decoder(16#e7#)) OR
 					(reg_q889 AND symb_decoder(16#08#)) OR
 					(reg_q889 AND symb_decoder(16#2c#)) OR
 					(reg_q889 AND symb_decoder(16#8c#)) OR
 					(reg_q889 AND symb_decoder(16#59#)) OR
 					(reg_q889 AND symb_decoder(16#f3#)) OR
 					(reg_q889 AND symb_decoder(16#e5#)) OR
 					(reg_q889 AND symb_decoder(16#4b#)) OR
 					(reg_q889 AND symb_decoder(16#8e#)) OR
 					(reg_q889 AND symb_decoder(16#48#)) OR
 					(reg_q889 AND symb_decoder(16#68#)) OR
 					(reg_q889 AND symb_decoder(16#d2#)) OR
 					(reg_q889 AND symb_decoder(16#0f#)) OR
 					(reg_q889 AND symb_decoder(16#57#)) OR
 					(reg_q889 AND symb_decoder(16#8d#)) OR
 					(reg_q889 AND symb_decoder(16#50#)) OR
 					(reg_q889 AND symb_decoder(16#97#)) OR
 					(reg_q889 AND symb_decoder(16#f4#)) OR
 					(reg_q889 AND symb_decoder(16#cb#)) OR
 					(reg_q889 AND symb_decoder(16#79#)) OR
 					(reg_q889 AND symb_decoder(16#ab#)) OR
 					(reg_q889 AND symb_decoder(16#89#)) OR
 					(reg_q889 AND symb_decoder(16#11#)) OR
 					(reg_q889 AND symb_decoder(16#ff#)) OR
 					(reg_q889 AND symb_decoder(16#49#)) OR
 					(reg_q889 AND symb_decoder(16#6d#)) OR
 					(reg_q889 AND symb_decoder(16#bd#)) OR
 					(reg_q889 AND symb_decoder(16#e0#)) OR
 					(reg_q889 AND symb_decoder(16#e3#)) OR
 					(reg_q889 AND symb_decoder(16#88#)) OR
 					(reg_q889 AND symb_decoder(16#70#)) OR
 					(reg_q889 AND symb_decoder(16#75#)) OR
 					(reg_q889 AND symb_decoder(16#91#)) OR
 					(reg_q889 AND symb_decoder(16#46#)) OR
 					(reg_q889 AND symb_decoder(16#1a#)) OR
 					(reg_q889 AND symb_decoder(16#9c#)) OR
 					(reg_q889 AND symb_decoder(16#7f#)) OR
 					(reg_q889 AND symb_decoder(16#b0#)) OR
 					(reg_q889 AND symb_decoder(16#84#)) OR
 					(reg_q889 AND symb_decoder(16#8f#)) OR
 					(reg_q889 AND symb_decoder(16#f0#)) OR
 					(reg_q889 AND symb_decoder(16#df#)) OR
 					(reg_q889 AND symb_decoder(16#74#)) OR
 					(reg_q889 AND symb_decoder(16#da#)) OR
 					(reg_q889 AND symb_decoder(16#63#)) OR
 					(reg_q889 AND symb_decoder(16#7a#)) OR
 					(reg_q889 AND symb_decoder(16#8a#)) OR
 					(reg_q889 AND symb_decoder(16#d6#)) OR
 					(reg_q889 AND symb_decoder(16#28#)) OR
 					(reg_q896 AND symb_decoder(16#5d#)) OR
 					(reg_q896 AND symb_decoder(16#c0#)) OR
 					(reg_q896 AND symb_decoder(16#74#)) OR
 					(reg_q896 AND symb_decoder(16#ed#)) OR
 					(reg_q896 AND symb_decoder(16#46#)) OR
 					(reg_q896 AND symb_decoder(16#ac#)) OR
 					(reg_q896 AND symb_decoder(16#bd#)) OR
 					(reg_q896 AND symb_decoder(16#5f#)) OR
 					(reg_q896 AND symb_decoder(16#f0#)) OR
 					(reg_q896 AND symb_decoder(16#ee#)) OR
 					(reg_q896 AND symb_decoder(16#66#)) OR
 					(reg_q896 AND symb_decoder(16#b0#)) OR
 					(reg_q896 AND symb_decoder(16#38#)) OR
 					(reg_q896 AND symb_decoder(16#6e#)) OR
 					(reg_q896 AND symb_decoder(16#52#)) OR
 					(reg_q896 AND symb_decoder(16#5c#)) OR
 					(reg_q896 AND symb_decoder(16#14#)) OR
 					(reg_q896 AND symb_decoder(16#3c#)) OR
 					(reg_q896 AND symb_decoder(16#91#)) OR
 					(reg_q896 AND symb_decoder(16#c3#)) OR
 					(reg_q896 AND symb_decoder(16#f2#)) OR
 					(reg_q896 AND symb_decoder(16#df#)) OR
 					(reg_q896 AND symb_decoder(16#87#)) OR
 					(reg_q896 AND symb_decoder(16#1b#)) OR
 					(reg_q896 AND symb_decoder(16#29#)) OR
 					(reg_q896 AND symb_decoder(16#b4#)) OR
 					(reg_q896 AND symb_decoder(16#4b#)) OR
 					(reg_q896 AND symb_decoder(16#82#)) OR
 					(reg_q896 AND symb_decoder(16#4f#)) OR
 					(reg_q896 AND symb_decoder(16#e9#)) OR
 					(reg_q896 AND symb_decoder(16#fe#)) OR
 					(reg_q896 AND symb_decoder(16#c9#)) OR
 					(reg_q896 AND symb_decoder(16#37#)) OR
 					(reg_q896 AND symb_decoder(16#28#)) OR
 					(reg_q896 AND symb_decoder(16#9c#)) OR
 					(reg_q896 AND symb_decoder(16#80#)) OR
 					(reg_q896 AND symb_decoder(16#12#)) OR
 					(reg_q896 AND symb_decoder(16#33#)) OR
 					(reg_q896 AND symb_decoder(16#15#)) OR
 					(reg_q896 AND symb_decoder(16#79#)) OR
 					(reg_q896 AND symb_decoder(16#4d#)) OR
 					(reg_q896 AND symb_decoder(16#78#)) OR
 					(reg_q896 AND symb_decoder(16#f9#)) OR
 					(reg_q896 AND symb_decoder(16#03#)) OR
 					(reg_q896 AND symb_decoder(16#4e#)) OR
 					(reg_q896 AND symb_decoder(16#bc#)) OR
 					(reg_q896 AND symb_decoder(16#71#)) OR
 					(reg_q896 AND symb_decoder(16#60#)) OR
 					(reg_q896 AND symb_decoder(16#a0#)) OR
 					(reg_q896 AND symb_decoder(16#55#)) OR
 					(reg_q896 AND symb_decoder(16#02#)) OR
 					(reg_q896 AND symb_decoder(16#36#)) OR
 					(reg_q896 AND symb_decoder(16#f5#)) OR
 					(reg_q896 AND symb_decoder(16#e5#)) OR
 					(reg_q896 AND symb_decoder(16#cc#)) OR
 					(reg_q896 AND symb_decoder(16#4c#)) OR
 					(reg_q896 AND symb_decoder(16#18#)) OR
 					(reg_q896 AND symb_decoder(16#2a#)) OR
 					(reg_q896 AND symb_decoder(16#08#)) OR
 					(reg_q896 AND symb_decoder(16#e2#)) OR
 					(reg_q896 AND symb_decoder(16#d0#)) OR
 					(reg_q896 AND symb_decoder(16#58#)) OR
 					(reg_q896 AND symb_decoder(16#e7#)) OR
 					(reg_q896 AND symb_decoder(16#3e#)) OR
 					(reg_q896 AND symb_decoder(16#00#)) OR
 					(reg_q896 AND symb_decoder(16#2d#)) OR
 					(reg_q896 AND symb_decoder(16#2f#)) OR
 					(reg_q896 AND symb_decoder(16#9f#)) OR
 					(reg_q896 AND symb_decoder(16#da#)) OR
 					(reg_q896 AND symb_decoder(16#c6#)) OR
 					(reg_q896 AND symb_decoder(16#a3#)) OR
 					(reg_q896 AND symb_decoder(16#c4#)) OR
 					(reg_q896 AND symb_decoder(16#0d#)) OR
 					(reg_q896 AND symb_decoder(16#fc#)) OR
 					(reg_q896 AND symb_decoder(16#ba#)) OR
 					(reg_q896 AND symb_decoder(16#76#)) OR
 					(reg_q896 AND symb_decoder(16#05#)) OR
 					(reg_q896 AND symb_decoder(16#ec#)) OR
 					(reg_q896 AND symb_decoder(16#39#)) OR
 					(reg_q896 AND symb_decoder(16#24#)) OR
 					(reg_q896 AND symb_decoder(16#7e#)) OR
 					(reg_q896 AND symb_decoder(16#d2#)) OR
 					(reg_q896 AND symb_decoder(16#45#)) OR
 					(reg_q896 AND symb_decoder(16#92#)) OR
 					(reg_q896 AND symb_decoder(16#1e#)) OR
 					(reg_q896 AND symb_decoder(16#34#)) OR
 					(reg_q896 AND symb_decoder(16#90#)) OR
 					(reg_q896 AND symb_decoder(16#cb#)) OR
 					(reg_q896 AND symb_decoder(16#0a#)) OR
 					(reg_q896 AND symb_decoder(16#35#)) OR
 					(reg_q896 AND symb_decoder(16#d7#)) OR
 					(reg_q896 AND symb_decoder(16#ff#)) OR
 					(reg_q896 AND symb_decoder(16#d1#)) OR
 					(reg_q896 AND symb_decoder(16#ab#)) OR
 					(reg_q896 AND symb_decoder(16#cd#)) OR
 					(reg_q896 AND symb_decoder(16#54#)) OR
 					(reg_q896 AND symb_decoder(16#f3#)) OR
 					(reg_q896 AND symb_decoder(16#8b#)) OR
 					(reg_q896 AND symb_decoder(16#72#)) OR
 					(reg_q896 AND symb_decoder(16#dd#)) OR
 					(reg_q896 AND symb_decoder(16#8a#)) OR
 					(reg_q896 AND symb_decoder(16#3a#)) OR
 					(reg_q896 AND symb_decoder(16#b1#)) OR
 					(reg_q896 AND symb_decoder(16#ef#)) OR
 					(reg_q896 AND symb_decoder(16#75#)) OR
 					(reg_q896 AND symb_decoder(16#09#)) OR
 					(reg_q896 AND symb_decoder(16#30#)) OR
 					(reg_q896 AND symb_decoder(16#53#)) OR
 					(reg_q896 AND symb_decoder(16#cf#)) OR
 					(reg_q896 AND symb_decoder(16#ce#)) OR
 					(reg_q896 AND symb_decoder(16#b9#)) OR
 					(reg_q896 AND symb_decoder(16#7b#)) OR
 					(reg_q896 AND symb_decoder(16#4a#)) OR
 					(reg_q896 AND symb_decoder(16#69#)) OR
 					(reg_q896 AND symb_decoder(16#97#)) OR
 					(reg_q896 AND symb_decoder(16#41#)) OR
 					(reg_q896 AND symb_decoder(16#1a#)) OR
 					(reg_q896 AND symb_decoder(16#44#)) OR
 					(reg_q896 AND symb_decoder(16#5a#)) OR
 					(reg_q896 AND symb_decoder(16#47#)) OR
 					(reg_q896 AND symb_decoder(16#d4#)) OR
 					(reg_q896 AND symb_decoder(16#e4#)) OR
 					(reg_q896 AND symb_decoder(16#bb#)) OR
 					(reg_q896 AND symb_decoder(16#84#)) OR
 					(reg_q896 AND symb_decoder(16#94#)) OR
 					(reg_q896 AND symb_decoder(16#13#)) OR
 					(reg_q896 AND symb_decoder(16#7a#)) OR
 					(reg_q896 AND symb_decoder(16#a8#)) OR
 					(reg_q896 AND symb_decoder(16#e8#)) OR
 					(reg_q896 AND symb_decoder(16#aa#)) OR
 					(reg_q896 AND symb_decoder(16#7d#)) OR
 					(reg_q896 AND symb_decoder(16#77#)) OR
 					(reg_q896 AND symb_decoder(16#f8#)) OR
 					(reg_q896 AND symb_decoder(16#86#)) OR
 					(reg_q896 AND symb_decoder(16#99#)) OR
 					(reg_q896 AND symb_decoder(16#9d#)) OR
 					(reg_q896 AND symb_decoder(16#e0#)) OR
 					(reg_q896 AND symb_decoder(16#a1#)) OR
 					(reg_q896 AND symb_decoder(16#f1#)) OR
 					(reg_q896 AND symb_decoder(16#0b#)) OR
 					(reg_q896 AND symb_decoder(16#31#)) OR
 					(reg_q896 AND symb_decoder(16#27#)) OR
 					(reg_q896 AND symb_decoder(16#0e#)) OR
 					(reg_q896 AND symb_decoder(16#a5#)) OR
 					(reg_q896 AND symb_decoder(16#bf#)) OR
 					(reg_q896 AND symb_decoder(16#63#)) OR
 					(reg_q896 AND symb_decoder(16#83#)) OR
 					(reg_q896 AND symb_decoder(16#04#)) OR
 					(reg_q896 AND symb_decoder(16#11#)) OR
 					(reg_q896 AND symb_decoder(16#ae#)) OR
 					(reg_q896 AND symb_decoder(16#64#)) OR
 					(reg_q896 AND symb_decoder(16#3d#)) OR
 					(reg_q896 AND symb_decoder(16#88#)) OR
 					(reg_q896 AND symb_decoder(16#b5#)) OR
 					(reg_q896 AND symb_decoder(16#b2#)) OR
 					(reg_q896 AND symb_decoder(16#67#)) OR
 					(reg_q896 AND symb_decoder(16#e3#)) OR
 					(reg_q896 AND symb_decoder(16#95#)) OR
 					(reg_q896 AND symb_decoder(16#68#)) OR
 					(reg_q896 AND symb_decoder(16#19#)) OR
 					(reg_q896 AND symb_decoder(16#61#)) OR
 					(reg_q896 AND symb_decoder(16#32#)) OR
 					(reg_q896 AND symb_decoder(16#e1#)) OR
 					(reg_q896 AND symb_decoder(16#1f#)) OR
 					(reg_q896 AND symb_decoder(16#0f#)) OR
 					(reg_q896 AND symb_decoder(16#23#)) OR
 					(reg_q896 AND symb_decoder(16#a9#)) OR
 					(reg_q896 AND symb_decoder(16#42#)) OR
 					(reg_q896 AND symb_decoder(16#b7#)) OR
 					(reg_q896 AND symb_decoder(16#b6#)) OR
 					(reg_q896 AND symb_decoder(16#5e#)) OR
 					(reg_q896 AND symb_decoder(16#ca#)) OR
 					(reg_q896 AND symb_decoder(16#eb#)) OR
 					(reg_q896 AND symb_decoder(16#3b#)) OR
 					(reg_q896 AND symb_decoder(16#a4#)) OR
 					(reg_q896 AND symb_decoder(16#2b#)) OR
 					(reg_q896 AND symb_decoder(16#6f#)) OR
 					(reg_q896 AND symb_decoder(16#22#)) OR
 					(reg_q896 AND symb_decoder(16#b3#)) OR
 					(reg_q896 AND symb_decoder(16#85#)) OR
 					(reg_q896 AND symb_decoder(16#62#)) OR
 					(reg_q896 AND symb_decoder(16#c7#)) OR
 					(reg_q896 AND symb_decoder(16#a2#)) OR
 					(reg_q896 AND symb_decoder(16#0c#)) OR
 					(reg_q896 AND symb_decoder(16#6a#)) OR
 					(reg_q896 AND symb_decoder(16#8c#)) OR
 					(reg_q896 AND symb_decoder(16#d9#)) OR
 					(reg_q896 AND symb_decoder(16#1d#)) OR
 					(reg_q896 AND symb_decoder(16#81#)) OR
 					(reg_q896 AND symb_decoder(16#8f#)) OR
 					(reg_q896 AND symb_decoder(16#db#)) OR
 					(reg_q896 AND symb_decoder(16#c8#)) OR
 					(reg_q896 AND symb_decoder(16#fb#)) OR
 					(reg_q896 AND symb_decoder(16#16#)) OR
 					(reg_q896 AND symb_decoder(16#07#)) OR
 					(reg_q896 AND symb_decoder(16#2e#)) OR
 					(reg_q896 AND symb_decoder(16#9b#)) OR
 					(reg_q896 AND symb_decoder(16#fa#)) OR
 					(reg_q896 AND symb_decoder(16#98#)) OR
 					(reg_q896 AND symb_decoder(16#de#)) OR
 					(reg_q896 AND symb_decoder(16#dc#)) OR
 					(reg_q896 AND symb_decoder(16#49#)) OR
 					(reg_q896 AND symb_decoder(16#89#)) OR
 					(reg_q896 AND symb_decoder(16#43#)) OR
 					(reg_q896 AND symb_decoder(16#b8#)) OR
 					(reg_q896 AND symb_decoder(16#f7#)) OR
 					(reg_q896 AND symb_decoder(16#06#)) OR
 					(reg_q896 AND symb_decoder(16#57#)) OR
 					(reg_q896 AND symb_decoder(16#21#)) OR
 					(reg_q896 AND symb_decoder(16#96#)) OR
 					(reg_q896 AND symb_decoder(16#d3#)) OR
 					(reg_q896 AND symb_decoder(16#20#)) OR
 					(reg_q896 AND symb_decoder(16#17#)) OR
 					(reg_q896 AND symb_decoder(16#d6#)) OR
 					(reg_q896 AND symb_decoder(16#be#)) OR
 					(reg_q896 AND symb_decoder(16#25#)) OR
 					(reg_q896 AND symb_decoder(16#51#)) OR
 					(reg_q896 AND symb_decoder(16#ad#)) OR
 					(reg_q896 AND symb_decoder(16#3f#)) OR
 					(reg_q896 AND symb_decoder(16#56#)) OR
 					(reg_q896 AND symb_decoder(16#65#)) OR
 					(reg_q896 AND symb_decoder(16#d8#)) OR
 					(reg_q896 AND symb_decoder(16#40#)) OR
 					(reg_q896 AND symb_decoder(16#6b#)) OR
 					(reg_q896 AND symb_decoder(16#a6#)) OR
 					(reg_q896 AND symb_decoder(16#7f#)) OR
 					(reg_q896 AND symb_decoder(16#93#)) OR
 					(reg_q896 AND symb_decoder(16#5b#)) OR
 					(reg_q896 AND symb_decoder(16#fd#)) OR
 					(reg_q896 AND symb_decoder(16#26#)) OR
 					(reg_q896 AND symb_decoder(16#6d#)) OR
 					(reg_q896 AND symb_decoder(16#1c#)) OR
 					(reg_q896 AND symb_decoder(16#e6#)) OR
 					(reg_q896 AND symb_decoder(16#c1#)) OR
 					(reg_q896 AND symb_decoder(16#9a#)) OR
 					(reg_q896 AND symb_decoder(16#50#)) OR
 					(reg_q896 AND symb_decoder(16#f6#)) OR
 					(reg_q896 AND symb_decoder(16#01#)) OR
 					(reg_q896 AND symb_decoder(16#8e#)) OR
 					(reg_q896 AND symb_decoder(16#9e#)) OR
 					(reg_q896 AND symb_decoder(16#d5#)) OR
 					(reg_q896 AND symb_decoder(16#af#)) OR
 					(reg_q896 AND symb_decoder(16#6c#)) OR
 					(reg_q896 AND symb_decoder(16#a7#)) OR
 					(reg_q896 AND symb_decoder(16#59#)) OR
 					(reg_q896 AND symb_decoder(16#7c#)) OR
 					(reg_q896 AND symb_decoder(16#f4#)) OR
 					(reg_q896 AND symb_decoder(16#73#)) OR
 					(reg_q896 AND symb_decoder(16#70#)) OR
 					(reg_q896 AND symb_decoder(16#c2#)) OR
 					(reg_q896 AND symb_decoder(16#ea#)) OR
 					(reg_q896 AND symb_decoder(16#48#)) OR
 					(reg_q896 AND symb_decoder(16#10#)) OR
 					(reg_q896 AND symb_decoder(16#8d#)) OR
 					(reg_q896 AND symb_decoder(16#c5#)) OR
 					(reg_q896 AND symb_decoder(16#2c#));
reg_q896_init <= '0' ;
	p_reg_q896: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q896 <= reg_q896_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q896 <= reg_q896_init;
        else
          reg_q896 <= reg_q896_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2000_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2000 AND symb_decoder(16#9b#)) OR
 					(reg_q2000 AND symb_decoder(16#a5#)) OR
 					(reg_q2000 AND symb_decoder(16#f7#)) OR
 					(reg_q2000 AND symb_decoder(16#d6#)) OR
 					(reg_q2000 AND symb_decoder(16#94#)) OR
 					(reg_q2000 AND symb_decoder(16#5a#)) OR
 					(reg_q2000 AND symb_decoder(16#b9#)) OR
 					(reg_q2000 AND symb_decoder(16#ac#)) OR
 					(reg_q2000 AND symb_decoder(16#46#)) OR
 					(reg_q2000 AND symb_decoder(16#ba#)) OR
 					(reg_q2000 AND symb_decoder(16#ce#)) OR
 					(reg_q2000 AND symb_decoder(16#ca#)) OR
 					(reg_q2000 AND symb_decoder(16#bb#)) OR
 					(reg_q2000 AND symb_decoder(16#88#)) OR
 					(reg_q2000 AND symb_decoder(16#2b#)) OR
 					(reg_q2000 AND symb_decoder(16#24#)) OR
 					(reg_q2000 AND symb_decoder(16#e3#)) OR
 					(reg_q2000 AND symb_decoder(16#63#)) OR
 					(reg_q2000 AND symb_decoder(16#d9#)) OR
 					(reg_q2000 AND symb_decoder(16#a9#)) OR
 					(reg_q2000 AND symb_decoder(16#a0#)) OR
 					(reg_q2000 AND symb_decoder(16#08#)) OR
 					(reg_q2000 AND symb_decoder(16#6b#)) OR
 					(reg_q2000 AND symb_decoder(16#6c#)) OR
 					(reg_q2000 AND symb_decoder(16#dc#)) OR
 					(reg_q2000 AND symb_decoder(16#01#)) OR
 					(reg_q2000 AND symb_decoder(16#e2#)) OR
 					(reg_q2000 AND symb_decoder(16#96#)) OR
 					(reg_q2000 AND symb_decoder(16#4e#)) OR
 					(reg_q2000 AND symb_decoder(16#32#)) OR
 					(reg_q2000 AND symb_decoder(16#33#)) OR
 					(reg_q2000 AND symb_decoder(16#15#)) OR
 					(reg_q2000 AND symb_decoder(16#c2#)) OR
 					(reg_q2000 AND symb_decoder(16#48#)) OR
 					(reg_q2000 AND symb_decoder(16#b5#)) OR
 					(reg_q2000 AND symb_decoder(16#b7#)) OR
 					(reg_q2000 AND symb_decoder(16#b4#)) OR
 					(reg_q2000 AND symb_decoder(16#e5#)) OR
 					(reg_q2000 AND symb_decoder(16#66#)) OR
 					(reg_q2000 AND symb_decoder(16#ec#)) OR
 					(reg_q2000 AND symb_decoder(16#d3#)) OR
 					(reg_q2000 AND symb_decoder(16#39#)) OR
 					(reg_q2000 AND symb_decoder(16#d4#)) OR
 					(reg_q2000 AND symb_decoder(16#be#)) OR
 					(reg_q2000 AND symb_decoder(16#0b#)) OR
 					(reg_q2000 AND symb_decoder(16#de#)) OR
 					(reg_q2000 AND symb_decoder(16#07#)) OR
 					(reg_q2000 AND symb_decoder(16#ae#)) OR
 					(reg_q2000 AND symb_decoder(16#db#)) OR
 					(reg_q2000 AND symb_decoder(16#76#)) OR
 					(reg_q2000 AND symb_decoder(16#7e#)) OR
 					(reg_q2000 AND symb_decoder(16#c4#)) OR
 					(reg_q2000 AND symb_decoder(16#77#)) OR
 					(reg_q2000 AND symb_decoder(16#69#)) OR
 					(reg_q2000 AND symb_decoder(16#25#)) OR
 					(reg_q2000 AND symb_decoder(16#a8#)) OR
 					(reg_q2000 AND symb_decoder(16#7f#)) OR
 					(reg_q2000 AND symb_decoder(16#84#)) OR
 					(reg_q2000 AND symb_decoder(16#c7#)) OR
 					(reg_q2000 AND symb_decoder(16#a1#)) OR
 					(reg_q2000 AND symb_decoder(16#5b#)) OR
 					(reg_q2000 AND symb_decoder(16#0f#)) OR
 					(reg_q2000 AND symb_decoder(16#8e#)) OR
 					(reg_q2000 AND symb_decoder(16#22#)) OR
 					(reg_q2000 AND symb_decoder(16#e8#)) OR
 					(reg_q2000 AND symb_decoder(16#3a#)) OR
 					(reg_q2000 AND symb_decoder(16#f6#)) OR
 					(reg_q2000 AND symb_decoder(16#53#)) OR
 					(reg_q2000 AND symb_decoder(16#5f#)) OR
 					(reg_q2000 AND symb_decoder(16#fd#)) OR
 					(reg_q2000 AND symb_decoder(16#04#)) OR
 					(reg_q2000 AND symb_decoder(16#93#)) OR
 					(reg_q2000 AND symb_decoder(16#2e#)) OR
 					(reg_q2000 AND symb_decoder(16#06#)) OR
 					(reg_q2000 AND symb_decoder(16#3b#)) OR
 					(reg_q2000 AND symb_decoder(16#f1#)) OR
 					(reg_q2000 AND symb_decoder(16#c8#)) OR
 					(reg_q2000 AND symb_decoder(16#0a#)) OR
 					(reg_q2000 AND symb_decoder(16#a4#)) OR
 					(reg_q2000 AND symb_decoder(16#95#)) OR
 					(reg_q2000 AND symb_decoder(16#98#)) OR
 					(reg_q2000 AND symb_decoder(16#8d#)) OR
 					(reg_q2000 AND symb_decoder(16#0d#)) OR
 					(reg_q2000 AND symb_decoder(16#6a#)) OR
 					(reg_q2000 AND symb_decoder(16#43#)) OR
 					(reg_q2000 AND symb_decoder(16#67#)) OR
 					(reg_q2000 AND symb_decoder(16#91#)) OR
 					(reg_q2000 AND symb_decoder(16#fb#)) OR
 					(reg_q2000 AND symb_decoder(16#70#)) OR
 					(reg_q2000 AND symb_decoder(16#47#)) OR
 					(reg_q2000 AND symb_decoder(16#71#)) OR
 					(reg_q2000 AND symb_decoder(16#44#)) OR
 					(reg_q2000 AND symb_decoder(16#9a#)) OR
 					(reg_q2000 AND symb_decoder(16#fa#)) OR
 					(reg_q2000 AND symb_decoder(16#d2#)) OR
 					(reg_q2000 AND symb_decoder(16#a7#)) OR
 					(reg_q2000 AND symb_decoder(16#75#)) OR
 					(reg_q2000 AND symb_decoder(16#73#)) OR
 					(reg_q2000 AND symb_decoder(16#cd#)) OR
 					(reg_q2000 AND symb_decoder(16#54#)) OR
 					(reg_q2000 AND symb_decoder(16#0c#)) OR
 					(reg_q2000 AND symb_decoder(16#f0#)) OR
 					(reg_q2000 AND symb_decoder(16#b0#)) OR
 					(reg_q2000 AND symb_decoder(16#74#)) OR
 					(reg_q2000 AND symb_decoder(16#00#)) OR
 					(reg_q2000 AND symb_decoder(16#03#)) OR
 					(reg_q2000 AND symb_decoder(16#92#)) OR
 					(reg_q2000 AND symb_decoder(16#c1#)) OR
 					(reg_q2000 AND symb_decoder(16#9f#)) OR
 					(reg_q2000 AND symb_decoder(16#51#)) OR
 					(reg_q2000 AND symb_decoder(16#2d#)) OR
 					(reg_q2000 AND symb_decoder(16#d1#)) OR
 					(reg_q2000 AND symb_decoder(16#af#)) OR
 					(reg_q2000 AND symb_decoder(16#11#)) OR
 					(reg_q2000 AND symb_decoder(16#3c#)) OR
 					(reg_q2000 AND symb_decoder(16#41#)) OR
 					(reg_q2000 AND symb_decoder(16#da#)) OR
 					(reg_q2000 AND symb_decoder(16#3d#)) OR
 					(reg_q2000 AND symb_decoder(16#9c#)) OR
 					(reg_q2000 AND symb_decoder(16#42#)) OR
 					(reg_q2000 AND symb_decoder(16#68#)) OR
 					(reg_q2000 AND symb_decoder(16#5c#)) OR
 					(reg_q2000 AND symb_decoder(16#1a#)) OR
 					(reg_q2000 AND symb_decoder(16#8c#)) OR
 					(reg_q2000 AND symb_decoder(16#35#)) OR
 					(reg_q2000 AND symb_decoder(16#4a#)) OR
 					(reg_q2000 AND symb_decoder(16#bf#)) OR
 					(reg_q2000 AND symb_decoder(16#4d#)) OR
 					(reg_q2000 AND symb_decoder(16#ef#)) OR
 					(reg_q2000 AND symb_decoder(16#55#)) OR
 					(reg_q2000 AND symb_decoder(16#2a#)) OR
 					(reg_q2000 AND symb_decoder(16#56#)) OR
 					(reg_q2000 AND symb_decoder(16#50#)) OR
 					(reg_q2000 AND symb_decoder(16#4c#)) OR
 					(reg_q2000 AND symb_decoder(16#c6#)) OR
 					(reg_q2000 AND symb_decoder(16#16#)) OR
 					(reg_q2000 AND symb_decoder(16#89#)) OR
 					(reg_q2000 AND symb_decoder(16#3f#)) OR
 					(reg_q2000 AND symb_decoder(16#c5#)) OR
 					(reg_q2000 AND symb_decoder(16#59#)) OR
 					(reg_q2000 AND symb_decoder(16#d0#)) OR
 					(reg_q2000 AND symb_decoder(16#7b#)) OR
 					(reg_q2000 AND symb_decoder(16#65#)) OR
 					(reg_q2000 AND symb_decoder(16#cf#)) OR
 					(reg_q2000 AND symb_decoder(16#37#)) OR
 					(reg_q2000 AND symb_decoder(16#17#)) OR
 					(reg_q2000 AND symb_decoder(16#4f#)) OR
 					(reg_q2000 AND symb_decoder(16#f3#)) OR
 					(reg_q2000 AND symb_decoder(16#5e#)) OR
 					(reg_q2000 AND symb_decoder(16#7d#)) OR
 					(reg_q2000 AND symb_decoder(16#38#)) OR
 					(reg_q2000 AND symb_decoder(16#dd#)) OR
 					(reg_q2000 AND symb_decoder(16#bd#)) OR
 					(reg_q2000 AND symb_decoder(16#e0#)) OR
 					(reg_q2000 AND symb_decoder(16#a3#)) OR
 					(reg_q2000 AND symb_decoder(16#9e#)) OR
 					(reg_q2000 AND symb_decoder(16#e4#)) OR
 					(reg_q2000 AND symb_decoder(16#21#)) OR
 					(reg_q2000 AND symb_decoder(16#23#)) OR
 					(reg_q2000 AND symb_decoder(16#97#)) OR
 					(reg_q2000 AND symb_decoder(16#12#)) OR
 					(reg_q2000 AND symb_decoder(16#09#)) OR
 					(reg_q2000 AND symb_decoder(16#36#)) OR
 					(reg_q2000 AND symb_decoder(16#df#)) OR
 					(reg_q2000 AND symb_decoder(16#18#)) OR
 					(reg_q2000 AND symb_decoder(16#6d#)) OR
 					(reg_q2000 AND symb_decoder(16#30#)) OR
 					(reg_q2000 AND symb_decoder(16#05#)) OR
 					(reg_q2000 AND symb_decoder(16#d7#)) OR
 					(reg_q2000 AND symb_decoder(16#99#)) OR
 					(reg_q2000 AND symb_decoder(16#78#)) OR
 					(reg_q2000 AND symb_decoder(16#cc#)) OR
 					(reg_q2000 AND symb_decoder(16#e7#)) OR
 					(reg_q2000 AND symb_decoder(16#d5#)) OR
 					(reg_q2000 AND symb_decoder(16#72#)) OR
 					(reg_q2000 AND symb_decoder(16#40#)) OR
 					(reg_q2000 AND symb_decoder(16#27#)) OR
 					(reg_q2000 AND symb_decoder(16#5d#)) OR
 					(reg_q2000 AND symb_decoder(16#7c#)) OR
 					(reg_q2000 AND symb_decoder(16#b8#)) OR
 					(reg_q2000 AND symb_decoder(16#aa#)) OR
 					(reg_q2000 AND symb_decoder(16#d8#)) OR
 					(reg_q2000 AND symb_decoder(16#31#)) OR
 					(reg_q2000 AND symb_decoder(16#b1#)) OR
 					(reg_q2000 AND symb_decoder(16#90#)) OR
 					(reg_q2000 AND symb_decoder(16#14#)) OR
 					(reg_q2000 AND symb_decoder(16#1e#)) OR
 					(reg_q2000 AND symb_decoder(16#1d#)) OR
 					(reg_q2000 AND symb_decoder(16#b6#)) OR
 					(reg_q2000 AND symb_decoder(16#1b#)) OR
 					(reg_q2000 AND symb_decoder(16#eb#)) OR
 					(reg_q2000 AND symb_decoder(16#85#)) OR
 					(reg_q2000 AND symb_decoder(16#e1#)) OR
 					(reg_q2000 AND symb_decoder(16#0e#)) OR
 					(reg_q2000 AND symb_decoder(16#f4#)) OR
 					(reg_q2000 AND symb_decoder(16#8f#)) OR
 					(reg_q2000 AND symb_decoder(16#8a#)) OR
 					(reg_q2000 AND symb_decoder(16#58#)) OR
 					(reg_q2000 AND symb_decoder(16#7a#)) OR
 					(reg_q2000 AND symb_decoder(16#ff#)) OR
 					(reg_q2000 AND symb_decoder(16#f8#)) OR
 					(reg_q2000 AND symb_decoder(16#ee#)) OR
 					(reg_q2000 AND symb_decoder(16#61#)) OR
 					(reg_q2000 AND symb_decoder(16#34#)) OR
 					(reg_q2000 AND symb_decoder(16#81#)) OR
 					(reg_q2000 AND symb_decoder(16#4b#)) OR
 					(reg_q2000 AND symb_decoder(16#52#)) OR
 					(reg_q2000 AND symb_decoder(16#c9#)) OR
 					(reg_q2000 AND symb_decoder(16#45#)) OR
 					(reg_q2000 AND symb_decoder(16#82#)) OR
 					(reg_q2000 AND symb_decoder(16#b2#)) OR
 					(reg_q2000 AND symb_decoder(16#57#)) OR
 					(reg_q2000 AND symb_decoder(16#2c#)) OR
 					(reg_q2000 AND symb_decoder(16#e6#)) OR
 					(reg_q2000 AND symb_decoder(16#6f#)) OR
 					(reg_q2000 AND symb_decoder(16#64#)) OR
 					(reg_q2000 AND symb_decoder(16#8b#)) OR
 					(reg_q2000 AND symb_decoder(16#ad#)) OR
 					(reg_q2000 AND symb_decoder(16#ea#)) OR
 					(reg_q2000 AND symb_decoder(16#49#)) OR
 					(reg_q2000 AND symb_decoder(16#80#)) OR
 					(reg_q2000 AND symb_decoder(16#87#)) OR
 					(reg_q2000 AND symb_decoder(16#1c#)) OR
 					(reg_q2000 AND symb_decoder(16#20#)) OR
 					(reg_q2000 AND symb_decoder(16#6e#)) OR
 					(reg_q2000 AND symb_decoder(16#2f#)) OR
 					(reg_q2000 AND symb_decoder(16#3e#)) OR
 					(reg_q2000 AND symb_decoder(16#60#)) OR
 					(reg_q2000 AND symb_decoder(16#cb#)) OR
 					(reg_q2000 AND symb_decoder(16#1f#)) OR
 					(reg_q2000 AND symb_decoder(16#79#)) OR
 					(reg_q2000 AND symb_decoder(16#28#)) OR
 					(reg_q2000 AND symb_decoder(16#c0#)) OR
 					(reg_q2000 AND symb_decoder(16#f9#)) OR
 					(reg_q2000 AND symb_decoder(16#a2#)) OR
 					(reg_q2000 AND symb_decoder(16#19#)) OR
 					(reg_q2000 AND symb_decoder(16#ed#)) OR
 					(reg_q2000 AND symb_decoder(16#f2#)) OR
 					(reg_q2000 AND symb_decoder(16#02#)) OR
 					(reg_q2000 AND symb_decoder(16#62#)) OR
 					(reg_q2000 AND symb_decoder(16#b3#)) OR
 					(reg_q2000 AND symb_decoder(16#83#)) OR
 					(reg_q2000 AND symb_decoder(16#f5#)) OR
 					(reg_q2000 AND symb_decoder(16#e9#)) OR
 					(reg_q2000 AND symb_decoder(16#fc#)) OR
 					(reg_q2000 AND symb_decoder(16#fe#)) OR
 					(reg_q2000 AND symb_decoder(16#13#)) OR
 					(reg_q2000 AND symb_decoder(16#c3#)) OR
 					(reg_q2000 AND symb_decoder(16#bc#)) OR
 					(reg_q2000 AND symb_decoder(16#ab#)) OR
 					(reg_q2000 AND symb_decoder(16#29#)) OR
 					(reg_q2000 AND symb_decoder(16#10#)) OR
 					(reg_q2000 AND symb_decoder(16#9d#)) OR
 					(reg_q2000 AND symb_decoder(16#86#)) OR
 					(reg_q2000 AND symb_decoder(16#a6#)) OR
 					(reg_q2000 AND symb_decoder(16#26#));
reg_q2000_init <= '0' ;
	p_reg_q2000: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2000 <= reg_q2000_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2000 <= reg_q2000_init;
        else
          reg_q2000 <= reg_q2000_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2533_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2533 AND symb_decoder(16#18#)) OR
 					(reg_q2533 AND symb_decoder(16#52#)) OR
 					(reg_q2533 AND symb_decoder(16#78#)) OR
 					(reg_q2533 AND symb_decoder(16#15#)) OR
 					(reg_q2533 AND symb_decoder(16#42#)) OR
 					(reg_q2533 AND symb_decoder(16#43#)) OR
 					(reg_q2533 AND symb_decoder(16#90#)) OR
 					(reg_q2533 AND symb_decoder(16#82#)) OR
 					(reg_q2533 AND symb_decoder(16#05#)) OR
 					(reg_q2533 AND symb_decoder(16#11#)) OR
 					(reg_q2533 AND symb_decoder(16#b9#)) OR
 					(reg_q2533 AND symb_decoder(16#58#)) OR
 					(reg_q2533 AND symb_decoder(16#5d#)) OR
 					(reg_q2533 AND symb_decoder(16#92#)) OR
 					(reg_q2533 AND symb_decoder(16#5a#)) OR
 					(reg_q2533 AND symb_decoder(16#1b#)) OR
 					(reg_q2533 AND symb_decoder(16#b6#)) OR
 					(reg_q2533 AND symb_decoder(16#bf#)) OR
 					(reg_q2533 AND symb_decoder(16#2b#)) OR
 					(reg_q2533 AND symb_decoder(16#ad#)) OR
 					(reg_q2533 AND symb_decoder(16#22#)) OR
 					(reg_q2533 AND symb_decoder(16#60#)) OR
 					(reg_q2533 AND symb_decoder(16#dd#)) OR
 					(reg_q2533 AND symb_decoder(16#63#)) OR
 					(reg_q2533 AND symb_decoder(16#f9#)) OR
 					(reg_q2533 AND symb_decoder(16#1f#)) OR
 					(reg_q2533 AND symb_decoder(16#24#)) OR
 					(reg_q2533 AND symb_decoder(16#e5#)) OR
 					(reg_q2533 AND symb_decoder(16#ee#)) OR
 					(reg_q2533 AND symb_decoder(16#4c#)) OR
 					(reg_q2533 AND symb_decoder(16#6a#)) OR
 					(reg_q2533 AND symb_decoder(16#84#)) OR
 					(reg_q2533 AND symb_decoder(16#7a#)) OR
 					(reg_q2533 AND symb_decoder(16#55#)) OR
 					(reg_q2533 AND symb_decoder(16#8f#)) OR
 					(reg_q2533 AND symb_decoder(16#46#)) OR
 					(reg_q2533 AND symb_decoder(16#aa#)) OR
 					(reg_q2533 AND symb_decoder(16#9c#)) OR
 					(reg_q2533 AND symb_decoder(16#c3#)) OR
 					(reg_q2533 AND symb_decoder(16#f5#)) OR
 					(reg_q2533 AND symb_decoder(16#3c#)) OR
 					(reg_q2533 AND symb_decoder(16#c8#)) OR
 					(reg_q2533 AND symb_decoder(16#49#)) OR
 					(reg_q2533 AND symb_decoder(16#98#)) OR
 					(reg_q2533 AND symb_decoder(16#e1#)) OR
 					(reg_q2533 AND symb_decoder(16#2c#)) OR
 					(reg_q2533 AND symb_decoder(16#e4#)) OR
 					(reg_q2533 AND symb_decoder(16#0e#)) OR
 					(reg_q2533 AND symb_decoder(16#4a#)) OR
 					(reg_q2533 AND symb_decoder(16#da#)) OR
 					(reg_q2533 AND symb_decoder(16#f0#)) OR
 					(reg_q2533 AND symb_decoder(16#59#)) OR
 					(reg_q2533 AND symb_decoder(16#02#)) OR
 					(reg_q2533 AND symb_decoder(16#30#)) OR
 					(reg_q2533 AND symb_decoder(16#03#)) OR
 					(reg_q2533 AND symb_decoder(16#fa#)) OR
 					(reg_q2533 AND symb_decoder(16#ab#)) OR
 					(reg_q2533 AND symb_decoder(16#cc#)) OR
 					(reg_q2533 AND symb_decoder(16#51#)) OR
 					(reg_q2533 AND symb_decoder(16#0f#)) OR
 					(reg_q2533 AND symb_decoder(16#d7#)) OR
 					(reg_q2533 AND symb_decoder(16#b8#)) OR
 					(reg_q2533 AND symb_decoder(16#ca#)) OR
 					(reg_q2533 AND symb_decoder(16#a7#)) OR
 					(reg_q2533 AND symb_decoder(16#0d#)) OR
 					(reg_q2533 AND symb_decoder(16#85#)) OR
 					(reg_q2533 AND symb_decoder(16#6c#)) OR
 					(reg_q2533 AND symb_decoder(16#7d#)) OR
 					(reg_q2533 AND symb_decoder(16#9e#)) OR
 					(reg_q2533 AND symb_decoder(16#ea#)) OR
 					(reg_q2533 AND symb_decoder(16#3f#)) OR
 					(reg_q2533 AND symb_decoder(16#17#)) OR
 					(reg_q2533 AND symb_decoder(16#a0#)) OR
 					(reg_q2533 AND symb_decoder(16#95#)) OR
 					(reg_q2533 AND symb_decoder(16#54#)) OR
 					(reg_q2533 AND symb_decoder(16#cd#)) OR
 					(reg_q2533 AND symb_decoder(16#06#)) OR
 					(reg_q2533 AND symb_decoder(16#d0#)) OR
 					(reg_q2533 AND symb_decoder(16#19#)) OR
 					(reg_q2533 AND symb_decoder(16#09#)) OR
 					(reg_q2533 AND symb_decoder(16#70#)) OR
 					(reg_q2533 AND symb_decoder(16#08#)) OR
 					(reg_q2533 AND symb_decoder(16#99#)) OR
 					(reg_q2533 AND symb_decoder(16#f4#)) OR
 					(reg_q2533 AND symb_decoder(16#20#)) OR
 					(reg_q2533 AND symb_decoder(16#45#)) OR
 					(reg_q2533 AND symb_decoder(16#e3#)) OR
 					(reg_q2533 AND symb_decoder(16#c7#)) OR
 					(reg_q2533 AND symb_decoder(16#29#)) OR
 					(reg_q2533 AND symb_decoder(16#79#)) OR
 					(reg_q2533 AND symb_decoder(16#21#)) OR
 					(reg_q2533 AND symb_decoder(16#c4#)) OR
 					(reg_q2533 AND symb_decoder(16#8d#)) OR
 					(reg_q2533 AND symb_decoder(16#34#)) OR
 					(reg_q2533 AND symb_decoder(16#dc#)) OR
 					(reg_q2533 AND symb_decoder(16#33#)) OR
 					(reg_q2533 AND symb_decoder(16#3d#)) OR
 					(reg_q2533 AND symb_decoder(16#07#)) OR
 					(reg_q2533 AND symb_decoder(16#7b#)) OR
 					(reg_q2533 AND symb_decoder(16#80#)) OR
 					(reg_q2533 AND symb_decoder(16#c6#)) OR
 					(reg_q2533 AND symb_decoder(16#9a#)) OR
 					(reg_q2533 AND symb_decoder(16#5e#)) OR
 					(reg_q2533 AND symb_decoder(16#14#)) OR
 					(reg_q2533 AND symb_decoder(16#39#)) OR
 					(reg_q2533 AND symb_decoder(16#38#)) OR
 					(reg_q2533 AND symb_decoder(16#56#)) OR
 					(reg_q2533 AND symb_decoder(16#4f#)) OR
 					(reg_q2533 AND symb_decoder(16#66#)) OR
 					(reg_q2533 AND symb_decoder(16#1a#)) OR
 					(reg_q2533 AND symb_decoder(16#5f#)) OR
 					(reg_q2533 AND symb_decoder(16#ac#)) OR
 					(reg_q2533 AND symb_decoder(16#0b#)) OR
 					(reg_q2533 AND symb_decoder(16#9d#)) OR
 					(reg_q2533 AND symb_decoder(16#1c#)) OR
 					(reg_q2533 AND symb_decoder(16#f3#)) OR
 					(reg_q2533 AND symb_decoder(16#0a#)) OR
 					(reg_q2533 AND symb_decoder(16#a3#)) OR
 					(reg_q2533 AND symb_decoder(16#35#)) OR
 					(reg_q2533 AND symb_decoder(16#27#)) OR
 					(reg_q2533 AND symb_decoder(16#7f#)) OR
 					(reg_q2533 AND symb_decoder(16#69#)) OR
 					(reg_q2533 AND symb_decoder(16#b7#)) OR
 					(reg_q2533 AND symb_decoder(16#36#)) OR
 					(reg_q2533 AND symb_decoder(16#2e#)) OR
 					(reg_q2533 AND symb_decoder(16#71#)) OR
 					(reg_q2533 AND symb_decoder(16#f8#)) OR
 					(reg_q2533 AND symb_decoder(16#b2#)) OR
 					(reg_q2533 AND symb_decoder(16#a8#)) OR
 					(reg_q2533 AND symb_decoder(16#d8#)) OR
 					(reg_q2533 AND symb_decoder(16#2f#)) OR
 					(reg_q2533 AND symb_decoder(16#23#)) OR
 					(reg_q2533 AND symb_decoder(16#db#)) OR
 					(reg_q2533 AND symb_decoder(16#13#)) OR
 					(reg_q2533 AND symb_decoder(16#c0#)) OR
 					(reg_q2533 AND symb_decoder(16#4b#)) OR
 					(reg_q2533 AND symb_decoder(16#c2#)) OR
 					(reg_q2533 AND symb_decoder(16#d9#)) OR
 					(reg_q2533 AND symb_decoder(16#88#)) OR
 					(reg_q2533 AND symb_decoder(16#bb#)) OR
 					(reg_q2533 AND symb_decoder(16#a1#)) OR
 					(reg_q2533 AND symb_decoder(16#1d#)) OR
 					(reg_q2533 AND symb_decoder(16#4d#)) OR
 					(reg_q2533 AND symb_decoder(16#48#)) OR
 					(reg_q2533 AND symb_decoder(16#a9#)) OR
 					(reg_q2533 AND symb_decoder(16#12#)) OR
 					(reg_q2533 AND symb_decoder(16#41#)) OR
 					(reg_q2533 AND symb_decoder(16#93#)) OR
 					(reg_q2533 AND symb_decoder(16#fe#)) OR
 					(reg_q2533 AND symb_decoder(16#d1#)) OR
 					(reg_q2533 AND symb_decoder(16#e7#)) OR
 					(reg_q2533 AND symb_decoder(16#c5#)) OR
 					(reg_q2533 AND symb_decoder(16#91#)) OR
 					(reg_q2533 AND symb_decoder(16#f6#)) OR
 					(reg_q2533 AND symb_decoder(16#fc#)) OR
 					(reg_q2533 AND symb_decoder(16#64#)) OR
 					(reg_q2533 AND symb_decoder(16#67#)) OR
 					(reg_q2533 AND symb_decoder(16#83#)) OR
 					(reg_q2533 AND symb_decoder(16#28#)) OR
 					(reg_q2533 AND symb_decoder(16#a6#)) OR
 					(reg_q2533 AND symb_decoder(16#8e#)) OR
 					(reg_q2533 AND symb_decoder(16#e2#)) OR
 					(reg_q2533 AND symb_decoder(16#01#)) OR
 					(reg_q2533 AND symb_decoder(16#76#)) OR
 					(reg_q2533 AND symb_decoder(16#65#)) OR
 					(reg_q2533 AND symb_decoder(16#ae#)) OR
 					(reg_q2533 AND symb_decoder(16#bd#)) OR
 					(reg_q2533 AND symb_decoder(16#87#)) OR
 					(reg_q2533 AND symb_decoder(16#6f#)) OR
 					(reg_q2533 AND symb_decoder(16#1e#)) OR
 					(reg_q2533 AND symb_decoder(16#73#)) OR
 					(reg_q2533 AND symb_decoder(16#6e#)) OR
 					(reg_q2533 AND symb_decoder(16#ff#)) OR
 					(reg_q2533 AND symb_decoder(16#f2#)) OR
 					(reg_q2533 AND symb_decoder(16#4e#)) OR
 					(reg_q2533 AND symb_decoder(16#8b#)) OR
 					(reg_q2533 AND symb_decoder(16#96#)) OR
 					(reg_q2533 AND symb_decoder(16#86#)) OR
 					(reg_q2533 AND symb_decoder(16#e9#)) OR
 					(reg_q2533 AND symb_decoder(16#f7#)) OR
 					(reg_q2533 AND symb_decoder(16#40#)) OR
 					(reg_q2533 AND symb_decoder(16#ec#)) OR
 					(reg_q2533 AND symb_decoder(16#cf#)) OR
 					(reg_q2533 AND symb_decoder(16#7c#)) OR
 					(reg_q2533 AND symb_decoder(16#c1#)) OR
 					(reg_q2533 AND symb_decoder(16#77#)) OR
 					(reg_q2533 AND symb_decoder(16#81#)) OR
 					(reg_q2533 AND symb_decoder(16#10#)) OR
 					(reg_q2533 AND symb_decoder(16#fb#)) OR
 					(reg_q2533 AND symb_decoder(16#53#)) OR
 					(reg_q2533 AND symb_decoder(16#8a#)) OR
 					(reg_q2533 AND symb_decoder(16#74#)) OR
 					(reg_q2533 AND symb_decoder(16#26#)) OR
 					(reg_q2533 AND symb_decoder(16#f1#)) OR
 					(reg_q2533 AND symb_decoder(16#97#)) OR
 					(reg_q2533 AND symb_decoder(16#61#)) OR
 					(reg_q2533 AND symb_decoder(16#a2#)) OR
 					(reg_q2533 AND symb_decoder(16#ef#)) OR
 					(reg_q2533 AND symb_decoder(16#5b#)) OR
 					(reg_q2533 AND symb_decoder(16#de#)) OR
 					(reg_q2533 AND symb_decoder(16#0c#)) OR
 					(reg_q2533 AND symb_decoder(16#44#)) OR
 					(reg_q2533 AND symb_decoder(16#fd#)) OR
 					(reg_q2533 AND symb_decoder(16#b1#)) OR
 					(reg_q2533 AND symb_decoder(16#eb#)) OR
 					(reg_q2533 AND symb_decoder(16#e6#)) OR
 					(reg_q2533 AND symb_decoder(16#47#)) OR
 					(reg_q2533 AND symb_decoder(16#df#)) OR
 					(reg_q2533 AND symb_decoder(16#a5#)) OR
 					(reg_q2533 AND symb_decoder(16#e0#)) OR
 					(reg_q2533 AND symb_decoder(16#72#)) OR
 					(reg_q2533 AND symb_decoder(16#2d#)) OR
 					(reg_q2533 AND symb_decoder(16#89#)) OR
 					(reg_q2533 AND symb_decoder(16#6b#)) OR
 					(reg_q2533 AND symb_decoder(16#31#)) OR
 					(reg_q2533 AND symb_decoder(16#b3#)) OR
 					(reg_q2533 AND symb_decoder(16#6d#)) OR
 					(reg_q2533 AND symb_decoder(16#ba#)) OR
 					(reg_q2533 AND symb_decoder(16#bc#)) OR
 					(reg_q2533 AND symb_decoder(16#c9#)) OR
 					(reg_q2533 AND symb_decoder(16#57#)) OR
 					(reg_q2533 AND symb_decoder(16#d3#)) OR
 					(reg_q2533 AND symb_decoder(16#62#)) OR
 					(reg_q2533 AND symb_decoder(16#5c#)) OR
 					(reg_q2533 AND symb_decoder(16#cb#)) OR
 					(reg_q2533 AND symb_decoder(16#3a#)) OR
 					(reg_q2533 AND symb_decoder(16#32#)) OR
 					(reg_q2533 AND symb_decoder(16#d6#)) OR
 					(reg_q2533 AND symb_decoder(16#b0#)) OR
 					(reg_q2533 AND symb_decoder(16#2a#)) OR
 					(reg_q2533 AND symb_decoder(16#a4#)) OR
 					(reg_q2533 AND symb_decoder(16#d4#)) OR
 					(reg_q2533 AND symb_decoder(16#3e#)) OR
 					(reg_q2533 AND symb_decoder(16#b5#)) OR
 					(reg_q2533 AND symb_decoder(16#ed#)) OR
 					(reg_q2533 AND symb_decoder(16#3b#)) OR
 					(reg_q2533 AND symb_decoder(16#7e#)) OR
 					(reg_q2533 AND symb_decoder(16#b4#)) OR
 					(reg_q2533 AND symb_decoder(16#16#)) OR
 					(reg_q2533 AND symb_decoder(16#ce#)) OR
 					(reg_q2533 AND symb_decoder(16#af#)) OR
 					(reg_q2533 AND symb_decoder(16#8c#)) OR
 					(reg_q2533 AND symb_decoder(16#e8#)) OR
 					(reg_q2533 AND symb_decoder(16#94#)) OR
 					(reg_q2533 AND symb_decoder(16#37#)) OR
 					(reg_q2533 AND symb_decoder(16#d5#)) OR
 					(reg_q2533 AND symb_decoder(16#68#)) OR
 					(reg_q2533 AND symb_decoder(16#d2#)) OR
 					(reg_q2533 AND symb_decoder(16#04#)) OR
 					(reg_q2533 AND symb_decoder(16#be#)) OR
 					(reg_q2533 AND symb_decoder(16#9f#)) OR
 					(reg_q2533 AND symb_decoder(16#75#)) OR
 					(reg_q2533 AND symb_decoder(16#25#)) OR
 					(reg_q2533 AND symb_decoder(16#50#)) OR
 					(reg_q2533 AND symb_decoder(16#9b#)) OR
 					(reg_q2533 AND symb_decoder(16#00#));
reg_q2533_init <= '0' ;
	p_reg_q2533: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2533 <= reg_q2533_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2533 <= reg_q2533_init;
        else
          reg_q2533 <= reg_q2533_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q303_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q303 AND symb_decoder(16#37#)) OR
 					(reg_q303 AND symb_decoder(16#24#)) OR
 					(reg_q303 AND symb_decoder(16#b8#)) OR
 					(reg_q303 AND symb_decoder(16#3a#)) OR
 					(reg_q303 AND symb_decoder(16#f2#)) OR
 					(reg_q303 AND symb_decoder(16#9a#)) OR
 					(reg_q303 AND symb_decoder(16#78#)) OR
 					(reg_q303 AND symb_decoder(16#d8#)) OR
 					(reg_q303 AND symb_decoder(16#89#)) OR
 					(reg_q303 AND symb_decoder(16#eb#)) OR
 					(reg_q303 AND symb_decoder(16#a1#)) OR
 					(reg_q303 AND symb_decoder(16#43#)) OR
 					(reg_q303 AND symb_decoder(16#7f#)) OR
 					(reg_q303 AND symb_decoder(16#c7#)) OR
 					(reg_q303 AND symb_decoder(16#d9#)) OR
 					(reg_q303 AND symb_decoder(16#b3#)) OR
 					(reg_q303 AND symb_decoder(16#f9#)) OR
 					(reg_q303 AND symb_decoder(16#3c#)) OR
 					(reg_q303 AND symb_decoder(16#de#)) OR
 					(reg_q303 AND symb_decoder(16#e4#)) OR
 					(reg_q303 AND symb_decoder(16#07#)) OR
 					(reg_q303 AND symb_decoder(16#7c#)) OR
 					(reg_q303 AND symb_decoder(16#33#)) OR
 					(reg_q303 AND symb_decoder(16#be#)) OR
 					(reg_q303 AND symb_decoder(16#50#)) OR
 					(reg_q303 AND symb_decoder(16#27#)) OR
 					(reg_q303 AND symb_decoder(16#1b#)) OR
 					(reg_q303 AND symb_decoder(16#55#)) OR
 					(reg_q303 AND symb_decoder(16#03#)) OR
 					(reg_q303 AND symb_decoder(16#09#)) OR
 					(reg_q303 AND symb_decoder(16#82#)) OR
 					(reg_q303 AND symb_decoder(16#5d#)) OR
 					(reg_q303 AND symb_decoder(16#7d#)) OR
 					(reg_q303 AND symb_decoder(16#96#)) OR
 					(reg_q303 AND symb_decoder(16#90#)) OR
 					(reg_q303 AND symb_decoder(16#52#)) OR
 					(reg_q303 AND symb_decoder(16#94#)) OR
 					(reg_q303 AND symb_decoder(16#16#)) OR
 					(reg_q303 AND symb_decoder(16#7a#)) OR
 					(reg_q303 AND symb_decoder(16#42#)) OR
 					(reg_q303 AND symb_decoder(16#1f#)) OR
 					(reg_q303 AND symb_decoder(16#71#)) OR
 					(reg_q303 AND symb_decoder(16#4a#)) OR
 					(reg_q303 AND symb_decoder(16#86#)) OR
 					(reg_q303 AND symb_decoder(16#c9#)) OR
 					(reg_q303 AND symb_decoder(16#22#)) OR
 					(reg_q303 AND symb_decoder(16#2d#)) OR
 					(reg_q303 AND symb_decoder(16#b9#)) OR
 					(reg_q303 AND symb_decoder(16#cc#)) OR
 					(reg_q303 AND symb_decoder(16#17#)) OR
 					(reg_q303 AND symb_decoder(16#93#)) OR
 					(reg_q303 AND symb_decoder(16#d1#)) OR
 					(reg_q303 AND symb_decoder(16#5a#)) OR
 					(reg_q303 AND symb_decoder(16#2a#)) OR
 					(reg_q303 AND symb_decoder(16#77#)) OR
 					(reg_q303 AND symb_decoder(16#fa#)) OR
 					(reg_q303 AND symb_decoder(16#5b#)) OR
 					(reg_q303 AND symb_decoder(16#e5#)) OR
 					(reg_q303 AND symb_decoder(16#f3#)) OR
 					(reg_q303 AND symb_decoder(16#ce#)) OR
 					(reg_q303 AND symb_decoder(16#bf#)) OR
 					(reg_q303 AND symb_decoder(16#8b#)) OR
 					(reg_q303 AND symb_decoder(16#d6#)) OR
 					(reg_q303 AND symb_decoder(16#d7#)) OR
 					(reg_q303 AND symb_decoder(16#9e#)) OR
 					(reg_q303 AND symb_decoder(16#c4#)) OR
 					(reg_q303 AND symb_decoder(16#cf#)) OR
 					(reg_q303 AND symb_decoder(16#26#)) OR
 					(reg_q303 AND symb_decoder(16#2f#)) OR
 					(reg_q303 AND symb_decoder(16#0c#)) OR
 					(reg_q303 AND symb_decoder(16#32#)) OR
 					(reg_q303 AND symb_decoder(16#97#)) OR
 					(reg_q303 AND symb_decoder(16#95#)) OR
 					(reg_q303 AND symb_decoder(16#84#)) OR
 					(reg_q303 AND symb_decoder(16#cd#)) OR
 					(reg_q303 AND symb_decoder(16#54#)) OR
 					(reg_q303 AND symb_decoder(16#10#)) OR
 					(reg_q303 AND symb_decoder(16#6e#)) OR
 					(reg_q303 AND symb_decoder(16#1d#)) OR
 					(reg_q303 AND symb_decoder(16#04#)) OR
 					(reg_q303 AND symb_decoder(16#48#)) OR
 					(reg_q303 AND symb_decoder(16#5e#)) OR
 					(reg_q303 AND symb_decoder(16#e0#)) OR
 					(reg_q303 AND symb_decoder(16#9f#)) OR
 					(reg_q303 AND symb_decoder(16#fc#)) OR
 					(reg_q303 AND symb_decoder(16#4b#)) OR
 					(reg_q303 AND symb_decoder(16#df#)) OR
 					(reg_q303 AND symb_decoder(16#a3#)) OR
 					(reg_q303 AND symb_decoder(16#0a#)) OR
 					(reg_q303 AND symb_decoder(16#1e#)) OR
 					(reg_q303 AND symb_decoder(16#5f#)) OR
 					(reg_q303 AND symb_decoder(16#91#)) OR
 					(reg_q303 AND symb_decoder(16#60#)) OR
 					(reg_q303 AND symb_decoder(16#57#)) OR
 					(reg_q303 AND symb_decoder(16#40#)) OR
 					(reg_q303 AND symb_decoder(16#d4#)) OR
 					(reg_q303 AND symb_decoder(16#9d#)) OR
 					(reg_q303 AND symb_decoder(16#99#)) OR
 					(reg_q303 AND symb_decoder(16#8d#)) OR
 					(reg_q303 AND symb_decoder(16#8c#)) OR
 					(reg_q303 AND symb_decoder(16#c1#)) OR
 					(reg_q303 AND symb_decoder(16#28#)) OR
 					(reg_q303 AND symb_decoder(16#f8#)) OR
 					(reg_q303 AND symb_decoder(16#dd#)) OR
 					(reg_q303 AND symb_decoder(16#0e#)) OR
 					(reg_q303 AND symb_decoder(16#ee#)) OR
 					(reg_q303 AND symb_decoder(16#fb#)) OR
 					(reg_q303 AND symb_decoder(16#64#)) OR
 					(reg_q303 AND symb_decoder(16#e2#)) OR
 					(reg_q303 AND symb_decoder(16#92#)) OR
 					(reg_q303 AND symb_decoder(16#56#)) OR
 					(reg_q303 AND symb_decoder(16#cb#)) OR
 					(reg_q303 AND symb_decoder(16#d0#)) OR
 					(reg_q303 AND symb_decoder(16#9c#)) OR
 					(reg_q303 AND symb_decoder(16#46#)) OR
 					(reg_q303 AND symb_decoder(16#20#)) OR
 					(reg_q303 AND symb_decoder(16#30#)) OR
 					(reg_q303 AND symb_decoder(16#ac#)) OR
 					(reg_q303 AND symb_decoder(16#2b#)) OR
 					(reg_q303 AND symb_decoder(16#7e#)) OR
 					(reg_q303 AND symb_decoder(16#0f#)) OR
 					(reg_q303 AND symb_decoder(16#34#)) OR
 					(reg_q303 AND symb_decoder(16#ec#)) OR
 					(reg_q303 AND symb_decoder(16#ef#)) OR
 					(reg_q303 AND symb_decoder(16#db#)) OR
 					(reg_q303 AND symb_decoder(16#bc#)) OR
 					(reg_q303 AND symb_decoder(16#21#)) OR
 					(reg_q303 AND symb_decoder(16#e6#)) OR
 					(reg_q303 AND symb_decoder(16#2c#)) OR
 					(reg_q303 AND symb_decoder(16#61#)) OR
 					(reg_q303 AND symb_decoder(16#f7#)) OR
 					(reg_q303 AND symb_decoder(16#b4#)) OR
 					(reg_q303 AND symb_decoder(16#ff#)) OR
 					(reg_q303 AND symb_decoder(16#12#)) OR
 					(reg_q303 AND symb_decoder(16#79#)) OR
 					(reg_q303 AND symb_decoder(16#23#)) OR
 					(reg_q303 AND symb_decoder(16#74#)) OR
 					(reg_q303 AND symb_decoder(16#a8#)) OR
 					(reg_q303 AND symb_decoder(16#aa#)) OR
 					(reg_q303 AND symb_decoder(16#b6#)) OR
 					(reg_q303 AND symb_decoder(16#83#)) OR
 					(reg_q303 AND symb_decoder(16#7b#)) OR
 					(reg_q303 AND symb_decoder(16#06#)) OR
 					(reg_q303 AND symb_decoder(16#fe#)) OR
 					(reg_q303 AND symb_decoder(16#3f#)) OR
 					(reg_q303 AND symb_decoder(16#bd#)) OR
 					(reg_q303 AND symb_decoder(16#0b#)) OR
 					(reg_q303 AND symb_decoder(16#dc#)) OR
 					(reg_q303 AND symb_decoder(16#f4#)) OR
 					(reg_q303 AND symb_decoder(16#76#)) OR
 					(reg_q303 AND symb_decoder(16#02#)) OR
 					(reg_q303 AND symb_decoder(16#a4#)) OR
 					(reg_q303 AND symb_decoder(16#72#)) OR
 					(reg_q303 AND symb_decoder(16#b0#)) OR
 					(reg_q303 AND symb_decoder(16#6a#)) OR
 					(reg_q303 AND symb_decoder(16#67#)) OR
 					(reg_q303 AND symb_decoder(16#f0#)) OR
 					(reg_q303 AND symb_decoder(16#8f#)) OR
 					(reg_q303 AND symb_decoder(16#8e#)) OR
 					(reg_q303 AND symb_decoder(16#bb#)) OR
 					(reg_q303 AND symb_decoder(16#41#)) OR
 					(reg_q303 AND symb_decoder(16#ca#)) OR
 					(reg_q303 AND symb_decoder(16#6d#)) OR
 					(reg_q303 AND symb_decoder(16#f6#)) OR
 					(reg_q303 AND symb_decoder(16#29#)) OR
 					(reg_q303 AND symb_decoder(16#ed#)) OR
 					(reg_q303 AND symb_decoder(16#a2#)) OR
 					(reg_q303 AND symb_decoder(16#88#)) OR
 					(reg_q303 AND symb_decoder(16#25#)) OR
 					(reg_q303 AND symb_decoder(16#3e#)) OR
 					(reg_q303 AND symb_decoder(16#45#)) OR
 					(reg_q303 AND symb_decoder(16#c3#)) OR
 					(reg_q303 AND symb_decoder(16#c6#)) OR
 					(reg_q303 AND symb_decoder(16#ae#)) OR
 					(reg_q303 AND symb_decoder(16#5c#)) OR
 					(reg_q303 AND symb_decoder(16#18#)) OR
 					(reg_q303 AND symb_decoder(16#36#)) OR
 					(reg_q303 AND symb_decoder(16#f1#)) OR
 					(reg_q303 AND symb_decoder(16#85#)) OR
 					(reg_q303 AND symb_decoder(16#66#)) OR
 					(reg_q303 AND symb_decoder(16#4c#)) OR
 					(reg_q303 AND symb_decoder(16#31#)) OR
 					(reg_q303 AND symb_decoder(16#4e#)) OR
 					(reg_q303 AND symb_decoder(16#80#)) OR
 					(reg_q303 AND symb_decoder(16#e8#)) OR
 					(reg_q303 AND symb_decoder(16#6b#)) OR
 					(reg_q303 AND symb_decoder(16#ba#)) OR
 					(reg_q303 AND symb_decoder(16#b2#)) OR
 					(reg_q303 AND symb_decoder(16#1a#)) OR
 					(reg_q303 AND symb_decoder(16#a5#)) OR
 					(reg_q303 AND symb_decoder(16#14#)) OR
 					(reg_q303 AND symb_decoder(16#d2#)) OR
 					(reg_q303 AND symb_decoder(16#e3#)) OR
 					(reg_q303 AND symb_decoder(16#11#)) OR
 					(reg_q303 AND symb_decoder(16#c5#)) OR
 					(reg_q303 AND symb_decoder(16#8a#)) OR
 					(reg_q303 AND symb_decoder(16#c2#)) OR
 					(reg_q303 AND symb_decoder(16#a7#)) OR
 					(reg_q303 AND symb_decoder(16#6c#)) OR
 					(reg_q303 AND symb_decoder(16#53#)) OR
 					(reg_q303 AND symb_decoder(16#4d#)) OR
 					(reg_q303 AND symb_decoder(16#38#)) OR
 					(reg_q303 AND symb_decoder(16#6f#)) OR
 					(reg_q303 AND symb_decoder(16#b7#)) OR
 					(reg_q303 AND symb_decoder(16#b1#)) OR
 					(reg_q303 AND symb_decoder(16#f5#)) OR
 					(reg_q303 AND symb_decoder(16#ad#)) OR
 					(reg_q303 AND symb_decoder(16#3d#)) OR
 					(reg_q303 AND symb_decoder(16#e1#)) OR
 					(reg_q303 AND symb_decoder(16#44#)) OR
 					(reg_q303 AND symb_decoder(16#58#)) OR
 					(reg_q303 AND symb_decoder(16#0d#)) OR
 					(reg_q303 AND symb_decoder(16#13#)) OR
 					(reg_q303 AND symb_decoder(16#3b#)) OR
 					(reg_q303 AND symb_decoder(16#af#)) OR
 					(reg_q303 AND symb_decoder(16#2e#)) OR
 					(reg_q303 AND symb_decoder(16#a6#)) OR
 					(reg_q303 AND symb_decoder(16#62#)) OR
 					(reg_q303 AND symb_decoder(16#15#)) OR
 					(reg_q303 AND symb_decoder(16#87#)) OR
 					(reg_q303 AND symb_decoder(16#e9#)) OR
 					(reg_q303 AND symb_decoder(16#73#)) OR
 					(reg_q303 AND symb_decoder(16#ab#)) OR
 					(reg_q303 AND symb_decoder(16#19#)) OR
 					(reg_q303 AND symb_decoder(16#ea#)) OR
 					(reg_q303 AND symb_decoder(16#c8#)) OR
 					(reg_q303 AND symb_decoder(16#e7#)) OR
 					(reg_q303 AND symb_decoder(16#da#)) OR
 					(reg_q303 AND symb_decoder(16#a0#)) OR
 					(reg_q303 AND symb_decoder(16#68#)) OR
 					(reg_q303 AND symb_decoder(16#1c#)) OR
 					(reg_q303 AND symb_decoder(16#c0#)) OR
 					(reg_q303 AND symb_decoder(16#05#)) OR
 					(reg_q303 AND symb_decoder(16#39#)) OR
 					(reg_q303 AND symb_decoder(16#35#)) OR
 					(reg_q303 AND symb_decoder(16#01#)) OR
 					(reg_q303 AND symb_decoder(16#98#)) OR
 					(reg_q303 AND symb_decoder(16#a9#)) OR
 					(reg_q303 AND symb_decoder(16#08#)) OR
 					(reg_q303 AND symb_decoder(16#b5#)) OR
 					(reg_q303 AND symb_decoder(16#d5#)) OR
 					(reg_q303 AND symb_decoder(16#63#)) OR
 					(reg_q303 AND symb_decoder(16#47#)) OR
 					(reg_q303 AND symb_decoder(16#49#)) OR
 					(reg_q303 AND symb_decoder(16#51#)) OR
 					(reg_q303 AND symb_decoder(16#75#)) OR
 					(reg_q303 AND symb_decoder(16#70#)) OR
 					(reg_q303 AND symb_decoder(16#59#)) OR
 					(reg_q303 AND symb_decoder(16#4f#)) OR
 					(reg_q303 AND symb_decoder(16#69#)) OR
 					(reg_q303 AND symb_decoder(16#00#)) OR
 					(reg_q303 AND symb_decoder(16#fd#)) OR
 					(reg_q303 AND symb_decoder(16#65#)) OR
 					(reg_q303 AND symb_decoder(16#9b#)) OR
 					(reg_q303 AND symb_decoder(16#d3#)) OR
 					(reg_q303 AND symb_decoder(16#81#));
reg_q303_init <= '0' ;
	p_reg_q303: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q303 <= reg_q303_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q303 <= reg_q303_init;
        else
          reg_q303 <= reg_q303_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q665_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q665 AND symb_decoder(16#bf#)) OR
 					(reg_q665 AND symb_decoder(16#70#)) OR
 					(reg_q665 AND symb_decoder(16#3f#)) OR
 					(reg_q665 AND symb_decoder(16#4a#)) OR
 					(reg_q665 AND symb_decoder(16#8d#)) OR
 					(reg_q665 AND symb_decoder(16#a7#)) OR
 					(reg_q665 AND symb_decoder(16#25#)) OR
 					(reg_q665 AND symb_decoder(16#75#)) OR
 					(reg_q665 AND symb_decoder(16#1a#)) OR
 					(reg_q665 AND symb_decoder(16#9d#)) OR
 					(reg_q665 AND symb_decoder(16#a6#)) OR
 					(reg_q665 AND symb_decoder(16#6d#)) OR
 					(reg_q665 AND symb_decoder(16#13#)) OR
 					(reg_q665 AND symb_decoder(16#20#)) OR
 					(reg_q665 AND symb_decoder(16#23#)) OR
 					(reg_q665 AND symb_decoder(16#0d#)) OR
 					(reg_q665 AND symb_decoder(16#28#)) OR
 					(reg_q665 AND symb_decoder(16#94#)) OR
 					(reg_q665 AND symb_decoder(16#6f#)) OR
 					(reg_q665 AND symb_decoder(16#31#)) OR
 					(reg_q665 AND symb_decoder(16#fe#)) OR
 					(reg_q665 AND symb_decoder(16#77#)) OR
 					(reg_q665 AND symb_decoder(16#73#)) OR
 					(reg_q665 AND symb_decoder(16#43#)) OR
 					(reg_q665 AND symb_decoder(16#ca#)) OR
 					(reg_q665 AND symb_decoder(16#c5#)) OR
 					(reg_q665 AND symb_decoder(16#12#)) OR
 					(reg_q665 AND symb_decoder(16#ab#)) OR
 					(reg_q665 AND symb_decoder(16#62#)) OR
 					(reg_q665 AND symb_decoder(16#69#)) OR
 					(reg_q665 AND symb_decoder(16#7d#)) OR
 					(reg_q665 AND symb_decoder(16#c0#)) OR
 					(reg_q665 AND symb_decoder(16#ee#)) OR
 					(reg_q665 AND symb_decoder(16#b2#)) OR
 					(reg_q665 AND symb_decoder(16#ff#)) OR
 					(reg_q665 AND symb_decoder(16#a0#)) OR
 					(reg_q665 AND symb_decoder(16#bc#)) OR
 					(reg_q665 AND symb_decoder(16#46#)) OR
 					(reg_q665 AND symb_decoder(16#6c#)) OR
 					(reg_q665 AND symb_decoder(16#9b#)) OR
 					(reg_q665 AND symb_decoder(16#51#)) OR
 					(reg_q665 AND symb_decoder(16#68#)) OR
 					(reg_q665 AND symb_decoder(16#a4#)) OR
 					(reg_q665 AND symb_decoder(16#99#)) OR
 					(reg_q665 AND symb_decoder(16#2d#)) OR
 					(reg_q665 AND symb_decoder(16#56#)) OR
 					(reg_q665 AND symb_decoder(16#be#)) OR
 					(reg_q665 AND symb_decoder(16#c3#)) OR
 					(reg_q665 AND symb_decoder(16#b4#)) OR
 					(reg_q665 AND symb_decoder(16#aa#)) OR
 					(reg_q665 AND symb_decoder(16#1c#)) OR
 					(reg_q665 AND symb_decoder(16#4c#)) OR
 					(reg_q665 AND symb_decoder(16#11#)) OR
 					(reg_q665 AND symb_decoder(16#5f#)) OR
 					(reg_q665 AND symb_decoder(16#6b#)) OR
 					(reg_q665 AND symb_decoder(16#82#)) OR
 					(reg_q665 AND symb_decoder(16#24#)) OR
 					(reg_q665 AND symb_decoder(16#93#)) OR
 					(reg_q665 AND symb_decoder(16#e6#)) OR
 					(reg_q665 AND symb_decoder(16#a5#)) OR
 					(reg_q665 AND symb_decoder(16#e1#)) OR
 					(reg_q665 AND symb_decoder(16#1d#)) OR
 					(reg_q665 AND symb_decoder(16#5c#)) OR
 					(reg_q665 AND symb_decoder(16#a2#)) OR
 					(reg_q665 AND symb_decoder(16#40#)) OR
 					(reg_q665 AND symb_decoder(16#bd#)) OR
 					(reg_q665 AND symb_decoder(16#7b#)) OR
 					(reg_q665 AND symb_decoder(16#41#)) OR
 					(reg_q665 AND symb_decoder(16#66#)) OR
 					(reg_q665 AND symb_decoder(16#5e#)) OR
 					(reg_q665 AND symb_decoder(16#9c#)) OR
 					(reg_q665 AND symb_decoder(16#3e#)) OR
 					(reg_q665 AND symb_decoder(16#64#)) OR
 					(reg_q665 AND symb_decoder(16#5b#)) OR
 					(reg_q665 AND symb_decoder(16#90#)) OR
 					(reg_q665 AND symb_decoder(16#7f#)) OR
 					(reg_q665 AND symb_decoder(16#fb#)) OR
 					(reg_q665 AND symb_decoder(16#02#)) OR
 					(reg_q665 AND symb_decoder(16#5d#)) OR
 					(reg_q665 AND symb_decoder(16#39#)) OR
 					(reg_q665 AND symb_decoder(16#48#)) OR
 					(reg_q665 AND symb_decoder(16#f5#)) OR
 					(reg_q665 AND symb_decoder(16#83#)) OR
 					(reg_q665 AND symb_decoder(16#86#)) OR
 					(reg_q665 AND symb_decoder(16#03#)) OR
 					(reg_q665 AND symb_decoder(16#57#)) OR
 					(reg_q665 AND symb_decoder(16#72#)) OR
 					(reg_q665 AND symb_decoder(16#61#)) OR
 					(reg_q665 AND symb_decoder(16#63#)) OR
 					(reg_q665 AND symb_decoder(16#fd#)) OR
 					(reg_q665 AND symb_decoder(16#ad#)) OR
 					(reg_q665 AND symb_decoder(16#dc#)) OR
 					(reg_q665 AND symb_decoder(16#cc#)) OR
 					(reg_q665 AND symb_decoder(16#8a#)) OR
 					(reg_q665 AND symb_decoder(16#c4#)) OR
 					(reg_q665 AND symb_decoder(16#71#)) OR
 					(reg_q665 AND symb_decoder(16#1f#)) OR
 					(reg_q665 AND symb_decoder(16#45#)) OR
 					(reg_q665 AND symb_decoder(16#5a#)) OR
 					(reg_q665 AND symb_decoder(16#27#)) OR
 					(reg_q665 AND symb_decoder(16#49#)) OR
 					(reg_q665 AND symb_decoder(16#17#)) OR
 					(reg_q665 AND symb_decoder(16#0a#)) OR
 					(reg_q665 AND symb_decoder(16#c1#)) OR
 					(reg_q665 AND symb_decoder(16#9e#)) OR
 					(reg_q665 AND symb_decoder(16#55#)) OR
 					(reg_q665 AND symb_decoder(16#15#)) OR
 					(reg_q665 AND symb_decoder(16#00#)) OR
 					(reg_q665 AND symb_decoder(16#d9#)) OR
 					(reg_q665 AND symb_decoder(16#d3#)) OR
 					(reg_q665 AND symb_decoder(16#b9#)) OR
 					(reg_q665 AND symb_decoder(16#ba#)) OR
 					(reg_q665 AND symb_decoder(16#78#)) OR
 					(reg_q665 AND symb_decoder(16#d1#)) OR
 					(reg_q665 AND symb_decoder(16#4d#)) OR
 					(reg_q665 AND symb_decoder(16#67#)) OR
 					(reg_q665 AND symb_decoder(16#22#)) OR
 					(reg_q665 AND symb_decoder(16#2b#)) OR
 					(reg_q665 AND symb_decoder(16#87#)) OR
 					(reg_q665 AND symb_decoder(16#36#)) OR
 					(reg_q665 AND symb_decoder(16#bb#)) OR
 					(reg_q665 AND symb_decoder(16#de#)) OR
 					(reg_q665 AND symb_decoder(16#f9#)) OR
 					(reg_q665 AND symb_decoder(16#e9#)) OR
 					(reg_q665 AND symb_decoder(16#81#)) OR
 					(reg_q665 AND symb_decoder(16#98#)) OR
 					(reg_q665 AND symb_decoder(16#c8#)) OR
 					(reg_q665 AND symb_decoder(16#b5#)) OR
 					(reg_q665 AND symb_decoder(16#c6#)) OR
 					(reg_q665 AND symb_decoder(16#88#)) OR
 					(reg_q665 AND symb_decoder(16#f3#)) OR
 					(reg_q665 AND symb_decoder(16#7c#)) OR
 					(reg_q665 AND symb_decoder(16#ae#)) OR
 					(reg_q665 AND symb_decoder(16#1b#)) OR
 					(reg_q665 AND symb_decoder(16#eb#)) OR
 					(reg_q665 AND symb_decoder(16#89#)) OR
 					(reg_q665 AND symb_decoder(16#d2#)) OR
 					(reg_q665 AND symb_decoder(16#7e#)) OR
 					(reg_q665 AND symb_decoder(16#18#)) OR
 					(reg_q665 AND symb_decoder(16#8e#)) OR
 					(reg_q665 AND symb_decoder(16#8f#)) OR
 					(reg_q665 AND symb_decoder(16#44#)) OR
 					(reg_q665 AND symb_decoder(16#07#)) OR
 					(reg_q665 AND symb_decoder(16#cf#)) OR
 					(reg_q665 AND symb_decoder(16#74#)) OR
 					(reg_q665 AND symb_decoder(16#37#)) OR
 					(reg_q665 AND symb_decoder(16#ec#)) OR
 					(reg_q665 AND symb_decoder(16#09#)) OR
 					(reg_q665 AND symb_decoder(16#4e#)) OR
 					(reg_q665 AND symb_decoder(16#96#)) OR
 					(reg_q665 AND symb_decoder(16#50#)) OR
 					(reg_q665 AND symb_decoder(16#58#)) OR
 					(reg_q665 AND symb_decoder(16#a9#)) OR
 					(reg_q665 AND symb_decoder(16#df#)) OR
 					(reg_q665 AND symb_decoder(16#f1#)) OR
 					(reg_q665 AND symb_decoder(16#2a#)) OR
 					(reg_q665 AND symb_decoder(16#3c#)) OR
 					(reg_q665 AND symb_decoder(16#ed#)) OR
 					(reg_q665 AND symb_decoder(16#f7#)) OR
 					(reg_q665 AND symb_decoder(16#e4#)) OR
 					(reg_q665 AND symb_decoder(16#6a#)) OR
 					(reg_q665 AND symb_decoder(16#7a#)) OR
 					(reg_q665 AND symb_decoder(16#b6#)) OR
 					(reg_q665 AND symb_decoder(16#c7#)) OR
 					(reg_q665 AND symb_decoder(16#3d#)) OR
 					(reg_q665 AND symb_decoder(16#db#)) OR
 					(reg_q665 AND symb_decoder(16#16#)) OR
 					(reg_q665 AND symb_decoder(16#59#)) OR
 					(reg_q665 AND symb_decoder(16#8b#)) OR
 					(reg_q665 AND symb_decoder(16#dd#)) OR
 					(reg_q665 AND symb_decoder(16#d0#)) OR
 					(reg_q665 AND symb_decoder(16#65#)) OR
 					(reg_q665 AND symb_decoder(16#38#)) OR
 					(reg_q665 AND symb_decoder(16#60#)) OR
 					(reg_q665 AND symb_decoder(16#b0#)) OR
 					(reg_q665 AND symb_decoder(16#b8#)) OR
 					(reg_q665 AND symb_decoder(16#01#)) OR
 					(reg_q665 AND symb_decoder(16#04#)) OR
 					(reg_q665 AND symb_decoder(16#0c#)) OR
 					(reg_q665 AND symb_decoder(16#0e#)) OR
 					(reg_q665 AND symb_decoder(16#10#)) OR
 					(reg_q665 AND symb_decoder(16#c9#)) OR
 					(reg_q665 AND symb_decoder(16#f8#)) OR
 					(reg_q665 AND symb_decoder(16#30#)) OR
 					(reg_q665 AND symb_decoder(16#32#)) OR
 					(reg_q665 AND symb_decoder(16#53#)) OR
 					(reg_q665 AND symb_decoder(16#9a#)) OR
 					(reg_q665 AND symb_decoder(16#92#)) OR
 					(reg_q665 AND symb_decoder(16#1e#)) OR
 					(reg_q665 AND symb_decoder(16#3a#)) OR
 					(reg_q665 AND symb_decoder(16#35#)) OR
 					(reg_q665 AND symb_decoder(16#05#)) OR
 					(reg_q665 AND symb_decoder(16#8c#)) OR
 					(reg_q665 AND symb_decoder(16#2f#)) OR
 					(reg_q665 AND symb_decoder(16#e0#)) OR
 					(reg_q665 AND symb_decoder(16#91#)) OR
 					(reg_q665 AND symb_decoder(16#42#)) OR
 					(reg_q665 AND symb_decoder(16#97#)) OR
 					(reg_q665 AND symb_decoder(16#80#)) OR
 					(reg_q665 AND symb_decoder(16#ac#)) OR
 					(reg_q665 AND symb_decoder(16#52#)) OR
 					(reg_q665 AND symb_decoder(16#d4#)) OR
 					(reg_q665 AND symb_decoder(16#ce#)) OR
 					(reg_q665 AND symb_decoder(16#b1#)) OR
 					(reg_q665 AND symb_decoder(16#fa#)) OR
 					(reg_q665 AND symb_decoder(16#34#)) OR
 					(reg_q665 AND symb_decoder(16#e2#)) OR
 					(reg_q665 AND symb_decoder(16#e7#)) OR
 					(reg_q665 AND symb_decoder(16#a3#)) OR
 					(reg_q665 AND symb_decoder(16#95#)) OR
 					(reg_q665 AND symb_decoder(16#a1#)) OR
 					(reg_q665 AND symb_decoder(16#3b#)) OR
 					(reg_q665 AND symb_decoder(16#f6#)) OR
 					(reg_q665 AND symb_decoder(16#84#)) OR
 					(reg_q665 AND symb_decoder(16#d5#)) OR
 					(reg_q665 AND symb_decoder(16#79#)) OR
 					(reg_q665 AND symb_decoder(16#cb#)) OR
 					(reg_q665 AND symb_decoder(16#21#)) OR
 					(reg_q665 AND symb_decoder(16#0f#)) OR
 					(reg_q665 AND symb_decoder(16#2c#)) OR
 					(reg_q665 AND symb_decoder(16#e3#)) OR
 					(reg_q665 AND symb_decoder(16#ea#)) OR
 					(reg_q665 AND symb_decoder(16#a8#)) OR
 					(reg_q665 AND symb_decoder(16#85#)) OR
 					(reg_q665 AND symb_decoder(16#4b#)) OR
 					(reg_q665 AND symb_decoder(16#d6#)) OR
 					(reg_q665 AND symb_decoder(16#d8#)) OR
 					(reg_q665 AND symb_decoder(16#9f#)) OR
 					(reg_q665 AND symb_decoder(16#08#)) OR
 					(reg_q665 AND symb_decoder(16#47#)) OR
 					(reg_q665 AND symb_decoder(16#0b#)) OR
 					(reg_q665 AND symb_decoder(16#ef#)) OR
 					(reg_q665 AND symb_decoder(16#76#)) OR
 					(reg_q665 AND symb_decoder(16#b7#)) OR
 					(reg_q665 AND symb_decoder(16#06#)) OR
 					(reg_q665 AND symb_decoder(16#14#)) OR
 					(reg_q665 AND symb_decoder(16#6e#)) OR
 					(reg_q665 AND symb_decoder(16#26#)) OR
 					(reg_q665 AND symb_decoder(16#f0#)) OR
 					(reg_q665 AND symb_decoder(16#19#)) OR
 					(reg_q665 AND symb_decoder(16#b3#)) OR
 					(reg_q665 AND symb_decoder(16#4f#)) OR
 					(reg_q665 AND symb_decoder(16#da#)) OR
 					(reg_q665 AND symb_decoder(16#af#)) OR
 					(reg_q665 AND symb_decoder(16#c2#)) OR
 					(reg_q665 AND symb_decoder(16#f4#)) OR
 					(reg_q665 AND symb_decoder(16#29#)) OR
 					(reg_q665 AND symb_decoder(16#fc#)) OR
 					(reg_q665 AND symb_decoder(16#33#)) OR
 					(reg_q665 AND symb_decoder(16#54#)) OR
 					(reg_q665 AND symb_decoder(16#cd#)) OR
 					(reg_q665 AND symb_decoder(16#2e#)) OR
 					(reg_q665 AND symb_decoder(16#e8#)) OR
 					(reg_q665 AND symb_decoder(16#d7#)) OR
 					(reg_q665 AND symb_decoder(16#f2#)) OR
 					(reg_q665 AND symb_decoder(16#e5#));
reg_q665_init <= '0' ;
	p_reg_q665: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q665 <= reg_q665_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q665 <= reg_q665_init;
        else
          reg_q665 <= reg_q665_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q703_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q703 AND symb_decoder(16#bb#)) OR
 					(reg_q703 AND symb_decoder(16#a7#)) OR
 					(reg_q703 AND symb_decoder(16#b1#)) OR
 					(reg_q703 AND symb_decoder(16#77#)) OR
 					(reg_q703 AND symb_decoder(16#2d#)) OR
 					(reg_q703 AND symb_decoder(16#64#)) OR
 					(reg_q703 AND symb_decoder(16#3f#)) OR
 					(reg_q703 AND symb_decoder(16#19#)) OR
 					(reg_q703 AND symb_decoder(16#cc#)) OR
 					(reg_q703 AND symb_decoder(16#dc#)) OR
 					(reg_q703 AND symb_decoder(16#c3#)) OR
 					(reg_q703 AND symb_decoder(16#f1#)) OR
 					(reg_q703 AND symb_decoder(16#ab#)) OR
 					(reg_q703 AND symb_decoder(16#a0#)) OR
 					(reg_q703 AND symb_decoder(16#5d#)) OR
 					(reg_q703 AND symb_decoder(16#2c#)) OR
 					(reg_q703 AND symb_decoder(16#92#)) OR
 					(reg_q703 AND symb_decoder(16#63#)) OR
 					(reg_q703 AND symb_decoder(16#52#)) OR
 					(reg_q703 AND symb_decoder(16#17#)) OR
 					(reg_q703 AND symb_decoder(16#fb#)) OR
 					(reg_q703 AND symb_decoder(16#30#)) OR
 					(reg_q703 AND symb_decoder(16#29#)) OR
 					(reg_q703 AND symb_decoder(16#31#)) OR
 					(reg_q703 AND symb_decoder(16#a3#)) OR
 					(reg_q703 AND symb_decoder(16#d5#)) OR
 					(reg_q703 AND symb_decoder(16#58#)) OR
 					(reg_q703 AND symb_decoder(16#98#)) OR
 					(reg_q703 AND symb_decoder(16#2e#)) OR
 					(reg_q703 AND symb_decoder(16#09#)) OR
 					(reg_q703 AND symb_decoder(16#fe#)) OR
 					(reg_q703 AND symb_decoder(16#8e#)) OR
 					(reg_q703 AND symb_decoder(16#0d#)) OR
 					(reg_q703 AND symb_decoder(16#1e#)) OR
 					(reg_q703 AND symb_decoder(16#83#)) OR
 					(reg_q703 AND symb_decoder(16#8c#)) OR
 					(reg_q703 AND symb_decoder(16#a5#)) OR
 					(reg_q703 AND symb_decoder(16#37#)) OR
 					(reg_q703 AND symb_decoder(16#78#)) OR
 					(reg_q703 AND symb_decoder(16#73#)) OR
 					(reg_q703 AND symb_decoder(16#20#)) OR
 					(reg_q703 AND symb_decoder(16#f7#)) OR
 					(reg_q703 AND symb_decoder(16#b5#)) OR
 					(reg_q703 AND symb_decoder(16#8a#)) OR
 					(reg_q703 AND symb_decoder(16#23#)) OR
 					(reg_q703 AND symb_decoder(16#99#)) OR
 					(reg_q703 AND symb_decoder(16#02#)) OR
 					(reg_q703 AND symb_decoder(16#96#)) OR
 					(reg_q703 AND symb_decoder(16#e7#)) OR
 					(reg_q703 AND symb_decoder(16#f2#)) OR
 					(reg_q703 AND symb_decoder(16#f9#)) OR
 					(reg_q703 AND symb_decoder(16#f5#)) OR
 					(reg_q703 AND symb_decoder(16#8f#)) OR
 					(reg_q703 AND symb_decoder(16#be#)) OR
 					(reg_q703 AND symb_decoder(16#ad#)) OR
 					(reg_q703 AND symb_decoder(16#8b#)) OR
 					(reg_q703 AND symb_decoder(16#56#)) OR
 					(reg_q703 AND symb_decoder(16#9f#)) OR
 					(reg_q703 AND symb_decoder(16#95#)) OR
 					(reg_q703 AND symb_decoder(16#df#)) OR
 					(reg_q703 AND symb_decoder(16#a6#)) OR
 					(reg_q703 AND symb_decoder(16#da#)) OR
 					(reg_q703 AND symb_decoder(16#e2#)) OR
 					(reg_q703 AND symb_decoder(16#ed#)) OR
 					(reg_q703 AND symb_decoder(16#32#)) OR
 					(reg_q703 AND symb_decoder(16#12#)) OR
 					(reg_q703 AND symb_decoder(16#4b#)) OR
 					(reg_q703 AND symb_decoder(16#c0#)) OR
 					(reg_q703 AND symb_decoder(16#2b#)) OR
 					(reg_q703 AND symb_decoder(16#2f#)) OR
 					(reg_q703 AND symb_decoder(16#e4#)) OR
 					(reg_q703 AND symb_decoder(16#d6#)) OR
 					(reg_q703 AND symb_decoder(16#06#)) OR
 					(reg_q703 AND symb_decoder(16#e3#)) OR
 					(reg_q703 AND symb_decoder(16#60#)) OR
 					(reg_q703 AND symb_decoder(16#4c#)) OR
 					(reg_q703 AND symb_decoder(16#24#)) OR
 					(reg_q703 AND symb_decoder(16#66#)) OR
 					(reg_q703 AND symb_decoder(16#57#)) OR
 					(reg_q703 AND symb_decoder(16#25#)) OR
 					(reg_q703 AND symb_decoder(16#ef#)) OR
 					(reg_q703 AND symb_decoder(16#cd#)) OR
 					(reg_q703 AND symb_decoder(16#54#)) OR
 					(reg_q703 AND symb_decoder(16#84#)) OR
 					(reg_q703 AND symb_decoder(16#b8#)) OR
 					(reg_q703 AND symb_decoder(16#4e#)) OR
 					(reg_q703 AND symb_decoder(16#d8#)) OR
 					(reg_q703 AND symb_decoder(16#fd#)) OR
 					(reg_q703 AND symb_decoder(16#0c#)) OR
 					(reg_q703 AND symb_decoder(16#ea#)) OR
 					(reg_q703 AND symb_decoder(16#0b#)) OR
 					(reg_q703 AND symb_decoder(16#07#)) OR
 					(reg_q703 AND symb_decoder(16#62#)) OR
 					(reg_q703 AND symb_decoder(16#70#)) OR
 					(reg_q703 AND symb_decoder(16#88#)) OR
 					(reg_q703 AND symb_decoder(16#72#)) OR
 					(reg_q703 AND symb_decoder(16#7b#)) OR
 					(reg_q703 AND symb_decoder(16#1d#)) OR
 					(reg_q703 AND symb_decoder(16#d4#)) OR
 					(reg_q703 AND symb_decoder(16#d3#)) OR
 					(reg_q703 AND symb_decoder(16#e1#)) OR
 					(reg_q703 AND symb_decoder(16#de#)) OR
 					(reg_q703 AND symb_decoder(16#fc#)) OR
 					(reg_q703 AND symb_decoder(16#6f#)) OR
 					(reg_q703 AND symb_decoder(16#c2#)) OR
 					(reg_q703 AND symb_decoder(16#5c#)) OR
 					(reg_q703 AND symb_decoder(16#50#)) OR
 					(reg_q703 AND symb_decoder(16#90#)) OR
 					(reg_q703 AND symb_decoder(16#dd#)) OR
 					(reg_q703 AND symb_decoder(16#9b#)) OR
 					(reg_q703 AND symb_decoder(16#28#)) OR
 					(reg_q703 AND symb_decoder(16#a8#)) OR
 					(reg_q703 AND symb_decoder(16#75#)) OR
 					(reg_q703 AND symb_decoder(16#53#)) OR
 					(reg_q703 AND symb_decoder(16#b0#)) OR
 					(reg_q703 AND symb_decoder(16#1a#)) OR
 					(reg_q703 AND symb_decoder(16#0a#)) OR
 					(reg_q703 AND symb_decoder(16#81#)) OR
 					(reg_q703 AND symb_decoder(16#c7#)) OR
 					(reg_q703 AND symb_decoder(16#89#)) OR
 					(reg_q703 AND symb_decoder(16#7a#)) OR
 					(reg_q703 AND symb_decoder(16#13#)) OR
 					(reg_q703 AND symb_decoder(16#87#)) OR
 					(reg_q703 AND symb_decoder(16#b6#)) OR
 					(reg_q703 AND symb_decoder(16#03#)) OR
 					(reg_q703 AND symb_decoder(16#67#)) OR
 					(reg_q703 AND symb_decoder(16#a9#)) OR
 					(reg_q703 AND symb_decoder(16#9d#)) OR
 					(reg_q703 AND symb_decoder(16#38#)) OR
 					(reg_q703 AND symb_decoder(16#00#)) OR
 					(reg_q703 AND symb_decoder(16#af#)) OR
 					(reg_q703 AND symb_decoder(16#bc#)) OR
 					(reg_q703 AND symb_decoder(16#cf#)) OR
 					(reg_q703 AND symb_decoder(16#71#)) OR
 					(reg_q703 AND symb_decoder(16#3d#)) OR
 					(reg_q703 AND symb_decoder(16#c4#)) OR
 					(reg_q703 AND symb_decoder(16#3b#)) OR
 					(reg_q703 AND symb_decoder(16#1b#)) OR
 					(reg_q703 AND symb_decoder(16#d0#)) OR
 					(reg_q703 AND symb_decoder(16#3a#)) OR
 					(reg_q703 AND symb_decoder(16#f4#)) OR
 					(reg_q703 AND symb_decoder(16#10#)) OR
 					(reg_q703 AND symb_decoder(16#ce#)) OR
 					(reg_q703 AND symb_decoder(16#35#)) OR
 					(reg_q703 AND symb_decoder(16#ee#)) OR
 					(reg_q703 AND symb_decoder(16#c8#)) OR
 					(reg_q703 AND symb_decoder(16#49#)) OR
 					(reg_q703 AND symb_decoder(16#bf#)) OR
 					(reg_q703 AND symb_decoder(16#9c#)) OR
 					(reg_q703 AND symb_decoder(16#91#)) OR
 					(reg_q703 AND symb_decoder(16#85#)) OR
 					(reg_q703 AND symb_decoder(16#ca#)) OR
 					(reg_q703 AND symb_decoder(16#d2#)) OR
 					(reg_q703 AND symb_decoder(16#4d#)) OR
 					(reg_q703 AND symb_decoder(16#0e#)) OR
 					(reg_q703 AND symb_decoder(16#65#)) OR
 					(reg_q703 AND symb_decoder(16#b3#)) OR
 					(reg_q703 AND symb_decoder(16#3e#)) OR
 					(reg_q703 AND symb_decoder(16#e5#)) OR
 					(reg_q703 AND symb_decoder(16#14#)) OR
 					(reg_q703 AND symb_decoder(16#bd#)) OR
 					(reg_q703 AND symb_decoder(16#ec#)) OR
 					(reg_q703 AND symb_decoder(16#34#)) OR
 					(reg_q703 AND symb_decoder(16#d1#)) OR
 					(reg_q703 AND symb_decoder(16#f6#)) OR
 					(reg_q703 AND symb_decoder(16#d9#)) OR
 					(reg_q703 AND symb_decoder(16#b4#)) OR
 					(reg_q703 AND symb_decoder(16#6a#)) OR
 					(reg_q703 AND symb_decoder(16#ac#)) OR
 					(reg_q703 AND symb_decoder(16#7c#)) OR
 					(reg_q703 AND symb_decoder(16#69#)) OR
 					(reg_q703 AND symb_decoder(16#e8#)) OR
 					(reg_q703 AND symb_decoder(16#e9#)) OR
 					(reg_q703 AND symb_decoder(16#6c#)) OR
 					(reg_q703 AND symb_decoder(16#7f#)) OR
 					(reg_q703 AND symb_decoder(16#42#)) OR
 					(reg_q703 AND symb_decoder(16#ae#)) OR
 					(reg_q703 AND symb_decoder(16#40#)) OR
 					(reg_q703 AND symb_decoder(16#1f#)) OR
 					(reg_q703 AND symb_decoder(16#94#)) OR
 					(reg_q703 AND symb_decoder(16#cb#)) OR
 					(reg_q703 AND symb_decoder(16#e6#)) OR
 					(reg_q703 AND symb_decoder(16#80#)) OR
 					(reg_q703 AND symb_decoder(16#7d#)) OR
 					(reg_q703 AND symb_decoder(16#f8#)) OR
 					(reg_q703 AND symb_decoder(16#16#)) OR
 					(reg_q703 AND symb_decoder(16#f3#)) OR
 					(reg_q703 AND symb_decoder(16#6e#)) OR
 					(reg_q703 AND symb_decoder(16#4f#)) OR
 					(reg_q703 AND symb_decoder(16#39#)) OR
 					(reg_q703 AND symb_decoder(16#97#)) OR
 					(reg_q703 AND symb_decoder(16#55#)) OR
 					(reg_q703 AND symb_decoder(16#9a#)) OR
 					(reg_q703 AND symb_decoder(16#21#)) OR
 					(reg_q703 AND symb_decoder(16#5a#)) OR
 					(reg_q703 AND symb_decoder(16#a2#)) OR
 					(reg_q703 AND symb_decoder(16#76#)) OR
 					(reg_q703 AND symb_decoder(16#f0#)) OR
 					(reg_q703 AND symb_decoder(16#33#)) OR
 					(reg_q703 AND symb_decoder(16#43#)) OR
 					(reg_q703 AND symb_decoder(16#18#)) OR
 					(reg_q703 AND symb_decoder(16#79#)) OR
 					(reg_q703 AND symb_decoder(16#5f#)) OR
 					(reg_q703 AND symb_decoder(16#48#)) OR
 					(reg_q703 AND symb_decoder(16#46#)) OR
 					(reg_q703 AND symb_decoder(16#44#)) OR
 					(reg_q703 AND symb_decoder(16#82#)) OR
 					(reg_q703 AND symb_decoder(16#61#)) OR
 					(reg_q703 AND symb_decoder(16#b7#)) OR
 					(reg_q703 AND symb_decoder(16#fa#)) OR
 					(reg_q703 AND symb_decoder(16#5b#)) OR
 					(reg_q703 AND symb_decoder(16#b9#)) OR
 					(reg_q703 AND symb_decoder(16#c1#)) OR
 					(reg_q703 AND symb_decoder(16#1c#)) OR
 					(reg_q703 AND symb_decoder(16#ba#)) OR
 					(reg_q703 AND symb_decoder(16#93#)) OR
 					(reg_q703 AND symb_decoder(16#01#)) OR
 					(reg_q703 AND symb_decoder(16#86#)) OR
 					(reg_q703 AND symb_decoder(16#11#)) OR
 					(reg_q703 AND symb_decoder(16#4a#)) OR
 					(reg_q703 AND symb_decoder(16#db#)) OR
 					(reg_q703 AND symb_decoder(16#ff#)) OR
 					(reg_q703 AND symb_decoder(16#eb#)) OR
 					(reg_q703 AND symb_decoder(16#26#)) OR
 					(reg_q703 AND symb_decoder(16#68#)) OR
 					(reg_q703 AND symb_decoder(16#45#)) OR
 					(reg_q703 AND symb_decoder(16#e0#)) OR
 					(reg_q703 AND symb_decoder(16#51#)) OR
 					(reg_q703 AND symb_decoder(16#c5#)) OR
 					(reg_q703 AND symb_decoder(16#c9#)) OR
 					(reg_q703 AND symb_decoder(16#47#)) OR
 					(reg_q703 AND symb_decoder(16#aa#)) OR
 					(reg_q703 AND symb_decoder(16#7e#)) OR
 					(reg_q703 AND symb_decoder(16#d7#)) OR
 					(reg_q703 AND symb_decoder(16#b2#)) OR
 					(reg_q703 AND symb_decoder(16#6d#)) OR
 					(reg_q703 AND symb_decoder(16#59#)) OR
 					(reg_q703 AND symb_decoder(16#0f#)) OR
 					(reg_q703 AND symb_decoder(16#41#)) OR
 					(reg_q703 AND symb_decoder(16#3c#)) OR
 					(reg_q703 AND symb_decoder(16#6b#)) OR
 					(reg_q703 AND symb_decoder(16#a4#)) OR
 					(reg_q703 AND symb_decoder(16#15#)) OR
 					(reg_q703 AND symb_decoder(16#8d#)) OR
 					(reg_q703 AND symb_decoder(16#36#)) OR
 					(reg_q703 AND symb_decoder(16#27#)) OR
 					(reg_q703 AND symb_decoder(16#a1#)) OR
 					(reg_q703 AND symb_decoder(16#2a#)) OR
 					(reg_q703 AND symb_decoder(16#74#)) OR
 					(reg_q703 AND symb_decoder(16#9e#)) OR
 					(reg_q703 AND symb_decoder(16#04#)) OR
 					(reg_q703 AND symb_decoder(16#5e#)) OR
 					(reg_q703 AND symb_decoder(16#05#)) OR
 					(reg_q703 AND symb_decoder(16#08#)) OR
 					(reg_q703 AND symb_decoder(16#22#)) OR
 					(reg_q703 AND symb_decoder(16#c6#));
reg_q703_init <= '0' ;
	p_reg_q703: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q703 <= reg_q703_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q703 <= reg_q703_init;
        else
          reg_q703 <= reg_q703_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q414_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q414 AND symb_decoder(16#f8#)) OR
 					(reg_q414 AND symb_decoder(16#8f#)) OR
 					(reg_q414 AND symb_decoder(16#8a#)) OR
 					(reg_q414 AND symb_decoder(16#fa#)) OR
 					(reg_q414 AND symb_decoder(16#2c#)) OR
 					(reg_q414 AND symb_decoder(16#f1#)) OR
 					(reg_q414 AND symb_decoder(16#3a#)) OR
 					(reg_q414 AND symb_decoder(16#79#)) OR
 					(reg_q414 AND symb_decoder(16#b3#)) OR
 					(reg_q414 AND symb_decoder(16#cf#)) OR
 					(reg_q414 AND symb_decoder(16#9c#)) OR
 					(reg_q414 AND symb_decoder(16#08#)) OR
 					(reg_q414 AND symb_decoder(16#5e#)) OR
 					(reg_q414 AND symb_decoder(16#dc#)) OR
 					(reg_q414 AND symb_decoder(16#27#)) OR
 					(reg_q414 AND symb_decoder(16#70#)) OR
 					(reg_q414 AND symb_decoder(16#7d#)) OR
 					(reg_q414 AND symb_decoder(16#11#)) OR
 					(reg_q414 AND symb_decoder(16#e4#)) OR
 					(reg_q414 AND symb_decoder(16#69#)) OR
 					(reg_q414 AND symb_decoder(16#aa#)) OR
 					(reg_q414 AND symb_decoder(16#c1#)) OR
 					(reg_q414 AND symb_decoder(16#9f#)) OR
 					(reg_q414 AND symb_decoder(16#0a#)) OR
 					(reg_q414 AND symb_decoder(16#0b#)) OR
 					(reg_q414 AND symb_decoder(16#6c#)) OR
 					(reg_q414 AND symb_decoder(16#84#)) OR
 					(reg_q414 AND symb_decoder(16#fd#)) OR
 					(reg_q414 AND symb_decoder(16#7b#)) OR
 					(reg_q414 AND symb_decoder(16#12#)) OR
 					(reg_q414 AND symb_decoder(16#13#)) OR
 					(reg_q414 AND symb_decoder(16#83#)) OR
 					(reg_q414 AND symb_decoder(16#dd#)) OR
 					(reg_q414 AND symb_decoder(16#25#)) OR
 					(reg_q414 AND symb_decoder(16#c0#)) OR
 					(reg_q414 AND symb_decoder(16#d4#)) OR
 					(reg_q414 AND symb_decoder(16#f2#)) OR
 					(reg_q414 AND symb_decoder(16#48#)) OR
 					(reg_q414 AND symb_decoder(16#6f#)) OR
 					(reg_q414 AND symb_decoder(16#3b#)) OR
 					(reg_q414 AND symb_decoder(16#db#)) OR
 					(reg_q414 AND symb_decoder(16#8d#)) OR
 					(reg_q414 AND symb_decoder(16#ec#)) OR
 					(reg_q414 AND symb_decoder(16#36#)) OR
 					(reg_q414 AND symb_decoder(16#6d#)) OR
 					(reg_q414 AND symb_decoder(16#a9#)) OR
 					(reg_q414 AND symb_decoder(16#c8#)) OR
 					(reg_q414 AND symb_decoder(16#64#)) OR
 					(reg_q414 AND symb_decoder(16#a3#)) OR
 					(reg_q414 AND symb_decoder(16#ba#)) OR
 					(reg_q414 AND symb_decoder(16#5c#)) OR
 					(reg_q414 AND symb_decoder(16#96#)) OR
 					(reg_q414 AND symb_decoder(16#42#)) OR
 					(reg_q414 AND symb_decoder(16#a6#)) OR
 					(reg_q414 AND symb_decoder(16#2f#)) OR
 					(reg_q414 AND symb_decoder(16#86#)) OR
 					(reg_q414 AND symb_decoder(16#9b#)) OR
 					(reg_q414 AND symb_decoder(16#c4#)) OR
 					(reg_q414 AND symb_decoder(16#65#)) OR
 					(reg_q414 AND symb_decoder(16#cc#)) OR
 					(reg_q414 AND symb_decoder(16#73#)) OR
 					(reg_q414 AND symb_decoder(16#09#)) OR
 					(reg_q414 AND symb_decoder(16#5a#)) OR
 					(reg_q414 AND symb_decoder(16#e7#)) OR
 					(reg_q414 AND symb_decoder(16#be#)) OR
 					(reg_q414 AND symb_decoder(16#04#)) OR
 					(reg_q414 AND symb_decoder(16#77#)) OR
 					(reg_q414 AND symb_decoder(16#1d#)) OR
 					(reg_q414 AND symb_decoder(16#78#)) OR
 					(reg_q414 AND symb_decoder(16#8b#)) OR
 					(reg_q414 AND symb_decoder(16#e2#)) OR
 					(reg_q414 AND symb_decoder(16#f6#)) OR
 					(reg_q414 AND symb_decoder(16#33#)) OR
 					(reg_q414 AND symb_decoder(16#ee#)) OR
 					(reg_q414 AND symb_decoder(16#8e#)) OR
 					(reg_q414 AND symb_decoder(16#b5#)) OR
 					(reg_q414 AND symb_decoder(16#6e#)) OR
 					(reg_q414 AND symb_decoder(16#2a#)) OR
 					(reg_q414 AND symb_decoder(16#00#)) OR
 					(reg_q414 AND symb_decoder(16#88#)) OR
 					(reg_q414 AND symb_decoder(16#bd#)) OR
 					(reg_q414 AND symb_decoder(16#54#)) OR
 					(reg_q414 AND symb_decoder(16#cd#)) OR
 					(reg_q414 AND symb_decoder(16#55#)) OR
 					(reg_q414 AND symb_decoder(16#6a#)) OR
 					(reg_q414 AND symb_decoder(16#66#)) OR
 					(reg_q414 AND symb_decoder(16#17#)) OR
 					(reg_q414 AND symb_decoder(16#35#)) OR
 					(reg_q414 AND symb_decoder(16#9a#)) OR
 					(reg_q414 AND symb_decoder(16#10#)) OR
 					(reg_q414 AND symb_decoder(16#21#)) OR
 					(reg_q414 AND symb_decoder(16#44#)) OR
 					(reg_q414 AND symb_decoder(16#82#)) OR
 					(reg_q414 AND symb_decoder(16#fe#)) OR
 					(reg_q414 AND symb_decoder(16#89#)) OR
 					(reg_q414 AND symb_decoder(16#1a#)) OR
 					(reg_q414 AND symb_decoder(16#bc#)) OR
 					(reg_q414 AND symb_decoder(16#71#)) OR
 					(reg_q414 AND symb_decoder(16#a0#)) OR
 					(reg_q414 AND symb_decoder(16#38#)) OR
 					(reg_q414 AND symb_decoder(16#1b#)) OR
 					(reg_q414 AND symb_decoder(16#0d#)) OR
 					(reg_q414 AND symb_decoder(16#7e#)) OR
 					(reg_q414 AND symb_decoder(16#b2#)) OR
 					(reg_q414 AND symb_decoder(16#d1#)) OR
 					(reg_q414 AND symb_decoder(16#e0#)) OR
 					(reg_q414 AND symb_decoder(16#ae#)) OR
 					(reg_q414 AND symb_decoder(16#d6#)) OR
 					(reg_q414 AND symb_decoder(16#95#)) OR
 					(reg_q414 AND symb_decoder(16#45#)) OR
 					(reg_q414 AND symb_decoder(16#37#)) OR
 					(reg_q414 AND symb_decoder(16#30#)) OR
 					(reg_q414 AND symb_decoder(16#0f#)) OR
 					(reg_q414 AND symb_decoder(16#5f#)) OR
 					(reg_q414 AND symb_decoder(16#d5#)) OR
 					(reg_q414 AND symb_decoder(16#3e#)) OR
 					(reg_q414 AND symb_decoder(16#1f#)) OR
 					(reg_q414 AND symb_decoder(16#18#)) OR
 					(reg_q414 AND symb_decoder(16#87#)) OR
 					(reg_q414 AND symb_decoder(16#fc#)) OR
 					(reg_q414 AND symb_decoder(16#32#)) OR
 					(reg_q414 AND symb_decoder(16#23#)) OR
 					(reg_q414 AND symb_decoder(16#a7#)) OR
 					(reg_q414 AND symb_decoder(16#c5#)) OR
 					(reg_q414 AND symb_decoder(16#34#)) OR
 					(reg_q414 AND symb_decoder(16#b6#)) OR
 					(reg_q414 AND symb_decoder(16#58#)) OR
 					(reg_q414 AND symb_decoder(16#9d#)) OR
 					(reg_q414 AND symb_decoder(16#d7#)) OR
 					(reg_q414 AND symb_decoder(16#f7#)) OR
 					(reg_q414 AND symb_decoder(16#e8#)) OR
 					(reg_q414 AND symb_decoder(16#50#)) OR
 					(reg_q414 AND symb_decoder(16#03#)) OR
 					(reg_q414 AND symb_decoder(16#b7#)) OR
 					(reg_q414 AND symb_decoder(16#2b#)) OR
 					(reg_q414 AND symb_decoder(16#c2#)) OR
 					(reg_q414 AND symb_decoder(16#4f#)) OR
 					(reg_q414 AND symb_decoder(16#df#)) OR
 					(reg_q414 AND symb_decoder(16#2e#)) OR
 					(reg_q414 AND symb_decoder(16#c3#)) OR
 					(reg_q414 AND symb_decoder(16#94#)) OR
 					(reg_q414 AND symb_decoder(16#7a#)) OR
 					(reg_q414 AND symb_decoder(16#af#)) OR
 					(reg_q414 AND symb_decoder(16#f9#)) OR
 					(reg_q414 AND symb_decoder(16#68#)) OR
 					(reg_q414 AND symb_decoder(16#f4#)) OR
 					(reg_q414 AND symb_decoder(16#39#)) OR
 					(reg_q414 AND symb_decoder(16#72#)) OR
 					(reg_q414 AND symb_decoder(16#19#)) OR
 					(reg_q414 AND symb_decoder(16#14#)) OR
 					(reg_q414 AND symb_decoder(16#76#)) OR
 					(reg_q414 AND symb_decoder(16#f3#)) OR
 					(reg_q414 AND symb_decoder(16#3c#)) OR
 					(reg_q414 AND symb_decoder(16#97#)) OR
 					(reg_q414 AND symb_decoder(16#15#)) OR
 					(reg_q414 AND symb_decoder(16#3f#)) OR
 					(reg_q414 AND symb_decoder(16#63#)) OR
 					(reg_q414 AND symb_decoder(16#c7#)) OR
 					(reg_q414 AND symb_decoder(16#a1#)) OR
 					(reg_q414 AND symb_decoder(16#40#)) OR
 					(reg_q414 AND symb_decoder(16#57#)) OR
 					(reg_q414 AND symb_decoder(16#b1#)) OR
 					(reg_q414 AND symb_decoder(16#9e#)) OR
 					(reg_q414 AND symb_decoder(16#47#)) OR
 					(reg_q414 AND symb_decoder(16#41#)) OR
 					(reg_q414 AND symb_decoder(16#c9#)) OR
 					(reg_q414 AND symb_decoder(16#60#)) OR
 					(reg_q414 AND symb_decoder(16#1c#)) OR
 					(reg_q414 AND symb_decoder(16#e1#)) OR
 					(reg_q414 AND symb_decoder(16#02#)) OR
 					(reg_q414 AND symb_decoder(16#80#)) OR
 					(reg_q414 AND symb_decoder(16#d0#)) OR
 					(reg_q414 AND symb_decoder(16#6b#)) OR
 					(reg_q414 AND symb_decoder(16#d8#)) OR
 					(reg_q414 AND symb_decoder(16#91#)) OR
 					(reg_q414 AND symb_decoder(16#61#)) OR
 					(reg_q414 AND symb_decoder(16#46#)) OR
 					(reg_q414 AND symb_decoder(16#06#)) OR
 					(reg_q414 AND symb_decoder(16#26#)) OR
 					(reg_q414 AND symb_decoder(16#d3#)) OR
 					(reg_q414 AND symb_decoder(16#4a#)) OR
 					(reg_q414 AND symb_decoder(16#ad#)) OR
 					(reg_q414 AND symb_decoder(16#28#)) OR
 					(reg_q414 AND symb_decoder(16#b8#)) OR
 					(reg_q414 AND symb_decoder(16#31#)) OR
 					(reg_q414 AND symb_decoder(16#4d#)) OR
 					(reg_q414 AND symb_decoder(16#62#)) OR
 					(reg_q414 AND symb_decoder(16#b4#)) OR
 					(reg_q414 AND symb_decoder(16#16#)) OR
 					(reg_q414 AND symb_decoder(16#a2#)) OR
 					(reg_q414 AND symb_decoder(16#67#)) OR
 					(reg_q414 AND symb_decoder(16#b9#)) OR
 					(reg_q414 AND symb_decoder(16#51#)) OR
 					(reg_q414 AND symb_decoder(16#a4#)) OR
 					(reg_q414 AND symb_decoder(16#f5#)) OR
 					(reg_q414 AND symb_decoder(16#2d#)) OR
 					(reg_q414 AND symb_decoder(16#ab#)) OR
 					(reg_q414 AND symb_decoder(16#ea#)) OR
 					(reg_q414 AND symb_decoder(16#81#)) OR
 					(reg_q414 AND symb_decoder(16#a5#)) OR
 					(reg_q414 AND symb_decoder(16#c6#)) OR
 					(reg_q414 AND symb_decoder(16#05#)) OR
 					(reg_q414 AND symb_decoder(16#bb#)) OR
 					(reg_q414 AND symb_decoder(16#01#)) OR
 					(reg_q414 AND symb_decoder(16#5b#)) OR
 					(reg_q414 AND symb_decoder(16#90#)) OR
 					(reg_q414 AND symb_decoder(16#93#)) OR
 					(reg_q414 AND symb_decoder(16#de#)) OR
 					(reg_q414 AND symb_decoder(16#f0#)) OR
 					(reg_q414 AND symb_decoder(16#ef#)) OR
 					(reg_q414 AND symb_decoder(16#ff#)) OR
 					(reg_q414 AND symb_decoder(16#e5#)) OR
 					(reg_q414 AND symb_decoder(16#75#)) OR
 					(reg_q414 AND symb_decoder(16#1e#)) OR
 					(reg_q414 AND symb_decoder(16#7f#)) OR
 					(reg_q414 AND symb_decoder(16#0c#)) OR
 					(reg_q414 AND symb_decoder(16#a8#)) OR
 					(reg_q414 AND symb_decoder(16#85#)) OR
 					(reg_q414 AND symb_decoder(16#4b#)) OR
 					(reg_q414 AND symb_decoder(16#fb#)) OR
 					(reg_q414 AND symb_decoder(16#22#)) OR
 					(reg_q414 AND symb_decoder(16#ca#)) OR
 					(reg_q414 AND symb_decoder(16#4c#)) OR
 					(reg_q414 AND symb_decoder(16#99#)) OR
 					(reg_q414 AND symb_decoder(16#20#)) OR
 					(reg_q414 AND symb_decoder(16#5d#)) OR
 					(reg_q414 AND symb_decoder(16#eb#)) OR
 					(reg_q414 AND symb_decoder(16#ce#)) OR
 					(reg_q414 AND symb_decoder(16#7c#)) OR
 					(reg_q414 AND symb_decoder(16#3d#)) OR
 					(reg_q414 AND symb_decoder(16#b0#)) OR
 					(reg_q414 AND symb_decoder(16#ed#)) OR
 					(reg_q414 AND symb_decoder(16#74#)) OR
 					(reg_q414 AND symb_decoder(16#cb#)) OR
 					(reg_q414 AND symb_decoder(16#e3#)) OR
 					(reg_q414 AND symb_decoder(16#59#)) OR
 					(reg_q414 AND symb_decoder(16#d2#)) OR
 					(reg_q414 AND symb_decoder(16#8c#)) OR
 					(reg_q414 AND symb_decoder(16#24#)) OR
 					(reg_q414 AND symb_decoder(16#07#)) OR
 					(reg_q414 AND symb_decoder(16#92#)) OR
 					(reg_q414 AND symb_decoder(16#43#)) OR
 					(reg_q414 AND symb_decoder(16#e9#)) OR
 					(reg_q414 AND symb_decoder(16#0e#)) OR
 					(reg_q414 AND symb_decoder(16#4e#)) OR
 					(reg_q414 AND symb_decoder(16#98#)) OR
 					(reg_q414 AND symb_decoder(16#29#)) OR
 					(reg_q414 AND symb_decoder(16#bf#)) OR
 					(reg_q414 AND symb_decoder(16#56#)) OR
 					(reg_q414 AND symb_decoder(16#52#)) OR
 					(reg_q414 AND symb_decoder(16#53#)) OR
 					(reg_q414 AND symb_decoder(16#da#)) OR
 					(reg_q414 AND symb_decoder(16#49#)) OR
 					(reg_q414 AND symb_decoder(16#ac#)) OR
 					(reg_q414 AND symb_decoder(16#d9#)) OR
 					(reg_q414 AND symb_decoder(16#e6#));
reg_q414_init <= '0' ;
	p_reg_q414: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q414 <= reg_q414_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q414 <= reg_q414_init;
        else
          reg_q414 <= reg_q414_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2252_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2252 AND symb_decoder(16#79#)) OR
 					(reg_q2252 AND symb_decoder(16#ad#)) OR
 					(reg_q2252 AND symb_decoder(16#07#)) OR
 					(reg_q2252 AND symb_decoder(16#a1#)) OR
 					(reg_q2252 AND symb_decoder(16#67#)) OR
 					(reg_q2252 AND symb_decoder(16#23#)) OR
 					(reg_q2252 AND symb_decoder(16#cc#)) OR
 					(reg_q2252 AND symb_decoder(16#43#)) OR
 					(reg_q2252 AND symb_decoder(16#48#)) OR
 					(reg_q2252 AND symb_decoder(16#3e#)) OR
 					(reg_q2252 AND symb_decoder(16#45#)) OR
 					(reg_q2252 AND symb_decoder(16#26#)) OR
 					(reg_q2252 AND symb_decoder(16#c3#)) OR
 					(reg_q2252 AND symb_decoder(16#e3#)) OR
 					(reg_q2252 AND symb_decoder(16#8b#)) OR
 					(reg_q2252 AND symb_decoder(16#e7#)) OR
 					(reg_q2252 AND symb_decoder(16#b8#)) OR
 					(reg_q2252 AND symb_decoder(16#ba#)) OR
 					(reg_q2252 AND symb_decoder(16#60#)) OR
 					(reg_q2252 AND symb_decoder(16#3b#)) OR
 					(reg_q2252 AND symb_decoder(16#b3#)) OR
 					(reg_q2252 AND symb_decoder(16#90#)) OR
 					(reg_q2252 AND symb_decoder(16#19#)) OR
 					(reg_q2252 AND symb_decoder(16#df#)) OR
 					(reg_q2252 AND symb_decoder(16#f8#)) OR
 					(reg_q2252 AND symb_decoder(16#0d#)) OR
 					(reg_q2252 AND symb_decoder(16#5f#)) OR
 					(reg_q2252 AND symb_decoder(16#8e#)) OR
 					(reg_q2252 AND symb_decoder(16#58#)) OR
 					(reg_q2252 AND symb_decoder(16#18#)) OR
 					(reg_q2252 AND symb_decoder(16#ab#)) OR
 					(reg_q2252 AND symb_decoder(16#61#)) OR
 					(reg_q2252 AND symb_decoder(16#25#)) OR
 					(reg_q2252 AND symb_decoder(16#13#)) OR
 					(reg_q2252 AND symb_decoder(16#1b#)) OR
 					(reg_q2252 AND symb_decoder(16#fd#)) OR
 					(reg_q2252 AND symb_decoder(16#22#)) OR
 					(reg_q2252 AND symb_decoder(16#2e#)) OR
 					(reg_q2252 AND symb_decoder(16#4e#)) OR
 					(reg_q2252 AND symb_decoder(16#7e#)) OR
 					(reg_q2252 AND symb_decoder(16#76#)) OR
 					(reg_q2252 AND symb_decoder(16#85#)) OR
 					(reg_q2252 AND symb_decoder(16#f1#)) OR
 					(reg_q2252 AND symb_decoder(16#a5#)) OR
 					(reg_q2252 AND symb_decoder(16#3f#)) OR
 					(reg_q2252 AND symb_decoder(16#0c#)) OR
 					(reg_q2252 AND symb_decoder(16#47#)) OR
 					(reg_q2252 AND symb_decoder(16#a8#)) OR
 					(reg_q2252 AND symb_decoder(16#f9#)) OR
 					(reg_q2252 AND symb_decoder(16#6f#)) OR
 					(reg_q2252 AND symb_decoder(16#b5#)) OR
 					(reg_q2252 AND symb_decoder(16#b2#)) OR
 					(reg_q2252 AND symb_decoder(16#27#)) OR
 					(reg_q2252 AND symb_decoder(16#64#)) OR
 					(reg_q2252 AND symb_decoder(16#77#)) OR
 					(reg_q2252 AND symb_decoder(16#c9#)) OR
 					(reg_q2252 AND symb_decoder(16#65#)) OR
 					(reg_q2252 AND symb_decoder(16#6b#)) OR
 					(reg_q2252 AND symb_decoder(16#c4#)) OR
 					(reg_q2252 AND symb_decoder(16#bf#)) OR
 					(reg_q2252 AND symb_decoder(16#96#)) OR
 					(reg_q2252 AND symb_decoder(16#fe#)) OR
 					(reg_q2252 AND symb_decoder(16#bc#)) OR
 					(reg_q2252 AND symb_decoder(16#1c#)) OR
 					(reg_q2252 AND symb_decoder(16#b4#)) OR
 					(reg_q2252 AND symb_decoder(16#40#)) OR
 					(reg_q2252 AND symb_decoder(16#8c#)) OR
 					(reg_q2252 AND symb_decoder(16#3c#)) OR
 					(reg_q2252 AND symb_decoder(16#6c#)) OR
 					(reg_q2252 AND symb_decoder(16#89#)) OR
 					(reg_q2252 AND symb_decoder(16#ec#)) OR
 					(reg_q2252 AND symb_decoder(16#4f#)) OR
 					(reg_q2252 AND symb_decoder(16#5e#)) OR
 					(reg_q2252 AND symb_decoder(16#1f#)) OR
 					(reg_q2252 AND symb_decoder(16#2d#)) OR
 					(reg_q2252 AND symb_decoder(16#80#)) OR
 					(reg_q2252 AND symb_decoder(16#69#)) OR
 					(reg_q2252 AND symb_decoder(16#0e#)) OR
 					(reg_q2252 AND symb_decoder(16#ed#)) OR
 					(reg_q2252 AND symb_decoder(16#4b#)) OR
 					(reg_q2252 AND symb_decoder(16#e5#)) OR
 					(reg_q2252 AND symb_decoder(16#5c#)) OR
 					(reg_q2252 AND symb_decoder(16#b6#)) OR
 					(reg_q2252 AND symb_decoder(16#d1#)) OR
 					(reg_q2252 AND symb_decoder(16#d9#)) OR
 					(reg_q2252 AND symb_decoder(16#32#)) OR
 					(reg_q2252 AND symb_decoder(16#ac#)) OR
 					(reg_q2252 AND symb_decoder(16#33#)) OR
 					(reg_q2252 AND symb_decoder(16#b1#)) OR
 					(reg_q2252 AND symb_decoder(16#36#)) OR
 					(reg_q2252 AND symb_decoder(16#28#)) OR
 					(reg_q2252 AND symb_decoder(16#d2#)) OR
 					(reg_q2252 AND symb_decoder(16#6a#)) OR
 					(reg_q2252 AND symb_decoder(16#f3#)) OR
 					(reg_q2252 AND symb_decoder(16#af#)) OR
 					(reg_q2252 AND symb_decoder(16#9a#)) OR
 					(reg_q2252 AND symb_decoder(16#49#)) OR
 					(reg_q2252 AND symb_decoder(16#c5#)) OR
 					(reg_q2252 AND symb_decoder(16#75#)) OR
 					(reg_q2252 AND symb_decoder(16#ee#)) OR
 					(reg_q2252 AND symb_decoder(16#81#)) OR
 					(reg_q2252 AND symb_decoder(16#63#)) OR
 					(reg_q2252 AND symb_decoder(16#ef#)) OR
 					(reg_q2252 AND symb_decoder(16#00#)) OR
 					(reg_q2252 AND symb_decoder(16#87#)) OR
 					(reg_q2252 AND symb_decoder(16#5a#)) OR
 					(reg_q2252 AND symb_decoder(16#38#)) OR
 					(reg_q2252 AND symb_decoder(16#b9#)) OR
 					(reg_q2252 AND symb_decoder(16#2c#)) OR
 					(reg_q2252 AND symb_decoder(16#db#)) OR
 					(reg_q2252 AND symb_decoder(16#f5#)) OR
 					(reg_q2252 AND symb_decoder(16#c7#)) OR
 					(reg_q2252 AND symb_decoder(16#d0#)) OR
 					(reg_q2252 AND symb_decoder(16#3d#)) OR
 					(reg_q2252 AND symb_decoder(16#72#)) OR
 					(reg_q2252 AND symb_decoder(16#31#)) OR
 					(reg_q2252 AND symb_decoder(16#78#)) OR
 					(reg_q2252 AND symb_decoder(16#e0#)) OR
 					(reg_q2252 AND symb_decoder(16#e6#)) OR
 					(reg_q2252 AND symb_decoder(16#54#)) OR
 					(reg_q2252 AND symb_decoder(16#cd#)) OR
 					(reg_q2252 AND symb_decoder(16#a0#)) OR
 					(reg_q2252 AND symb_decoder(16#f0#)) OR
 					(reg_q2252 AND symb_decoder(16#99#)) OR
 					(reg_q2252 AND symb_decoder(16#d8#)) OR
 					(reg_q2252 AND symb_decoder(16#94#)) OR
 					(reg_q2252 AND symb_decoder(16#95#)) OR
 					(reg_q2252 AND symb_decoder(16#cf#)) OR
 					(reg_q2252 AND symb_decoder(16#12#)) OR
 					(reg_q2252 AND symb_decoder(16#d4#)) OR
 					(reg_q2252 AND symb_decoder(16#c0#)) OR
 					(reg_q2252 AND symb_decoder(16#92#)) OR
 					(reg_q2252 AND symb_decoder(16#24#)) OR
 					(reg_q2252 AND symb_decoder(16#a4#)) OR
 					(reg_q2252 AND symb_decoder(16#01#)) OR
 					(reg_q2252 AND symb_decoder(16#ea#)) OR
 					(reg_q2252 AND symb_decoder(16#70#)) OR
 					(reg_q2252 AND symb_decoder(16#44#)) OR
 					(reg_q2252 AND symb_decoder(16#2a#)) OR
 					(reg_q2252 AND symb_decoder(16#39#)) OR
 					(reg_q2252 AND symb_decoder(16#f6#)) OR
 					(reg_q2252 AND symb_decoder(16#aa#)) OR
 					(reg_q2252 AND symb_decoder(16#1e#)) OR
 					(reg_q2252 AND symb_decoder(16#fa#)) OR
 					(reg_q2252 AND symb_decoder(16#bd#)) OR
 					(reg_q2252 AND symb_decoder(16#10#)) OR
 					(reg_q2252 AND symb_decoder(16#ff#)) OR
 					(reg_q2252 AND symb_decoder(16#30#)) OR
 					(reg_q2252 AND symb_decoder(16#9e#)) OR
 					(reg_q2252 AND symb_decoder(16#71#)) OR
 					(reg_q2252 AND symb_decoder(16#0f#)) OR
 					(reg_q2252 AND symb_decoder(16#05#)) OR
 					(reg_q2252 AND symb_decoder(16#50#)) OR
 					(reg_q2252 AND symb_decoder(16#62#)) OR
 					(reg_q2252 AND symb_decoder(16#be#)) OR
 					(reg_q2252 AND symb_decoder(16#ce#)) OR
 					(reg_q2252 AND symb_decoder(16#f7#)) OR
 					(reg_q2252 AND symb_decoder(16#82#)) OR
 					(reg_q2252 AND symb_decoder(16#4a#)) OR
 					(reg_q2252 AND symb_decoder(16#9b#)) OR
 					(reg_q2252 AND symb_decoder(16#2b#)) OR
 					(reg_q2252 AND symb_decoder(16#b0#)) OR
 					(reg_q2252 AND symb_decoder(16#7a#)) OR
 					(reg_q2252 AND symb_decoder(16#08#)) OR
 					(reg_q2252 AND symb_decoder(16#e9#)) OR
 					(reg_q2252 AND symb_decoder(16#59#)) OR
 					(reg_q2252 AND symb_decoder(16#3a#)) OR
 					(reg_q2252 AND symb_decoder(16#c8#)) OR
 					(reg_q2252 AND symb_decoder(16#a3#)) OR
 					(reg_q2252 AND symb_decoder(16#11#)) OR
 					(reg_q2252 AND symb_decoder(16#29#)) OR
 					(reg_q2252 AND symb_decoder(16#6d#)) OR
 					(reg_q2252 AND symb_decoder(16#66#)) OR
 					(reg_q2252 AND symb_decoder(16#57#)) OR
 					(reg_q2252 AND symb_decoder(16#14#)) OR
 					(reg_q2252 AND symb_decoder(16#51#)) OR
 					(reg_q2252 AND symb_decoder(16#c1#)) OR
 					(reg_q2252 AND symb_decoder(16#da#)) OR
 					(reg_q2252 AND symb_decoder(16#37#)) OR
 					(reg_q2252 AND symb_decoder(16#56#)) OR
 					(reg_q2252 AND symb_decoder(16#17#)) OR
 					(reg_q2252 AND symb_decoder(16#91#)) OR
 					(reg_q2252 AND symb_decoder(16#9c#)) OR
 					(reg_q2252 AND symb_decoder(16#9d#)) OR
 					(reg_q2252 AND symb_decoder(16#a6#)) OR
 					(reg_q2252 AND symb_decoder(16#ca#)) OR
 					(reg_q2252 AND symb_decoder(16#2f#)) OR
 					(reg_q2252 AND symb_decoder(16#e2#)) OR
 					(reg_q2252 AND symb_decoder(16#74#)) OR
 					(reg_q2252 AND symb_decoder(16#8a#)) OR
 					(reg_q2252 AND symb_decoder(16#35#)) OR
 					(reg_q2252 AND symb_decoder(16#03#)) OR
 					(reg_q2252 AND symb_decoder(16#f2#)) OR
 					(reg_q2252 AND symb_decoder(16#bb#)) OR
 					(reg_q2252 AND symb_decoder(16#84#)) OR
 					(reg_q2252 AND symb_decoder(16#e1#)) OR
 					(reg_q2252 AND symb_decoder(16#0a#)) OR
 					(reg_q2252 AND symb_decoder(16#5d#)) OR
 					(reg_q2252 AND symb_decoder(16#eb#)) OR
 					(reg_q2252 AND symb_decoder(16#88#)) OR
 					(reg_q2252 AND symb_decoder(16#53#)) OR
 					(reg_q2252 AND symb_decoder(16#02#)) OR
 					(reg_q2252 AND symb_decoder(16#98#)) OR
 					(reg_q2252 AND symb_decoder(16#55#)) OR
 					(reg_q2252 AND symb_decoder(16#e8#)) OR
 					(reg_q2252 AND symb_decoder(16#6e#)) OR
 					(reg_q2252 AND symb_decoder(16#fc#)) OR
 					(reg_q2252 AND symb_decoder(16#c6#)) OR
 					(reg_q2252 AND symb_decoder(16#04#)) OR
 					(reg_q2252 AND symb_decoder(16#c2#)) OR
 					(reg_q2252 AND symb_decoder(16#1a#)) OR
 					(reg_q2252 AND symb_decoder(16#68#)) OR
 					(reg_q2252 AND symb_decoder(16#f4#)) OR
 					(reg_q2252 AND symb_decoder(16#4c#)) OR
 					(reg_q2252 AND symb_decoder(16#4d#)) OR
 					(reg_q2252 AND symb_decoder(16#83#)) OR
 					(reg_q2252 AND symb_decoder(16#ae#)) OR
 					(reg_q2252 AND symb_decoder(16#7c#)) OR
 					(reg_q2252 AND symb_decoder(16#d6#)) OR
 					(reg_q2252 AND symb_decoder(16#fb#)) OR
 					(reg_q2252 AND symb_decoder(16#34#)) OR
 					(reg_q2252 AND symb_decoder(16#e4#)) OR
 					(reg_q2252 AND symb_decoder(16#7d#)) OR
 					(reg_q2252 AND symb_decoder(16#8d#)) OR
 					(reg_q2252 AND symb_decoder(16#a7#)) OR
 					(reg_q2252 AND symb_decoder(16#93#)) OR
 					(reg_q2252 AND symb_decoder(16#0b#)) OR
 					(reg_q2252 AND symb_decoder(16#73#)) OR
 					(reg_q2252 AND symb_decoder(16#b7#)) OR
 					(reg_q2252 AND symb_decoder(16#20#)) OR
 					(reg_q2252 AND symb_decoder(16#15#)) OR
 					(reg_q2252 AND symb_decoder(16#42#)) OR
 					(reg_q2252 AND symb_decoder(16#d5#)) OR
 					(reg_q2252 AND symb_decoder(16#7b#)) OR
 					(reg_q2252 AND symb_decoder(16#dd#)) OR
 					(reg_q2252 AND symb_decoder(16#52#)) OR
 					(reg_q2252 AND symb_decoder(16#8f#)) OR
 					(reg_q2252 AND symb_decoder(16#de#)) OR
 					(reg_q2252 AND symb_decoder(16#21#)) OR
 					(reg_q2252 AND symb_decoder(16#a9#)) OR
 					(reg_q2252 AND symb_decoder(16#d3#)) OR
 					(reg_q2252 AND symb_decoder(16#dc#)) OR
 					(reg_q2252 AND symb_decoder(16#cb#)) OR
 					(reg_q2252 AND symb_decoder(16#9f#)) OR
 					(reg_q2252 AND symb_decoder(16#5b#)) OR
 					(reg_q2252 AND symb_decoder(16#41#)) OR
 					(reg_q2252 AND symb_decoder(16#97#)) OR
 					(reg_q2252 AND symb_decoder(16#d7#)) OR
 					(reg_q2252 AND symb_decoder(16#06#)) OR
 					(reg_q2252 AND symb_decoder(16#a2#)) OR
 					(reg_q2252 AND symb_decoder(16#7f#)) OR
 					(reg_q2252 AND symb_decoder(16#86#)) OR
 					(reg_q2252 AND symb_decoder(16#09#)) OR
 					(reg_q2252 AND symb_decoder(16#46#)) OR
 					(reg_q2252 AND symb_decoder(16#16#)) OR
 					(reg_q2252 AND symb_decoder(16#1d#));
reg_q2252_init <= '0' ;
	p_reg_q2252: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2252 <= reg_q2252_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2252 <= reg_q2252_init;
        else
          reg_q2252 <= reg_q2252_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph43

reg_q1772_in <= (reg_q1770 AND symb_decoder(16#0a#)) OR
 					(reg_q1770 AND symb_decoder(16#20#)) OR
 					(reg_q1770 AND symb_decoder(16#09#)) OR
 					(reg_q1770 AND symb_decoder(16#0c#)) OR
 					(reg_q1770 AND symb_decoder(16#0d#));
reg_q618_in <= (reg_q616 AND symb_decoder(16#16#)) OR
 					(reg_q616 AND symb_decoder(16#01#)) OR
 					(reg_q616 AND symb_decoder(16#17#)) OR
 					(reg_q616 AND symb_decoder(16#31#)) OR
 					(reg_q616 AND symb_decoder(16#5c#)) OR
 					(reg_q616 AND symb_decoder(16#a1#)) OR
 					(reg_q616 AND symb_decoder(16#e6#)) OR
 					(reg_q616 AND symb_decoder(16#58#)) OR
 					(reg_q616 AND symb_decoder(16#ae#)) OR
 					(reg_q616 AND symb_decoder(16#00#)) OR
 					(reg_q616 AND symb_decoder(16#1f#)) OR
 					(reg_q616 AND symb_decoder(16#b9#)) OR
 					(reg_q616 AND symb_decoder(16#fb#)) OR
 					(reg_q616 AND symb_decoder(16#b0#)) OR
 					(reg_q616 AND symb_decoder(16#de#)) OR
 					(reg_q616 AND symb_decoder(16#35#)) OR
 					(reg_q616 AND symb_decoder(16#a0#)) OR
 					(reg_q616 AND symb_decoder(16#aa#)) OR
 					(reg_q616 AND symb_decoder(16#db#)) OR
 					(reg_q616 AND symb_decoder(16#2d#)) OR
 					(reg_q616 AND symb_decoder(16#57#)) OR
 					(reg_q616 AND symb_decoder(16#cc#)) OR
 					(reg_q616 AND symb_decoder(16#1b#)) OR
 					(reg_q616 AND symb_decoder(16#88#)) OR
 					(reg_q616 AND symb_decoder(16#48#)) OR
 					(reg_q616 AND symb_decoder(16#6b#)) OR
 					(reg_q616 AND symb_decoder(16#30#)) OR
 					(reg_q616 AND symb_decoder(16#e5#)) OR
 					(reg_q616 AND symb_decoder(16#98#)) OR
 					(reg_q616 AND symb_decoder(16#63#)) OR
 					(reg_q616 AND symb_decoder(16#f4#)) OR
 					(reg_q616 AND symb_decoder(16#d7#)) OR
 					(reg_q616 AND symb_decoder(16#f8#)) OR
 					(reg_q616 AND symb_decoder(16#8f#)) OR
 					(reg_q616 AND symb_decoder(16#e7#)) OR
 					(reg_q616 AND symb_decoder(16#0e#)) OR
 					(reg_q616 AND symb_decoder(16#bd#)) OR
 					(reg_q616 AND symb_decoder(16#d4#)) OR
 					(reg_q616 AND symb_decoder(16#9f#)) OR
 					(reg_q616 AND symb_decoder(16#84#)) OR
 					(reg_q616 AND symb_decoder(16#1e#)) OR
 					(reg_q616 AND symb_decoder(16#ff#)) OR
 					(reg_q616 AND symb_decoder(16#f1#)) OR
 					(reg_q616 AND symb_decoder(16#a7#)) OR
 					(reg_q616 AND symb_decoder(16#56#)) OR
 					(reg_q616 AND symb_decoder(16#32#)) OR
 					(reg_q616 AND symb_decoder(16#94#)) OR
 					(reg_q616 AND symb_decoder(16#7e#)) OR
 					(reg_q616 AND symb_decoder(16#d9#)) OR
 					(reg_q616 AND symb_decoder(16#a8#)) OR
 					(reg_q616 AND symb_decoder(16#7f#)) OR
 					(reg_q616 AND symb_decoder(16#ef#)) OR
 					(reg_q616 AND symb_decoder(16#87#)) OR
 					(reg_q616 AND symb_decoder(16#5f#)) OR
 					(reg_q616 AND symb_decoder(16#cd#)) OR
 					(reg_q616 AND symb_decoder(16#54#)) OR
 					(reg_q616 AND symb_decoder(16#fa#)) OR
 					(reg_q616 AND symb_decoder(16#b7#)) OR
 					(reg_q616 AND symb_decoder(16#10#)) OR
 					(reg_q616 AND symb_decoder(16#51#)) OR
 					(reg_q616 AND symb_decoder(16#52#)) OR
 					(reg_q616 AND symb_decoder(16#be#)) OR
 					(reg_q616 AND symb_decoder(16#8a#)) OR
 					(reg_q616 AND symb_decoder(16#7d#)) OR
 					(reg_q616 AND symb_decoder(16#4a#)) OR
 					(reg_q616 AND symb_decoder(16#38#)) OR
 					(reg_q616 AND symb_decoder(16#03#)) OR
 					(reg_q616 AND symb_decoder(16#fd#)) OR
 					(reg_q616 AND symb_decoder(16#85#)) OR
 					(reg_q616 AND symb_decoder(16#92#)) OR
 					(reg_q616 AND symb_decoder(16#33#)) OR
 					(reg_q616 AND symb_decoder(16#42#)) OR
 					(reg_q616 AND symb_decoder(16#c2#)) OR
 					(reg_q616 AND symb_decoder(16#eb#)) OR
 					(reg_q616 AND symb_decoder(16#d2#)) OR
 					(reg_q616 AND symb_decoder(16#b8#)) OR
 					(reg_q616 AND symb_decoder(16#ec#)) OR
 					(reg_q616 AND symb_decoder(16#45#)) OR
 					(reg_q616 AND symb_decoder(16#91#)) OR
 					(reg_q616 AND symb_decoder(16#71#)) OR
 					(reg_q616 AND symb_decoder(16#5e#)) OR
 					(reg_q616 AND symb_decoder(16#24#)) OR
 					(reg_q616 AND symb_decoder(16#21#)) OR
 					(reg_q616 AND symb_decoder(16#75#)) OR
 					(reg_q616 AND symb_decoder(16#a2#)) OR
 					(reg_q616 AND symb_decoder(16#50#)) OR
 					(reg_q616 AND symb_decoder(16#2a#)) OR
 					(reg_q616 AND symb_decoder(16#c0#)) OR
 					(reg_q616 AND symb_decoder(16#59#)) OR
 					(reg_q616 AND symb_decoder(16#c5#)) OR
 					(reg_q616 AND symb_decoder(16#11#)) OR
 					(reg_q616 AND symb_decoder(16#14#)) OR
 					(reg_q616 AND symb_decoder(16#0b#)) OR
 					(reg_q616 AND symb_decoder(16#18#)) OR
 					(reg_q616 AND symb_decoder(16#41#)) OR
 					(reg_q616 AND symb_decoder(16#3f#)) OR
 					(reg_q616 AND symb_decoder(16#8e#)) OR
 					(reg_q616 AND symb_decoder(16#74#)) OR
 					(reg_q616 AND symb_decoder(16#c8#)) OR
 					(reg_q616 AND symb_decoder(16#a9#)) OR
 					(reg_q616 AND symb_decoder(16#89#)) OR
 					(reg_q616 AND symb_decoder(16#49#)) OR
 					(reg_q616 AND symb_decoder(16#fe#)) OR
 					(reg_q616 AND symb_decoder(16#60#)) OR
 					(reg_q616 AND symb_decoder(16#44#)) OR
 					(reg_q616 AND symb_decoder(16#ab#)) OR
 					(reg_q616 AND symb_decoder(16#ce#)) OR
 					(reg_q616 AND symb_decoder(16#68#)) OR
 					(reg_q616 AND symb_decoder(16#cb#)) OR
 					(reg_q616 AND symb_decoder(16#cf#)) OR
 					(reg_q616 AND symb_decoder(16#43#)) OR
 					(reg_q616 AND symb_decoder(16#28#)) OR
 					(reg_q616 AND symb_decoder(16#a6#)) OR
 					(reg_q616 AND symb_decoder(16#04#)) OR
 					(reg_q616 AND symb_decoder(16#90#)) OR
 					(reg_q616 AND symb_decoder(16#bf#)) OR
 					(reg_q616 AND symb_decoder(16#64#)) OR
 					(reg_q616 AND symb_decoder(16#df#)) OR
 					(reg_q616 AND symb_decoder(16#c9#)) OR
 					(reg_q616 AND symb_decoder(16#23#)) OR
 					(reg_q616 AND symb_decoder(16#15#)) OR
 					(reg_q616 AND symb_decoder(16#d6#)) OR
 					(reg_q616 AND symb_decoder(16#6f#)) OR
 					(reg_q616 AND symb_decoder(16#b5#)) OR
 					(reg_q616 AND symb_decoder(16#4d#)) OR
 					(reg_q616 AND symb_decoder(16#e8#)) OR
 					(reg_q616 AND symb_decoder(16#b2#)) OR
 					(reg_q616 AND symb_decoder(16#ea#)) OR
 					(reg_q616 AND symb_decoder(16#86#)) OR
 					(reg_q616 AND symb_decoder(16#08#)) OR
 					(reg_q616 AND symb_decoder(16#47#)) OR
 					(reg_q616 AND symb_decoder(16#6d#)) OR
 					(reg_q616 AND symb_decoder(16#37#)) OR
 					(reg_q616 AND symb_decoder(16#7c#)) OR
 					(reg_q616 AND symb_decoder(16#0f#)) OR
 					(reg_q616 AND symb_decoder(16#53#)) OR
 					(reg_q616 AND symb_decoder(16#79#)) OR
 					(reg_q616 AND symb_decoder(16#76#)) OR
 					(reg_q616 AND symb_decoder(16#06#)) OR
 					(reg_q616 AND symb_decoder(16#4c#)) OR
 					(reg_q616 AND symb_decoder(16#83#)) OR
 					(reg_q616 AND symb_decoder(16#9a#)) OR
 					(reg_q616 AND symb_decoder(16#19#)) OR
 					(reg_q616 AND symb_decoder(16#7a#)) OR
 					(reg_q616 AND symb_decoder(16#6a#)) OR
 					(reg_q616 AND symb_decoder(16#05#)) OR
 					(reg_q616 AND symb_decoder(16#e2#)) OR
 					(reg_q616 AND symb_decoder(16#3c#)) OR
 					(reg_q616 AND symb_decoder(16#9d#)) OR
 					(reg_q616 AND symb_decoder(16#95#)) OR
 					(reg_q616 AND symb_decoder(16#8c#)) OR
 					(reg_q616 AND symb_decoder(16#39#)) OR
 					(reg_q616 AND symb_decoder(16#3e#)) OR
 					(reg_q616 AND symb_decoder(16#7b#)) OR
 					(reg_q616 AND symb_decoder(16#81#)) OR
 					(reg_q616 AND symb_decoder(16#2e#)) OR
 					(reg_q616 AND symb_decoder(16#25#)) OR
 					(reg_q616 AND symb_decoder(16#8b#)) OR
 					(reg_q616 AND symb_decoder(16#5a#)) OR
 					(reg_q616 AND symb_decoder(16#4f#)) OR
 					(reg_q616 AND symb_decoder(16#97#)) OR
 					(reg_q616 AND symb_decoder(16#2f#)) OR
 					(reg_q616 AND symb_decoder(16#da#)) OR
 					(reg_q616 AND symb_decoder(16#8d#)) OR
 					(reg_q616 AND symb_decoder(16#e3#)) OR
 					(reg_q616 AND symb_decoder(16#ee#)) OR
 					(reg_q616 AND symb_decoder(16#70#)) OR
 					(reg_q616 AND symb_decoder(16#f6#)) OR
 					(reg_q616 AND symb_decoder(16#40#)) OR
 					(reg_q616 AND symb_decoder(16#93#)) OR
 					(reg_q616 AND symb_decoder(16#e0#)) OR
 					(reg_q616 AND symb_decoder(16#ac#)) OR
 					(reg_q616 AND symb_decoder(16#e9#)) OR
 					(reg_q616 AND symb_decoder(16#ad#)) OR
 					(reg_q616 AND symb_decoder(16#c3#)) OR
 					(reg_q616 AND symb_decoder(16#d8#)) OR
 					(reg_q616 AND symb_decoder(16#34#)) OR
 					(reg_q616 AND symb_decoder(16#02#)) OR
 					(reg_q616 AND symb_decoder(16#f3#)) OR
 					(reg_q616 AND symb_decoder(16#f5#)) OR
 					(reg_q616 AND symb_decoder(16#1d#)) OR
 					(reg_q616 AND symb_decoder(16#5b#)) OR
 					(reg_q616 AND symb_decoder(16#4e#)) OR
 					(reg_q616 AND symb_decoder(16#a4#)) OR
 					(reg_q616 AND symb_decoder(16#69#)) OR
 					(reg_q616 AND symb_decoder(16#b3#)) OR
 					(reg_q616 AND symb_decoder(16#6c#)) OR
 					(reg_q616 AND symb_decoder(16#66#)) OR
 					(reg_q616 AND symb_decoder(16#f0#)) OR
 					(reg_q616 AND symb_decoder(16#82#)) OR
 					(reg_q616 AND symb_decoder(16#46#)) OR
 					(reg_q616 AND symb_decoder(16#af#)) OR
 					(reg_q616 AND symb_decoder(16#f7#)) OR
 					(reg_q616 AND symb_decoder(16#1c#)) OR
 					(reg_q616 AND symb_decoder(16#e4#)) OR
 					(reg_q616 AND symb_decoder(16#dc#)) OR
 					(reg_q616 AND symb_decoder(16#27#)) OR
 					(reg_q616 AND symb_decoder(16#3d#)) OR
 					(reg_q616 AND symb_decoder(16#b6#)) OR
 					(reg_q616 AND symb_decoder(16#4b#)) OR
 					(reg_q616 AND symb_decoder(16#65#)) OR
 					(reg_q616 AND symb_decoder(16#36#)) OR
 					(reg_q616 AND symb_decoder(16#61#)) OR
 					(reg_q616 AND symb_decoder(16#ba#)) OR
 					(reg_q616 AND symb_decoder(16#c6#)) OR
 					(reg_q616 AND symb_decoder(16#f9#)) OR
 					(reg_q616 AND symb_decoder(16#07#)) OR
 					(reg_q616 AND symb_decoder(16#96#)) OR
 					(reg_q616 AND symb_decoder(16#13#)) OR
 					(reg_q616 AND symb_decoder(16#67#)) OR
 					(reg_q616 AND symb_decoder(16#dd#)) OR
 					(reg_q616 AND symb_decoder(16#2b#)) OR
 					(reg_q616 AND symb_decoder(16#c7#)) OR
 					(reg_q616 AND symb_decoder(16#3a#)) OR
 					(reg_q616 AND symb_decoder(16#bc#)) OR
 					(reg_q616 AND symb_decoder(16#78#)) OR
 					(reg_q616 AND symb_decoder(16#9e#)) OR
 					(reg_q616 AND symb_decoder(16#1a#)) OR
 					(reg_q616 AND symb_decoder(16#e1#)) OR
 					(reg_q616 AND symb_decoder(16#bb#)) OR
 					(reg_q616 AND symb_decoder(16#62#)) OR
 					(reg_q616 AND symb_decoder(16#a3#)) OR
 					(reg_q616 AND symb_decoder(16#d1#)) OR
 					(reg_q616 AND symb_decoder(16#5d#)) OR
 					(reg_q616 AND symb_decoder(16#9c#)) OR
 					(reg_q616 AND symb_decoder(16#d3#)) OR
 					(reg_q616 AND symb_decoder(16#ed#)) OR
 					(reg_q616 AND symb_decoder(16#a5#)) OR
 					(reg_q616 AND symb_decoder(16#c1#)) OR
 					(reg_q616 AND symb_decoder(16#99#)) OR
 					(reg_q616 AND symb_decoder(16#26#)) OR
 					(reg_q616 AND symb_decoder(16#12#)) OR
 					(reg_q616 AND symb_decoder(16#29#)) OR
 					(reg_q616 AND symb_decoder(16#77#)) OR
 					(reg_q616 AND symb_decoder(16#d0#)) OR
 					(reg_q616 AND symb_decoder(16#9b#)) OR
 					(reg_q616 AND symb_decoder(16#2c#)) OR
 					(reg_q616 AND symb_decoder(16#c4#)) OR
 					(reg_q616 AND symb_decoder(16#f2#)) OR
 					(reg_q616 AND symb_decoder(16#b4#)) OR
 					(reg_q616 AND symb_decoder(16#72#)) OR
 					(reg_q616 AND symb_decoder(16#b1#)) OR
 					(reg_q616 AND symb_decoder(16#80#)) OR
 					(reg_q616 AND symb_decoder(16#6e#)) OR
 					(reg_q616 AND symb_decoder(16#55#)) OR
 					(reg_q616 AND symb_decoder(16#73#)) OR
 					(reg_q616 AND symb_decoder(16#fc#)) OR
 					(reg_q616 AND symb_decoder(16#3b#)) OR
 					(reg_q616 AND symb_decoder(16#d5#)) OR
 					(reg_q616 AND symb_decoder(16#22#)) OR
 					(reg_q616 AND symb_decoder(16#ca#)) OR
 					(reg_q618 AND symb_decoder(16#fc#)) OR
 					(reg_q618 AND symb_decoder(16#e9#)) OR
 					(reg_q618 AND symb_decoder(16#e0#)) OR
 					(reg_q618 AND symb_decoder(16#4b#)) OR
 					(reg_q618 AND symb_decoder(16#b7#)) OR
 					(reg_q618 AND symb_decoder(16#02#)) OR
 					(reg_q618 AND symb_decoder(16#71#)) OR
 					(reg_q618 AND symb_decoder(16#e2#)) OR
 					(reg_q618 AND symb_decoder(16#51#)) OR
 					(reg_q618 AND symb_decoder(16#48#)) OR
 					(reg_q618 AND symb_decoder(16#6c#)) OR
 					(reg_q618 AND symb_decoder(16#59#)) OR
 					(reg_q618 AND symb_decoder(16#5f#)) OR
 					(reg_q618 AND symb_decoder(16#d3#)) OR
 					(reg_q618 AND symb_decoder(16#70#)) OR
 					(reg_q618 AND symb_decoder(16#36#)) OR
 					(reg_q618 AND symb_decoder(16#68#)) OR
 					(reg_q618 AND symb_decoder(16#fe#)) OR
 					(reg_q618 AND symb_decoder(16#55#)) OR
 					(reg_q618 AND symb_decoder(16#73#)) OR
 					(reg_q618 AND symb_decoder(16#f3#)) OR
 					(reg_q618 AND symb_decoder(16#dc#)) OR
 					(reg_q618 AND symb_decoder(16#d9#)) OR
 					(reg_q618 AND symb_decoder(16#bb#)) OR
 					(reg_q618 AND symb_decoder(16#47#)) OR
 					(reg_q618 AND symb_decoder(16#ba#)) OR
 					(reg_q618 AND symb_decoder(16#14#)) OR
 					(reg_q618 AND symb_decoder(16#45#)) OR
 					(reg_q618 AND symb_decoder(16#b5#)) OR
 					(reg_q618 AND symb_decoder(16#03#)) OR
 					(reg_q618 AND symb_decoder(16#5d#)) OR
 					(reg_q618 AND symb_decoder(16#87#)) OR
 					(reg_q618 AND symb_decoder(16#c2#)) OR
 					(reg_q618 AND symb_decoder(16#2a#)) OR
 					(reg_q618 AND symb_decoder(16#dd#)) OR
 					(reg_q618 AND symb_decoder(16#bf#)) OR
 					(reg_q618 AND symb_decoder(16#fd#)) OR
 					(reg_q618 AND symb_decoder(16#c8#)) OR
 					(reg_q618 AND symb_decoder(16#07#)) OR
 					(reg_q618 AND symb_decoder(16#eb#)) OR
 					(reg_q618 AND symb_decoder(16#2f#)) OR
 					(reg_q618 AND symb_decoder(16#18#)) OR
 					(reg_q618 AND symb_decoder(16#97#)) OR
 					(reg_q618 AND symb_decoder(16#13#)) OR
 					(reg_q618 AND symb_decoder(16#58#)) OR
 					(reg_q618 AND symb_decoder(16#af#)) OR
 					(reg_q618 AND symb_decoder(16#9b#)) OR
 					(reg_q618 AND symb_decoder(16#28#)) OR
 					(reg_q618 AND symb_decoder(16#16#)) OR
 					(reg_q618 AND symb_decoder(16#e8#)) OR
 					(reg_q618 AND symb_decoder(16#cd#)) OR
 					(reg_q618 AND symb_decoder(16#54#)) OR
 					(reg_q618 AND symb_decoder(16#15#)) OR
 					(reg_q618 AND symb_decoder(16#65#)) OR
 					(reg_q618 AND symb_decoder(16#ca#)) OR
 					(reg_q618 AND symb_decoder(16#ae#)) OR
 					(reg_q618 AND symb_decoder(16#74#)) OR
 					(reg_q618 AND symb_decoder(16#3b#)) OR
 					(reg_q618 AND symb_decoder(16#40#)) OR
 					(reg_q618 AND symb_decoder(16#3f#)) OR
 					(reg_q618 AND symb_decoder(16#be#)) OR
 					(reg_q618 AND symb_decoder(16#6f#)) OR
 					(reg_q618 AND symb_decoder(16#12#)) OR
 					(reg_q618 AND symb_decoder(16#ab#)) OR
 					(reg_q618 AND symb_decoder(16#c4#)) OR
 					(reg_q618 AND symb_decoder(16#89#)) OR
 					(reg_q618 AND symb_decoder(16#31#)) OR
 					(reg_q618 AND symb_decoder(16#1f#)) OR
 					(reg_q618 AND symb_decoder(16#ed#)) OR
 					(reg_q618 AND symb_decoder(16#4c#)) OR
 					(reg_q618 AND symb_decoder(16#6b#)) OR
 					(reg_q618 AND symb_decoder(16#1c#)) OR
 					(reg_q618 AND symb_decoder(16#f2#)) OR
 					(reg_q618 AND symb_decoder(16#c9#)) OR
 					(reg_q618 AND symb_decoder(16#8c#)) OR
 					(reg_q618 AND symb_decoder(16#4d#)) OR
 					(reg_q618 AND symb_decoder(16#5e#)) OR
 					(reg_q618 AND symb_decoder(16#22#)) OR
 					(reg_q618 AND symb_decoder(16#e4#)) OR
 					(reg_q618 AND symb_decoder(16#60#)) OR
 					(reg_q618 AND symb_decoder(16#01#)) OR
 					(reg_q618 AND symb_decoder(16#c0#)) OR
 					(reg_q618 AND symb_decoder(16#b9#)) OR
 					(reg_q618 AND symb_decoder(16#83#)) OR
 					(reg_q618 AND symb_decoder(16#e6#)) OR
 					(reg_q618 AND symb_decoder(16#11#)) OR
 					(reg_q618 AND symb_decoder(16#04#)) OR
 					(reg_q618 AND symb_decoder(16#9f#)) OR
 					(reg_q618 AND symb_decoder(16#c6#)) OR
 					(reg_q618 AND symb_decoder(16#a4#)) OR
 					(reg_q618 AND symb_decoder(16#37#)) OR
 					(reg_q618 AND symb_decoder(16#de#)) OR
 					(reg_q618 AND symb_decoder(16#2d#)) OR
 					(reg_q618 AND symb_decoder(16#f4#)) OR
 					(reg_q618 AND symb_decoder(16#d4#)) OR
 					(reg_q618 AND symb_decoder(16#d2#)) OR
 					(reg_q618 AND symb_decoder(16#fb#)) OR
 					(reg_q618 AND symb_decoder(16#86#)) OR
 					(reg_q618 AND symb_decoder(16#39#)) OR
 					(reg_q618 AND symb_decoder(16#53#)) OR
 					(reg_q618 AND symb_decoder(16#94#)) OR
 					(reg_q618 AND symb_decoder(16#4f#)) OR
 					(reg_q618 AND symb_decoder(16#8b#)) OR
 					(reg_q618 AND symb_decoder(16#6a#)) OR
 					(reg_q618 AND symb_decoder(16#f6#)) OR
 					(reg_q618 AND symb_decoder(16#95#)) OR
 					(reg_q618 AND symb_decoder(16#cf#)) OR
 					(reg_q618 AND symb_decoder(16#57#)) OR
 					(reg_q618 AND symb_decoder(16#78#)) OR
 					(reg_q618 AND symb_decoder(16#98#)) OR
 					(reg_q618 AND symb_decoder(16#56#)) OR
 					(reg_q618 AND symb_decoder(16#e5#)) OR
 					(reg_q618 AND symb_decoder(16#a6#)) OR
 					(reg_q618 AND symb_decoder(16#32#)) OR
 					(reg_q618 AND symb_decoder(16#91#)) OR
 					(reg_q618 AND symb_decoder(16#10#)) OR
 					(reg_q618 AND symb_decoder(16#81#)) OR
 					(reg_q618 AND symb_decoder(16#7b#)) OR
 					(reg_q618 AND symb_decoder(16#d7#)) OR
 					(reg_q618 AND symb_decoder(16#19#)) OR
 					(reg_q618 AND symb_decoder(16#b0#)) OR
 					(reg_q618 AND symb_decoder(16#d8#)) OR
 					(reg_q618 AND symb_decoder(16#a7#)) OR
 					(reg_q618 AND symb_decoder(16#06#)) OR
 					(reg_q618 AND symb_decoder(16#fa#)) OR
 					(reg_q618 AND symb_decoder(16#30#)) OR
 					(reg_q618 AND symb_decoder(16#69#)) OR
 					(reg_q618 AND symb_decoder(16#c3#)) OR
 					(reg_q618 AND symb_decoder(16#85#)) OR
 					(reg_q618 AND symb_decoder(16#b4#)) OR
 					(reg_q618 AND symb_decoder(16#f8#)) OR
 					(reg_q618 AND symb_decoder(16#cc#)) OR
 					(reg_q618 AND symb_decoder(16#ad#)) OR
 					(reg_q618 AND symb_decoder(16#3a#)) OR
 					(reg_q618 AND symb_decoder(16#8a#)) OR
 					(reg_q618 AND symb_decoder(16#ea#)) OR
 					(reg_q618 AND symb_decoder(16#ec#)) OR
 					(reg_q618 AND symb_decoder(16#3d#)) OR
 					(reg_q618 AND symb_decoder(16#ac#)) OR
 					(reg_q618 AND symb_decoder(16#7c#)) OR
 					(reg_q618 AND symb_decoder(16#6d#)) OR
 					(reg_q618 AND symb_decoder(16#f7#)) OR
 					(reg_q618 AND symb_decoder(16#7d#)) OR
 					(reg_q618 AND symb_decoder(16#a1#)) OR
 					(reg_q618 AND symb_decoder(16#21#)) OR
 					(reg_q618 AND symb_decoder(16#1e#)) OR
 					(reg_q618 AND symb_decoder(16#a2#)) OR
 					(reg_q618 AND symb_decoder(16#96#)) OR
 					(reg_q618 AND symb_decoder(16#2b#)) OR
 					(reg_q618 AND symb_decoder(16#0e#)) OR
 					(reg_q618 AND symb_decoder(16#27#)) OR
 					(reg_q618 AND symb_decoder(16#f0#)) OR
 					(reg_q618 AND symb_decoder(16#9c#)) OR
 					(reg_q618 AND symb_decoder(16#9e#)) OR
 					(reg_q618 AND symb_decoder(16#a8#)) OR
 					(reg_q618 AND symb_decoder(16#42#)) OR
 					(reg_q618 AND symb_decoder(16#b2#)) OR
 					(reg_q618 AND symb_decoder(16#e1#)) OR
 					(reg_q618 AND symb_decoder(16#50#)) OR
 					(reg_q618 AND symb_decoder(16#cb#)) OR
 					(reg_q618 AND symb_decoder(16#67#)) OR
 					(reg_q618 AND symb_decoder(16#62#)) OR
 					(reg_q618 AND symb_decoder(16#4e#)) OR
 					(reg_q618 AND symb_decoder(16#c5#)) OR
 					(reg_q618 AND symb_decoder(16#bc#)) OR
 					(reg_q618 AND symb_decoder(16#b6#)) OR
 					(reg_q618 AND symb_decoder(16#33#)) OR
 					(reg_q618 AND symb_decoder(16#61#)) OR
 					(reg_q618 AND symb_decoder(16#64#)) OR
 					(reg_q618 AND symb_decoder(16#0f#)) OR
 					(reg_q618 AND symb_decoder(16#ef#)) OR
 					(reg_q618 AND symb_decoder(16#99#)) OR
 					(reg_q618 AND symb_decoder(16#82#)) OR
 					(reg_q618 AND symb_decoder(16#93#)) OR
 					(reg_q618 AND symb_decoder(16#8e#)) OR
 					(reg_q618 AND symb_decoder(16#b8#)) OR
 					(reg_q618 AND symb_decoder(16#f9#)) OR
 					(reg_q618 AND symb_decoder(16#a5#)) OR
 					(reg_q618 AND symb_decoder(16#41#)) OR
 					(reg_q618 AND symb_decoder(16#5b#)) OR
 					(reg_q618 AND symb_decoder(16#17#)) OR
 					(reg_q618 AND symb_decoder(16#0b#)) OR
 					(reg_q618 AND symb_decoder(16#38#)) OR
 					(reg_q618 AND symb_decoder(16#72#)) OR
 					(reg_q618 AND symb_decoder(16#c1#)) OR
 					(reg_q618 AND symb_decoder(16#26#)) OR
 					(reg_q618 AND symb_decoder(16#80#)) OR
 					(reg_q618 AND symb_decoder(16#2e#)) OR
 					(reg_q618 AND symb_decoder(16#2c#)) OR
 					(reg_q618 AND symb_decoder(16#1a#)) OR
 					(reg_q618 AND symb_decoder(16#9a#)) OR
 					(reg_q618 AND symb_decoder(16#e7#)) OR
 					(reg_q618 AND symb_decoder(16#d1#)) OR
 					(reg_q618 AND symb_decoder(16#a9#)) OR
 					(reg_q618 AND symb_decoder(16#c7#)) OR
 					(reg_q618 AND symb_decoder(16#f1#)) OR
 					(reg_q618 AND symb_decoder(16#84#)) OR
 					(reg_q618 AND symb_decoder(16#ee#)) OR
 					(reg_q618 AND symb_decoder(16#29#)) OR
 					(reg_q618 AND symb_decoder(16#90#)) OR
 					(reg_q618 AND symb_decoder(16#34#)) OR
 					(reg_q618 AND symb_decoder(16#79#)) OR
 					(reg_q618 AND symb_decoder(16#5c#)) OR
 					(reg_q618 AND symb_decoder(16#43#)) OR
 					(reg_q618 AND symb_decoder(16#a0#)) OR
 					(reg_q618 AND symb_decoder(16#76#)) OR
 					(reg_q618 AND symb_decoder(16#df#)) OR
 					(reg_q618 AND symb_decoder(16#63#)) OR
 					(reg_q618 AND symb_decoder(16#f5#)) OR
 					(reg_q618 AND symb_decoder(16#05#)) OR
 					(reg_q618 AND symb_decoder(16#db#)) OR
 					(reg_q618 AND symb_decoder(16#24#)) OR
 					(reg_q618 AND symb_decoder(16#9d#)) OR
 					(reg_q618 AND symb_decoder(16#d6#)) OR
 					(reg_q618 AND symb_decoder(16#00#)) OR
 					(reg_q618 AND symb_decoder(16#8f#)) OR
 					(reg_q618 AND symb_decoder(16#08#)) OR
 					(reg_q618 AND symb_decoder(16#aa#)) OR
 					(reg_q618 AND symb_decoder(16#23#)) OR
 					(reg_q618 AND symb_decoder(16#6e#)) OR
 					(reg_q618 AND symb_decoder(16#e3#)) OR
 					(reg_q618 AND symb_decoder(16#77#)) OR
 					(reg_q618 AND symb_decoder(16#7a#)) OR
 					(reg_q618 AND symb_decoder(16#66#)) OR
 					(reg_q618 AND symb_decoder(16#ce#)) OR
 					(reg_q618 AND symb_decoder(16#bd#)) OR
 					(reg_q618 AND symb_decoder(16#1b#)) OR
 					(reg_q618 AND symb_decoder(16#3e#)) OR
 					(reg_q618 AND symb_decoder(16#44#)) OR
 					(reg_q618 AND symb_decoder(16#7f#)) OR
 					(reg_q618 AND symb_decoder(16#88#)) OR
 					(reg_q618 AND symb_decoder(16#b3#)) OR
 					(reg_q618 AND symb_decoder(16#d5#)) OR
 					(reg_q618 AND symb_decoder(16#5a#)) OR
 					(reg_q618 AND symb_decoder(16#75#)) OR
 					(reg_q618 AND symb_decoder(16#1d#)) OR
 					(reg_q618 AND symb_decoder(16#7e#)) OR
 					(reg_q618 AND symb_decoder(16#d0#)) OR
 					(reg_q618 AND symb_decoder(16#ff#)) OR
 					(reg_q618 AND symb_decoder(16#52#)) OR
 					(reg_q618 AND symb_decoder(16#46#)) OR
 					(reg_q618 AND symb_decoder(16#3c#)) OR
 					(reg_q618 AND symb_decoder(16#8d#)) OR
 					(reg_q618 AND symb_decoder(16#b1#)) OR
 					(reg_q618 AND symb_decoder(16#92#)) OR
 					(reg_q618 AND symb_decoder(16#25#)) OR
 					(reg_q618 AND symb_decoder(16#35#)) OR
 					(reg_q618 AND symb_decoder(16#da#)) OR
 					(reg_q618 AND symb_decoder(16#a3#)) OR
 					(reg_q618 AND symb_decoder(16#4a#)) OR
 					(reg_q618 AND symb_decoder(16#49#));
reg_q48_in <= (reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q47 AND symb_decoder(16#30#));
reg_q227_in <= (reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q226 AND symb_decoder(16#36#));
reg_q229_in <= (reg_q227 AND symb_decoder(16#36#));
reg_q233_in <= (reg_q233 AND symb_decoder(16#31#)) OR
 					(reg_q233 AND symb_decoder(16#37#)) OR
 					(reg_q233 AND symb_decoder(16#33#)) OR
 					(reg_q233 AND symb_decoder(16#39#)) OR
 					(reg_q233 AND symb_decoder(16#32#)) OR
 					(reg_q233 AND symb_decoder(16#34#)) OR
 					(reg_q233 AND symb_decoder(16#36#)) OR
 					(reg_q233 AND symb_decoder(16#35#)) OR
 					(reg_q233 AND symb_decoder(16#30#)) OR
 					(reg_q233 AND symb_decoder(16#38#)) OR
 					(reg_q231 AND symb_decoder(16#34#)) OR
 					(reg_q231 AND symb_decoder(16#30#)) OR
 					(reg_q231 AND symb_decoder(16#33#)) OR
 					(reg_q231 AND symb_decoder(16#38#)) OR
 					(reg_q231 AND symb_decoder(16#39#)) OR
 					(reg_q231 AND symb_decoder(16#31#)) OR
 					(reg_q231 AND symb_decoder(16#36#)) OR
 					(reg_q231 AND symb_decoder(16#35#)) OR
 					(reg_q231 AND symb_decoder(16#32#)) OR
 					(reg_q231 AND symb_decoder(16#37#));
reg_q182_in <= (reg_q180 AND symb_decoder(16#30#));
reg_q184_in <= (reg_q182 AND symb_decoder(16#30#));
reg_q231_in <= (reg_q229 AND symb_decoder(16#36#));
reg_q1790_in <= (reg_q1788 AND symb_decoder(16#44#)) OR
 					(reg_q1788 AND symb_decoder(16#64#));
reg_q1385_in <= (reg_q1383 AND symb_decoder(16#6e#)) OR
 					(reg_q1383 AND symb_decoder(16#4e#));
reg_q1211_in <= (reg_q1209 AND symb_decoder(16#54#)) OR
 					(reg_q1209 AND symb_decoder(16#74#));
reg_q2451_in <= (reg_q2449 AND symb_decoder(16#32#));
reg_q2453_in <= (reg_q2451 AND symb_decoder(16#23#));
reg_q1015_in <= (reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q1014 AND symb_decoder(16#45#)) OR
 					(reg_q1014 AND symb_decoder(16#65#));
reg_q2128_in <= (reg_q2126 AND symb_decoder(16#45#)) OR
 					(reg_q2126 AND symb_decoder(16#65#));
reg_q2213_in <= (reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2212 AND symb_decoder(16#57#)) OR
 					(reg_q2212 AND symb_decoder(16#77#));
reg_q264_in <= (reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q263 AND symb_decoder(16#61#)) OR
 					(reg_q263 AND symb_decoder(16#41#));
reg_q705_in <= (reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q704 AND symb_decoder(16#63#)) OR
 					(reg_q704 AND symb_decoder(16#43#));
reg_q2132_in <= (reg_q2130 AND symb_decoder(16#47#)) OR
 					(reg_q2130 AND symb_decoder(16#67#));
reg_q1957_in <= (reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q1956 AND symb_decoder(16#53#)) OR
 					(reg_q1956 AND symb_decoder(16#73#));
reg_q2455_in <= (reg_q2453 AND symb_decoder(16#23#));
reg_q50_in <= (reg_q48 AND symb_decoder(16#30#));
reg_q52_in <= (reg_q50 AND symb_decoder(16#30#));
reg_q186_in <= (reg_q184 AND symb_decoder(16#30#));
reg_q1906_in <= (reg_q1904 AND symb_decoder(16#72#)) OR
 					(reg_q1904 AND symb_decoder(16#52#));
reg_q188_in <= (reg_q186 AND symb_decoder(16#31#));
reg_q190_in <= (reg_q188 AND symb_decoder(16#33#));
reg_q2068_in <= (reg_q2066 AND symb_decoder(16#46#));
reg_q2449_in <= (reg_q2447 AND symb_decoder(16#23#));
reg_q1377_in <= (reg_q1375 AND symb_decoder(16#49#)) OR
 					(reg_q1375 AND symb_decoder(16#69#));
reg_q180_in <= (reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q179 AND symb_decoder(16#31#));
reg_q416_in <= (reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q415 AND symb_decoder(16#42#)) OR
 					(reg_q415 AND symb_decoder(16#62#));
reg_q1694_in <= (reg_q1692 AND symb_decoder(16#47#)) OR
 					(reg_q1692 AND symb_decoder(16#67#));
reg_q718_in <= (reg_q716 AND symb_decoder(16#49#)) OR
 					(reg_q716 AND symb_decoder(16#69#));
reg_q2461_in <= (reg_q2459 AND symb_decoder(16#23#));
reg_q2070_in <= (reg_q2068 AND symb_decoder(16#54#));
reg_q2457_in <= (reg_q2455 AND symb_decoder(16#33#));
reg_q2459_in <= (reg_q2457 AND symb_decoder(16#23#));
reg_q2150_in <= (reg_q2148 AND symb_decoder(16#67#)) OR
 					(reg_q2148 AND symb_decoder(16#47#));
reg_q1375_in <= (reg_q1373 AND symb_decoder(16#46#)) OR
 					(reg_q1373 AND symb_decoder(16#66#));
reg_q97_in <= (reg_q95 AND symb_decoder(16#31#));
reg_q2465_in <= (reg_q2463 AND symb_decoder(16#23#));
reg_fullgraph43_init <= "000000";

reg_fullgraph43_sel <= "000000000000000000000" & reg_q2465_in & reg_q97_in & reg_q1375_in & reg_q2150_in & reg_q2459_in & reg_q2457_in & reg_q2070_in & reg_q2461_in & reg_q718_in & reg_q1694_in & reg_q416_in & reg_q180_in & reg_q1377_in & reg_q2449_in & reg_q2068_in & reg_q190_in & reg_q188_in & reg_q1906_in & reg_q186_in & reg_q52_in & reg_q50_in & reg_q2455_in & reg_q1957_in & reg_q2132_in & reg_q705_in & reg_q264_in & reg_q2213_in & reg_q2128_in & reg_q1015_in & reg_q2453_in & reg_q2451_in & reg_q1211_in & reg_q1385_in & reg_q1790_in & reg_q231_in & reg_q184_in & reg_q182_in & reg_q233_in & reg_q229_in & reg_q227_in & reg_q48_in & reg_q618_in & reg_q1772_in;

	--coder fullgraph43
with reg_fullgraph43_sel select
reg_fullgraph43_in <=
	"000001" when "0000000000000000000000000000000000000000000000000000000000000001",
	"000010" when "0000000000000000000000000000000000000000000000000000000000000010",
	"000011" when "0000000000000000000000000000000000000000000000000000000000000100",
	"000100" when "0000000000000000000000000000000000000000000000000000000000001000",
	"000101" when "0000000000000000000000000000000000000000000000000000000000010000",
	"000110" when "0000000000000000000000000000000000000000000000000000000000100000",
	"000111" when "0000000000000000000000000000000000000000000000000000000001000000",
	"001000" when "0000000000000000000000000000000000000000000000000000000010000000",
	"001001" when "0000000000000000000000000000000000000000000000000000000100000000",
	"001010" when "0000000000000000000000000000000000000000000000000000001000000000",
	"001011" when "0000000000000000000000000000000000000000000000000000010000000000",
	"001100" when "0000000000000000000000000000000000000000000000000000100000000000",
	"001101" when "0000000000000000000000000000000000000000000000000001000000000000",
	"001110" when "0000000000000000000000000000000000000000000000000010000000000000",
	"001111" when "0000000000000000000000000000000000000000000000000100000000000000",
	"010000" when "0000000000000000000000000000000000000000000000001000000000000000",
	"010001" when "0000000000000000000000000000000000000000000000010000000000000000",
	"010010" when "0000000000000000000000000000000000000000000000100000000000000000",
	"010011" when "0000000000000000000000000000000000000000000001000000000000000000",
	"010100" when "0000000000000000000000000000000000000000000010000000000000000000",
	"010101" when "0000000000000000000000000000000000000000000100000000000000000000",
	"010110" when "0000000000000000000000000000000000000000001000000000000000000000",
	"010111" when "0000000000000000000000000000000000000000010000000000000000000000",
	"011000" when "0000000000000000000000000000000000000000100000000000000000000000",
	"011001" when "0000000000000000000000000000000000000001000000000000000000000000",
	"011010" when "0000000000000000000000000000000000000010000000000000000000000000",
	"011011" when "0000000000000000000000000000000000000100000000000000000000000000",
	"011100" when "0000000000000000000000000000000000001000000000000000000000000000",
	"011101" when "0000000000000000000000000000000000010000000000000000000000000000",
	"011110" when "0000000000000000000000000000000000100000000000000000000000000000",
	"011111" when "0000000000000000000000000000000001000000000000000000000000000000",
	"100000" when "0000000000000000000000000000000010000000000000000000000000000000",
	"100001" when "0000000000000000000000000000000100000000000000000000000000000000",
	"100010" when "0000000000000000000000000000001000000000000000000000000000000000",
	"100011" when "0000000000000000000000000000010000000000000000000000000000000000",
	"100100" when "0000000000000000000000000000100000000000000000000000000000000000",
	"100101" when "0000000000000000000000000001000000000000000000000000000000000000",
	"100110" when "0000000000000000000000000010000000000000000000000000000000000000",
	"100111" when "0000000000000000000000000100000000000000000000000000000000000000",
	"101000" when "0000000000000000000000001000000000000000000000000000000000000000",
	"101001" when "0000000000000000000000010000000000000000000000000000000000000000",
	"101010" when "0000000000000000000000100000000000000000000000000000000000000000",
	"101011" when "0000000000000000000001000000000000000000000000000000000000000000",
	"000000" when others;
 --end coder

	p_reg_fullgraph43: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph43 <= reg_fullgraph43_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph43 <= reg_fullgraph43_init;
        else
          reg_fullgraph43 <= reg_fullgraph43_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph43

		reg_q1772 <= '1' when reg_fullgraph43 = "000001" else '0'; 
		reg_q618 <= '1' when reg_fullgraph43 = "000010" else '0'; 
		reg_q48 <= '1' when reg_fullgraph43 = "000011" else '0'; 
		reg_q227 <= '1' when reg_fullgraph43 = "000100" else '0'; 
		reg_q229 <= '1' when reg_fullgraph43 = "000101" else '0'; 
		reg_q233 <= '1' when reg_fullgraph43 = "000110" else '0'; 
		reg_q182 <= '1' when reg_fullgraph43 = "000111" else '0'; 
		reg_q184 <= '1' when reg_fullgraph43 = "001000" else '0'; 
		reg_q231 <= '1' when reg_fullgraph43 = "001001" else '0'; 
		reg_q1790 <= '1' when reg_fullgraph43 = "001010" else '0'; 
		reg_q1385 <= '1' when reg_fullgraph43 = "001011" else '0'; 
		reg_q1211 <= '1' when reg_fullgraph43 = "001100" else '0'; 
		reg_q2451 <= '1' when reg_fullgraph43 = "001101" else '0'; 
		reg_q2453 <= '1' when reg_fullgraph43 = "001110" else '0'; 
		reg_q1015 <= '1' when reg_fullgraph43 = "001111" else '0'; 
		reg_q2128 <= '1' when reg_fullgraph43 = "010000" else '0'; 
		reg_q2213 <= '1' when reg_fullgraph43 = "010001" else '0'; 
		reg_q264 <= '1' when reg_fullgraph43 = "010010" else '0'; 
		reg_q705 <= '1' when reg_fullgraph43 = "010011" else '0'; 
		reg_q2132 <= '1' when reg_fullgraph43 = "010100" else '0'; 
		reg_q1957 <= '1' when reg_fullgraph43 = "010101" else '0'; 
		reg_q2455 <= '1' when reg_fullgraph43 = "010110" else '0'; 
		reg_q50 <= '1' when reg_fullgraph43 = "010111" else '0'; 
		reg_q52 <= '1' when reg_fullgraph43 = "011000" else '0'; 
		reg_q186 <= '1' when reg_fullgraph43 = "011001" else '0'; 
		reg_q1906 <= '1' when reg_fullgraph43 = "011010" else '0'; 
		reg_q188 <= '1' when reg_fullgraph43 = "011011" else '0'; 
		reg_q190 <= '1' when reg_fullgraph43 = "011100" else '0'; 
		reg_q2068 <= '1' when reg_fullgraph43 = "011101" else '0'; 
		reg_q2449 <= '1' when reg_fullgraph43 = "011110" else '0'; 
		reg_q1377 <= '1' when reg_fullgraph43 = "011111" else '0'; 
		reg_q180 <= '1' when reg_fullgraph43 = "100000" else '0'; 
		reg_q416 <= '1' when reg_fullgraph43 = "100001" else '0'; 
		reg_q1694 <= '1' when reg_fullgraph43 = "100010" else '0'; 
		reg_q718 <= '1' when reg_fullgraph43 = "100011" else '0'; 
		reg_q2461 <= '1' when reg_fullgraph43 = "100100" else '0'; 
		reg_q2070 <= '1' when reg_fullgraph43 = "100101" else '0'; 
		reg_q2457 <= '1' when reg_fullgraph43 = "100110" else '0'; 
		reg_q2459 <= '1' when reg_fullgraph43 = "100111" else '0'; 
		reg_q2150 <= '1' when reg_fullgraph43 = "101000" else '0'; 
		reg_q1375 <= '1' when reg_fullgraph43 = "101001" else '0'; 
		reg_q97 <= '1' when reg_fullgraph43 = "101010" else '0'; 
		reg_q2465 <= '1' when reg_fullgraph43 = "101011" else '0'; 
--end decoder 

reg_q2211_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2211 AND symb_decoder(16#f3#)) OR
 					(reg_q2211 AND symb_decoder(16#7f#)) OR
 					(reg_q2211 AND symb_decoder(16#ac#)) OR
 					(reg_q2211 AND symb_decoder(16#01#)) OR
 					(reg_q2211 AND symb_decoder(16#a0#)) OR
 					(reg_q2211 AND symb_decoder(16#38#)) OR
 					(reg_q2211 AND symb_decoder(16#fb#)) OR
 					(reg_q2211 AND symb_decoder(16#83#)) OR
 					(reg_q2211 AND symb_decoder(16#b1#)) OR
 					(reg_q2211 AND symb_decoder(16#e7#)) OR
 					(reg_q2211 AND symb_decoder(16#fa#)) OR
 					(reg_q2211 AND symb_decoder(16#d6#)) OR
 					(reg_q2211 AND symb_decoder(16#9c#)) OR
 					(reg_q2211 AND symb_decoder(16#d2#)) OR
 					(reg_q2211 AND symb_decoder(16#ab#)) OR
 					(reg_q2211 AND symb_decoder(16#52#)) OR
 					(reg_q2211 AND symb_decoder(16#37#)) OR
 					(reg_q2211 AND symb_decoder(16#5a#)) OR
 					(reg_q2211 AND symb_decoder(16#42#)) OR
 					(reg_q2211 AND symb_decoder(16#e5#)) OR
 					(reg_q2211 AND symb_decoder(16#fd#)) OR
 					(reg_q2211 AND symb_decoder(16#49#)) OR
 					(reg_q2211 AND symb_decoder(16#1c#)) OR
 					(reg_q2211 AND symb_decoder(16#1d#)) OR
 					(reg_q2211 AND symb_decoder(16#04#)) OR
 					(reg_q2211 AND symb_decoder(16#7e#)) OR
 					(reg_q2211 AND symb_decoder(16#75#)) OR
 					(reg_q2211 AND symb_decoder(16#76#)) OR
 					(reg_q2211 AND symb_decoder(16#dc#)) OR
 					(reg_q2211 AND symb_decoder(16#46#)) OR
 					(reg_q2211 AND symb_decoder(16#5b#)) OR
 					(reg_q2211 AND symb_decoder(16#a2#)) OR
 					(reg_q2211 AND symb_decoder(16#89#)) OR
 					(reg_q2211 AND symb_decoder(16#64#)) OR
 					(reg_q2211 AND symb_decoder(16#43#)) OR
 					(reg_q2211 AND symb_decoder(16#e3#)) OR
 					(reg_q2211 AND symb_decoder(16#06#)) OR
 					(reg_q2211 AND symb_decoder(16#1f#)) OR
 					(reg_q2211 AND symb_decoder(16#47#)) OR
 					(reg_q2211 AND symb_decoder(16#af#)) OR
 					(reg_q2211 AND symb_decoder(16#2a#)) OR
 					(reg_q2211 AND symb_decoder(16#26#)) OR
 					(reg_q2211 AND symb_decoder(16#a3#)) OR
 					(reg_q2211 AND symb_decoder(16#72#)) OR
 					(reg_q2211 AND symb_decoder(16#71#)) OR
 					(reg_q2211 AND symb_decoder(16#32#)) OR
 					(reg_q2211 AND symb_decoder(16#ae#)) OR
 					(reg_q2211 AND symb_decoder(16#fe#)) OR
 					(reg_q2211 AND symb_decoder(16#4b#)) OR
 					(reg_q2211 AND symb_decoder(16#4f#)) OR
 					(reg_q2211 AND symb_decoder(16#e6#)) OR
 					(reg_q2211 AND symb_decoder(16#4d#)) OR
 					(reg_q2211 AND symb_decoder(16#c9#)) OR
 					(reg_q2211 AND symb_decoder(16#4a#)) OR
 					(reg_q2211 AND symb_decoder(16#c7#)) OR
 					(reg_q2211 AND symb_decoder(16#a8#)) OR
 					(reg_q2211 AND symb_decoder(16#81#)) OR
 					(reg_q2211 AND symb_decoder(16#c0#)) OR
 					(reg_q2211 AND symb_decoder(16#2c#)) OR
 					(reg_q2211 AND symb_decoder(16#07#)) OR
 					(reg_q2211 AND symb_decoder(16#60#)) OR
 					(reg_q2211 AND symb_decoder(16#15#)) OR
 					(reg_q2211 AND symb_decoder(16#70#)) OR
 					(reg_q2211 AND symb_decoder(16#78#)) OR
 					(reg_q2211 AND symb_decoder(16#ec#)) OR
 					(reg_q2211 AND symb_decoder(16#51#)) OR
 					(reg_q2211 AND symb_decoder(16#f7#)) OR
 					(reg_q2211 AND symb_decoder(16#9f#)) OR
 					(reg_q2211 AND symb_decoder(16#b7#)) OR
 					(reg_q2211 AND symb_decoder(16#ce#)) OR
 					(reg_q2211 AND symb_decoder(16#69#)) OR
 					(reg_q2211 AND symb_decoder(16#21#)) OR
 					(reg_q2211 AND symb_decoder(16#00#)) OR
 					(reg_q2211 AND symb_decoder(16#92#)) OR
 					(reg_q2211 AND symb_decoder(16#b9#)) OR
 					(reg_q2211 AND symb_decoder(16#4e#)) OR
 					(reg_q2211 AND symb_decoder(16#bc#)) OR
 					(reg_q2211 AND symb_decoder(16#1b#)) OR
 					(reg_q2211 AND symb_decoder(16#bf#)) OR
 					(reg_q2211 AND symb_decoder(16#9d#)) OR
 					(reg_q2211 AND symb_decoder(16#6d#)) OR
 					(reg_q2211 AND symb_decoder(16#c5#)) OR
 					(reg_q2211 AND symb_decoder(16#18#)) OR
 					(reg_q2211 AND symb_decoder(16#99#)) OR
 					(reg_q2211 AND symb_decoder(16#84#)) OR
 					(reg_q2211 AND symb_decoder(16#2e#)) OR
 					(reg_q2211 AND symb_decoder(16#5f#)) OR
 					(reg_q2211 AND symb_decoder(16#8a#)) OR
 					(reg_q2211 AND symb_decoder(16#80#)) OR
 					(reg_q2211 AND symb_decoder(16#ee#)) OR
 					(reg_q2211 AND symb_decoder(16#0d#)) OR
 					(reg_q2211 AND symb_decoder(16#d7#)) OR
 					(reg_q2211 AND symb_decoder(16#23#)) OR
 					(reg_q2211 AND symb_decoder(16#e1#)) OR
 					(reg_q2211 AND symb_decoder(16#30#)) OR
 					(reg_q2211 AND symb_decoder(16#7b#)) OR
 					(reg_q2211 AND symb_decoder(16#96#)) OR
 					(reg_q2211 AND symb_decoder(16#b8#)) OR
 					(reg_q2211 AND symb_decoder(16#53#)) OR
 					(reg_q2211 AND symb_decoder(16#0f#)) OR
 					(reg_q2211 AND symb_decoder(16#8b#)) OR
 					(reg_q2211 AND symb_decoder(16#35#)) OR
 					(reg_q2211 AND symb_decoder(16#6b#)) OR
 					(reg_q2211 AND symb_decoder(16#16#)) OR
 					(reg_q2211 AND symb_decoder(16#20#)) OR
 					(reg_q2211 AND symb_decoder(16#2f#)) OR
 					(reg_q2211 AND symb_decoder(16#9e#)) OR
 					(reg_q2211 AND symb_decoder(16#df#)) OR
 					(reg_q2211 AND symb_decoder(16#8c#)) OR
 					(reg_q2211 AND symb_decoder(16#41#)) OR
 					(reg_q2211 AND symb_decoder(16#82#)) OR
 					(reg_q2211 AND symb_decoder(16#19#)) OR
 					(reg_q2211 AND symb_decoder(16#f4#)) OR
 					(reg_q2211 AND symb_decoder(16#f8#)) OR
 					(reg_q2211 AND symb_decoder(16#f1#)) OR
 					(reg_q2211 AND symb_decoder(16#40#)) OR
 					(reg_q2211 AND symb_decoder(16#3a#)) OR
 					(reg_q2211 AND symb_decoder(16#f2#)) OR
 					(reg_q2211 AND symb_decoder(16#0a#)) OR
 					(reg_q2211 AND symb_decoder(16#f0#)) OR
 					(reg_q2211 AND symb_decoder(16#57#)) OR
 					(reg_q2211 AND symb_decoder(16#4c#)) OR
 					(reg_q2211 AND symb_decoder(16#db#)) OR
 					(reg_q2211 AND symb_decoder(16#6e#)) OR
 					(reg_q2211 AND symb_decoder(16#6f#)) OR
 					(reg_q2211 AND symb_decoder(16#08#)) OR
 					(reg_q2211 AND symb_decoder(16#10#)) OR
 					(reg_q2211 AND symb_decoder(16#59#)) OR
 					(reg_q2211 AND symb_decoder(16#9a#)) OR
 					(reg_q2211 AND symb_decoder(16#09#)) OR
 					(reg_q2211 AND symb_decoder(16#a9#)) OR
 					(reg_q2211 AND symb_decoder(16#3c#)) OR
 					(reg_q2211 AND symb_decoder(16#33#)) OR
 					(reg_q2211 AND symb_decoder(16#d4#)) OR
 					(reg_q2211 AND symb_decoder(16#50#)) OR
 					(reg_q2211 AND symb_decoder(16#93#)) OR
 					(reg_q2211 AND symb_decoder(16#d3#)) OR
 					(reg_q2211 AND symb_decoder(16#14#)) OR
 					(reg_q2211 AND symb_decoder(16#8f#)) OR
 					(reg_q2211 AND symb_decoder(16#7a#)) OR
 					(reg_q2211 AND symb_decoder(16#17#)) OR
 					(reg_q2211 AND symb_decoder(16#b5#)) OR
 					(reg_q2211 AND symb_decoder(16#ea#)) OR
 					(reg_q2211 AND symb_decoder(16#ed#)) OR
 					(reg_q2211 AND symb_decoder(16#c4#)) OR
 					(reg_q2211 AND symb_decoder(16#cb#)) OR
 					(reg_q2211 AND symb_decoder(16#a5#)) OR
 					(reg_q2211 AND symb_decoder(16#d8#)) OR
 					(reg_q2211 AND symb_decoder(16#90#)) OR
 					(reg_q2211 AND symb_decoder(16#11#)) OR
 					(reg_q2211 AND symb_decoder(16#b4#)) OR
 					(reg_q2211 AND symb_decoder(16#9b#)) OR
 					(reg_q2211 AND symb_decoder(16#d0#)) OR
 					(reg_q2211 AND symb_decoder(16#f9#)) OR
 					(reg_q2211 AND symb_decoder(16#27#)) OR
 					(reg_q2211 AND symb_decoder(16#d5#)) OR
 					(reg_q2211 AND symb_decoder(16#91#)) OR
 					(reg_q2211 AND symb_decoder(16#48#)) OR
 					(reg_q2211 AND symb_decoder(16#ad#)) OR
 					(reg_q2211 AND symb_decoder(16#65#)) OR
 					(reg_q2211 AND symb_decoder(16#c1#)) OR
 					(reg_q2211 AND symb_decoder(16#0e#)) OR
 					(reg_q2211 AND symb_decoder(16#44#)) OR
 					(reg_q2211 AND symb_decoder(16#e4#)) OR
 					(reg_q2211 AND symb_decoder(16#3f#)) OR
 					(reg_q2211 AND symb_decoder(16#77#)) OR
 					(reg_q2211 AND symb_decoder(16#66#)) OR
 					(reg_q2211 AND symb_decoder(16#8d#)) OR
 					(reg_q2211 AND symb_decoder(16#1e#)) OR
 					(reg_q2211 AND symb_decoder(16#3e#)) OR
 					(reg_q2211 AND symb_decoder(16#a4#)) OR
 					(reg_q2211 AND symb_decoder(16#2d#)) OR
 					(reg_q2211 AND symb_decoder(16#36#)) OR
 					(reg_q2211 AND symb_decoder(16#94#)) OR
 					(reg_q2211 AND symb_decoder(16#79#)) OR
 					(reg_q2211 AND symb_decoder(16#aa#)) OR
 					(reg_q2211 AND symb_decoder(16#f6#)) OR
 					(reg_q2211 AND symb_decoder(16#25#)) OR
 					(reg_q2211 AND symb_decoder(16#68#)) OR
 					(reg_q2211 AND symb_decoder(16#c2#)) OR
 					(reg_q2211 AND symb_decoder(16#be#)) OR
 					(reg_q2211 AND symb_decoder(16#5c#)) OR
 					(reg_q2211 AND symb_decoder(16#b3#)) OR
 					(reg_q2211 AND symb_decoder(16#0c#)) OR
 					(reg_q2211 AND symb_decoder(16#fc#)) OR
 					(reg_q2211 AND symb_decoder(16#ba#)) OR
 					(reg_q2211 AND symb_decoder(16#dd#)) OR
 					(reg_q2211 AND symb_decoder(16#12#)) OR
 					(reg_q2211 AND symb_decoder(16#97#)) OR
 					(reg_q2211 AND symb_decoder(16#c8#)) OR
 					(reg_q2211 AND symb_decoder(16#eb#)) OR
 					(reg_q2211 AND symb_decoder(16#29#)) OR
 					(reg_q2211 AND symb_decoder(16#ff#)) OR
 					(reg_q2211 AND symb_decoder(16#ef#)) OR
 					(reg_q2211 AND symb_decoder(16#45#)) OR
 					(reg_q2211 AND symb_decoder(16#39#)) OR
 					(reg_q2211 AND symb_decoder(16#b2#)) OR
 					(reg_q2211 AND symb_decoder(16#7c#)) OR
 					(reg_q2211 AND symb_decoder(16#e0#)) OR
 					(reg_q2211 AND symb_decoder(16#74#)) OR
 					(reg_q2211 AND symb_decoder(16#13#)) OR
 					(reg_q2211 AND symb_decoder(16#3b#)) OR
 					(reg_q2211 AND symb_decoder(16#cc#)) OR
 					(reg_q2211 AND symb_decoder(16#22#)) OR
 					(reg_q2211 AND symb_decoder(16#0b#)) OR
 					(reg_q2211 AND symb_decoder(16#a7#)) OR
 					(reg_q2211 AND symb_decoder(16#a6#)) OR
 					(reg_q2211 AND symb_decoder(16#62#)) OR
 					(reg_q2211 AND symb_decoder(16#87#)) OR
 					(reg_q2211 AND symb_decoder(16#d9#)) OR
 					(reg_q2211 AND symb_decoder(16#56#)) OR
 					(reg_q2211 AND symb_decoder(16#c6#)) OR
 					(reg_q2211 AND symb_decoder(16#02#)) OR
 					(reg_q2211 AND symb_decoder(16#ca#)) OR
 					(reg_q2211 AND symb_decoder(16#d1#)) OR
 					(reg_q2211 AND symb_decoder(16#34#)) OR
 					(reg_q2211 AND symb_decoder(16#bb#)) OR
 					(reg_q2211 AND symb_decoder(16#85#)) OR
 					(reg_q2211 AND symb_decoder(16#e8#)) OR
 					(reg_q2211 AND symb_decoder(16#2b#)) OR
 					(reg_q2211 AND symb_decoder(16#de#)) OR
 					(reg_q2211 AND symb_decoder(16#f5#)) OR
 					(reg_q2211 AND symb_decoder(16#55#)) OR
 					(reg_q2211 AND symb_decoder(16#3d#)) OR
 					(reg_q2211 AND symb_decoder(16#31#)) OR
 					(reg_q2211 AND symb_decoder(16#95#)) OR
 					(reg_q2211 AND symb_decoder(16#5d#)) OR
 					(reg_q2211 AND symb_decoder(16#28#)) OR
 					(reg_q2211 AND symb_decoder(16#b0#)) OR
 					(reg_q2211 AND symb_decoder(16#98#)) OR
 					(reg_q2211 AND symb_decoder(16#86#)) OR
 					(reg_q2211 AND symb_decoder(16#63#)) OR
 					(reg_q2211 AND symb_decoder(16#8e#)) OR
 					(reg_q2211 AND symb_decoder(16#cf#)) OR
 					(reg_q2211 AND symb_decoder(16#05#)) OR
 					(reg_q2211 AND symb_decoder(16#24#)) OR
 					(reg_q2211 AND symb_decoder(16#c3#)) OR
 					(reg_q2211 AND symb_decoder(16#67#)) OR
 					(reg_q2211 AND symb_decoder(16#5e#)) OR
 					(reg_q2211 AND symb_decoder(16#73#)) OR
 					(reg_q2211 AND symb_decoder(16#7d#)) OR
 					(reg_q2211 AND symb_decoder(16#a1#)) OR
 					(reg_q2211 AND symb_decoder(16#61#)) OR
 					(reg_q2211 AND symb_decoder(16#da#)) OR
 					(reg_q2211 AND symb_decoder(16#b6#)) OR
 					(reg_q2211 AND symb_decoder(16#6a#)) OR
 					(reg_q2211 AND symb_decoder(16#bd#)) OR
 					(reg_q2211 AND symb_decoder(16#58#)) OR
 					(reg_q2211 AND symb_decoder(16#03#)) OR
 					(reg_q2211 AND symb_decoder(16#6c#)) OR
 					(reg_q2211 AND symb_decoder(16#88#)) OR
 					(reg_q2211 AND symb_decoder(16#e9#)) OR
 					(reg_q2211 AND symb_decoder(16#e2#)) OR
 					(reg_q2211 AND symb_decoder(16#1a#)) OR
 					(reg_q2211 AND symb_decoder(16#cd#)) OR
 					(reg_q2211 AND symb_decoder(16#54#));
reg_q2211_init <= '0' ;
	p_reg_q2211: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2211 <= reg_q2211_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2211 <= reg_q2211_init;
        else
          reg_q2211 <= reg_q2211_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph45

reg_q813_in <= (reg_q813 AND symb_decoder(16#47#)) OR
 					(reg_q813 AND symb_decoder(16#87#)) OR
 					(reg_q813 AND symb_decoder(16#d6#)) OR
 					(reg_q813 AND symb_decoder(16#7e#)) OR
 					(reg_q813 AND symb_decoder(16#dd#)) OR
 					(reg_q813 AND symb_decoder(16#ce#)) OR
 					(reg_q813 AND symb_decoder(16#ea#)) OR
 					(reg_q813 AND symb_decoder(16#2d#)) OR
 					(reg_q813 AND symb_decoder(16#f2#)) OR
 					(reg_q813 AND symb_decoder(16#62#)) OR
 					(reg_q813 AND symb_decoder(16#37#)) OR
 					(reg_q813 AND symb_decoder(16#8c#)) OR
 					(reg_q813 AND symb_decoder(16#2e#)) OR
 					(reg_q813 AND symb_decoder(16#75#)) OR
 					(reg_q813 AND symb_decoder(16#1c#)) OR
 					(reg_q813 AND symb_decoder(16#f4#)) OR
 					(reg_q813 AND symb_decoder(16#d7#)) OR
 					(reg_q813 AND symb_decoder(16#bb#)) OR
 					(reg_q813 AND symb_decoder(16#2b#)) OR
 					(reg_q813 AND symb_decoder(16#a5#)) OR
 					(reg_q813 AND symb_decoder(16#ab#)) OR
 					(reg_q813 AND symb_decoder(16#94#)) OR
 					(reg_q813 AND symb_decoder(16#dc#)) OR
 					(reg_q813 AND symb_decoder(16#71#)) OR
 					(reg_q813 AND symb_decoder(16#cc#)) OR
 					(reg_q813 AND symb_decoder(16#04#)) OR
 					(reg_q813 AND symb_decoder(16#6e#)) OR
 					(reg_q813 AND symb_decoder(16#43#)) OR
 					(reg_q813 AND symb_decoder(16#b9#)) OR
 					(reg_q813 AND symb_decoder(16#e8#)) OR
 					(reg_q813 AND symb_decoder(16#d8#)) OR
 					(reg_q813 AND symb_decoder(16#6c#)) OR
 					(reg_q813 AND symb_decoder(16#9c#)) OR
 					(reg_q813 AND symb_decoder(16#e0#)) OR
 					(reg_q813 AND symb_decoder(16#44#)) OR
 					(reg_q813 AND symb_decoder(16#66#)) OR
 					(reg_q813 AND symb_decoder(16#bc#)) OR
 					(reg_q813 AND symb_decoder(16#17#)) OR
 					(reg_q813 AND symb_decoder(16#3e#)) OR
 					(reg_q813 AND symb_decoder(16#ff#)) OR
 					(reg_q813 AND symb_decoder(16#b7#)) OR
 					(reg_q813 AND symb_decoder(16#3d#)) OR
 					(reg_q813 AND symb_decoder(16#5f#)) OR
 					(reg_q813 AND symb_decoder(16#84#)) OR
 					(reg_q813 AND symb_decoder(16#39#)) OR
 					(reg_q813 AND symb_decoder(16#01#)) OR
 					(reg_q813 AND symb_decoder(16#82#)) OR
 					(reg_q813 AND symb_decoder(16#a6#)) OR
 					(reg_q813 AND symb_decoder(16#68#)) OR
 					(reg_q813 AND symb_decoder(16#59#)) OR
 					(reg_q813 AND symb_decoder(16#f1#)) OR
 					(reg_q813 AND symb_decoder(16#2f#)) OR
 					(reg_q813 AND symb_decoder(16#35#)) OR
 					(reg_q813 AND symb_decoder(16#3a#)) OR
 					(reg_q813 AND symb_decoder(16#7b#)) OR
 					(reg_q813 AND symb_decoder(16#8e#)) OR
 					(reg_q813 AND symb_decoder(16#15#)) OR
 					(reg_q813 AND symb_decoder(16#65#)) OR
 					(reg_q813 AND symb_decoder(16#fc#)) OR
 					(reg_q813 AND symb_decoder(16#6f#)) OR
 					(reg_q813 AND symb_decoder(16#03#)) OR
 					(reg_q813 AND symb_decoder(16#e3#)) OR
 					(reg_q813 AND symb_decoder(16#9b#)) OR
 					(reg_q813 AND symb_decoder(16#0c#)) OR
 					(reg_q813 AND symb_decoder(16#88#)) OR
 					(reg_q813 AND symb_decoder(16#f3#)) OR
 					(reg_q813 AND symb_decoder(16#c4#)) OR
 					(reg_q813 AND symb_decoder(16#45#)) OR
 					(reg_q813 AND symb_decoder(16#b3#)) OR
 					(reg_q813 AND symb_decoder(16#c0#)) OR
 					(reg_q813 AND symb_decoder(16#51#)) OR
 					(reg_q813 AND symb_decoder(16#fe#)) OR
 					(reg_q813 AND symb_decoder(16#a8#)) OR
 					(reg_q813 AND symb_decoder(16#61#)) OR
 					(reg_q813 AND symb_decoder(16#18#)) OR
 					(reg_q813 AND symb_decoder(16#14#)) OR
 					(reg_q813 AND symb_decoder(16#73#)) OR
 					(reg_q813 AND symb_decoder(16#aa#)) OR
 					(reg_q813 AND symb_decoder(16#ba#)) OR
 					(reg_q813 AND symb_decoder(16#09#)) OR
 					(reg_q813 AND symb_decoder(16#0f#)) OR
 					(reg_q813 AND symb_decoder(16#8b#)) OR
 					(reg_q813 AND symb_decoder(16#80#)) OR
 					(reg_q813 AND symb_decoder(16#77#)) OR
 					(reg_q813 AND symb_decoder(16#f5#)) OR
 					(reg_q813 AND symb_decoder(16#49#)) OR
 					(reg_q813 AND symb_decoder(16#d4#)) OR
 					(reg_q813 AND symb_decoder(16#b0#)) OR
 					(reg_q813 AND symb_decoder(16#cb#)) OR
 					(reg_q813 AND symb_decoder(16#a1#)) OR
 					(reg_q813 AND symb_decoder(16#1a#)) OR
 					(reg_q813 AND symb_decoder(16#f9#)) OR
 					(reg_q813 AND symb_decoder(16#60#)) OR
 					(reg_q813 AND symb_decoder(16#c9#)) OR
 					(reg_q813 AND symb_decoder(16#90#)) OR
 					(reg_q813 AND symb_decoder(16#5e#)) OR
 					(reg_q813 AND symb_decoder(16#7a#)) OR
 					(reg_q813 AND symb_decoder(16#f7#)) OR
 					(reg_q813 AND symb_decoder(16#5b#)) OR
 					(reg_q813 AND symb_decoder(16#a3#)) OR
 					(reg_q813 AND symb_decoder(16#67#)) OR
 					(reg_q813 AND symb_decoder(16#40#)) OR
 					(reg_q813 AND symb_decoder(16#e1#)) OR
 					(reg_q813 AND symb_decoder(16#23#)) OR
 					(reg_q813 AND symb_decoder(16#48#)) OR
 					(reg_q813 AND symb_decoder(16#da#)) OR
 					(reg_q813 AND symb_decoder(16#b4#)) OR
 					(reg_q813 AND symb_decoder(16#d0#)) OR
 					(reg_q813 AND symb_decoder(16#56#)) OR
 					(reg_q813 AND symb_decoder(16#22#)) OR
 					(reg_q813 AND symb_decoder(16#85#)) OR
 					(reg_q813 AND symb_decoder(16#cd#)) OR
 					(reg_q813 AND symb_decoder(16#54#)) OR
 					(reg_q813 AND symb_decoder(16#c5#)) OR
 					(reg_q813 AND symb_decoder(16#b2#)) OR
 					(reg_q813 AND symb_decoder(16#d5#)) OR
 					(reg_q813 AND symb_decoder(16#c7#)) OR
 					(reg_q813 AND symb_decoder(16#3c#)) OR
 					(reg_q813 AND symb_decoder(16#ef#)) OR
 					(reg_q813 AND symb_decoder(16#21#)) OR
 					(reg_q813 AND symb_decoder(16#a9#)) OR
 					(reg_q813 AND symb_decoder(16#a4#)) OR
 					(reg_q813 AND symb_decoder(16#b8#)) OR
 					(reg_q813 AND symb_decoder(16#31#)) OR
 					(reg_q813 AND symb_decoder(16#36#)) OR
 					(reg_q813 AND symb_decoder(16#41#)) OR
 					(reg_q813 AND symb_decoder(16#fd#)) OR
 					(reg_q813 AND symb_decoder(16#5a#)) OR
 					(reg_q813 AND symb_decoder(16#0e#)) OR
 					(reg_q813 AND symb_decoder(16#be#)) OR
 					(reg_q813 AND symb_decoder(16#a0#)) OR
 					(reg_q813 AND symb_decoder(16#30#)) OR
 					(reg_q813 AND symb_decoder(16#08#)) OR
 					(reg_q813 AND symb_decoder(16#fa#)) OR
 					(reg_q813 AND symb_decoder(16#11#)) OR
 					(reg_q813 AND symb_decoder(16#91#)) OR
 					(reg_q813 AND symb_decoder(16#72#)) OR
 					(reg_q813 AND symb_decoder(16#7d#)) OR
 					(reg_q813 AND symb_decoder(16#ae#)) OR
 					(reg_q813 AND symb_decoder(16#02#)) OR
 					(reg_q813 AND symb_decoder(16#7c#)) OR
 					(reg_q813 AND symb_decoder(16#db#)) OR
 					(reg_q813 AND symb_decoder(16#53#)) OR
 					(reg_q813 AND symb_decoder(16#f8#)) OR
 					(reg_q813 AND symb_decoder(16#de#)) OR
 					(reg_q813 AND symb_decoder(16#a2#)) OR
 					(reg_q813 AND symb_decoder(16#16#)) OR
 					(reg_q813 AND symb_decoder(16#d1#)) OR
 					(reg_q813 AND symb_decoder(16#8d#)) OR
 					(reg_q813 AND symb_decoder(16#ed#)) OR
 					(reg_q813 AND symb_decoder(16#57#)) OR
 					(reg_q813 AND symb_decoder(16#70#)) OR
 					(reg_q813 AND symb_decoder(16#46#)) OR
 					(reg_q813 AND symb_decoder(16#69#)) OR
 					(reg_q813 AND symb_decoder(16#e5#)) OR
 					(reg_q813 AND symb_decoder(16#e6#)) OR
 					(reg_q813 AND symb_decoder(16#c2#)) OR
 					(reg_q813 AND symb_decoder(16#4b#)) OR
 					(reg_q813 AND symb_decoder(16#55#)) OR
 					(reg_q813 AND symb_decoder(16#bd#)) OR
 					(reg_q813 AND symb_decoder(16#df#)) OR
 					(reg_q813 AND symb_decoder(16#07#)) OR
 					(reg_q813 AND symb_decoder(16#8a#)) OR
 					(reg_q813 AND symb_decoder(16#9d#)) OR
 					(reg_q813 AND symb_decoder(16#83#)) OR
 					(reg_q813 AND symb_decoder(16#ad#)) OR
 					(reg_q813 AND symb_decoder(16#05#)) OR
 					(reg_q813 AND symb_decoder(16#06#)) OR
 					(reg_q813 AND symb_decoder(16#a7#)) OR
 					(reg_q813 AND symb_decoder(16#ca#)) OR
 					(reg_q813 AND symb_decoder(16#1d#)) OR
 					(reg_q813 AND symb_decoder(16#27#)) OR
 					(reg_q813 AND symb_decoder(16#0b#)) OR
 					(reg_q813 AND symb_decoder(16#9a#)) OR
 					(reg_q813 AND symb_decoder(16#5d#)) OR
 					(reg_q813 AND symb_decoder(16#92#)) OR
 					(reg_q813 AND symb_decoder(16#e2#)) OR
 					(reg_q813 AND symb_decoder(16#6b#)) OR
 					(reg_q813 AND symb_decoder(16#c3#)) OR
 					(reg_q813 AND symb_decoder(16#33#)) OR
 					(reg_q813 AND symb_decoder(16#6d#)) OR
 					(reg_q813 AND symb_decoder(16#13#)) OR
 					(reg_q813 AND symb_decoder(16#34#)) OR
 					(reg_q813 AND symb_decoder(16#2a#)) OR
 					(reg_q813 AND symb_decoder(16#95#)) OR
 					(reg_q813 AND symb_decoder(16#1e#)) OR
 					(reg_q813 AND symb_decoder(16#4a#)) OR
 					(reg_q813 AND symb_decoder(16#52#)) OR
 					(reg_q813 AND symb_decoder(16#3f#)) OR
 					(reg_q813 AND symb_decoder(16#00#)) OR
 					(reg_q813 AND symb_decoder(16#50#)) OR
 					(reg_q813 AND symb_decoder(16#2c#)) OR
 					(reg_q813 AND symb_decoder(16#ec#)) OR
 					(reg_q813 AND symb_decoder(16#86#)) OR
 					(reg_q813 AND symb_decoder(16#64#)) OR
 					(reg_q813 AND symb_decoder(16#ac#)) OR
 					(reg_q813 AND symb_decoder(16#4f#)) OR
 					(reg_q813 AND symb_decoder(16#fb#)) OR
 					(reg_q813 AND symb_decoder(16#4c#)) OR
 					(reg_q813 AND symb_decoder(16#ee#)) OR
 					(reg_q813 AND symb_decoder(16#5c#)) OR
 					(reg_q813 AND symb_decoder(16#99#)) OR
 					(reg_q813 AND symb_decoder(16#79#)) OR
 					(reg_q813 AND symb_decoder(16#c1#)) OR
 					(reg_q813 AND symb_decoder(16#20#)) OR
 					(reg_q813 AND symb_decoder(16#96#)) OR
 					(reg_q813 AND symb_decoder(16#d3#)) OR
 					(reg_q813 AND symb_decoder(16#98#)) OR
 					(reg_q813 AND symb_decoder(16#78#)) OR
 					(reg_q813 AND symb_decoder(16#e9#)) OR
 					(reg_q813 AND symb_decoder(16#eb#)) OR
 					(reg_q813 AND symb_decoder(16#6a#)) OR
 					(reg_q813 AND symb_decoder(16#19#)) OR
 					(reg_q813 AND symb_decoder(16#81#)) OR
 					(reg_q813 AND symb_decoder(16#63#)) OR
 					(reg_q813 AND symb_decoder(16#c8#)) OR
 					(reg_q813 AND symb_decoder(16#9e#)) OR
 					(reg_q813 AND symb_decoder(16#e7#)) OR
 					(reg_q813 AND symb_decoder(16#26#)) OR
 					(reg_q813 AND symb_decoder(16#28#)) OR
 					(reg_q813 AND symb_decoder(16#8f#)) OR
 					(reg_q813 AND symb_decoder(16#74#)) OR
 					(reg_q813 AND symb_decoder(16#b6#)) OR
 					(reg_q813 AND symb_decoder(16#93#)) OR
 					(reg_q813 AND symb_decoder(16#10#)) OR
 					(reg_q813 AND symb_decoder(16#58#)) OR
 					(reg_q813 AND symb_decoder(16#38#)) OR
 					(reg_q813 AND symb_decoder(16#b1#)) OR
 					(reg_q813 AND symb_decoder(16#bf#)) OR
 					(reg_q813 AND symb_decoder(16#9f#)) OR
 					(reg_q813 AND symb_decoder(16#1b#)) OR
 					(reg_q813 AND symb_decoder(16#cf#)) OR
 					(reg_q813 AND symb_decoder(16#12#)) OR
 					(reg_q813 AND symb_decoder(16#25#)) OR
 					(reg_q813 AND symb_decoder(16#f0#)) OR
 					(reg_q813 AND symb_decoder(16#7f#)) OR
 					(reg_q813 AND symb_decoder(16#42#)) OR
 					(reg_q813 AND symb_decoder(16#4d#)) OR
 					(reg_q813 AND symb_decoder(16#97#)) OR
 					(reg_q813 AND symb_decoder(16#af#)) OR
 					(reg_q813 AND symb_decoder(16#e4#)) OR
 					(reg_q813 AND symb_decoder(16#24#)) OR
 					(reg_q813 AND symb_decoder(16#76#)) OR
 					(reg_q813 AND symb_decoder(16#d2#)) OR
 					(reg_q813 AND symb_decoder(16#d9#)) OR
 					(reg_q813 AND symb_decoder(16#b5#)) OR
 					(reg_q813 AND symb_decoder(16#32#)) OR
 					(reg_q813 AND symb_decoder(16#c6#)) OR
 					(reg_q813 AND symb_decoder(16#1f#)) OR
 					(reg_q813 AND symb_decoder(16#89#)) OR
 					(reg_q813 AND symb_decoder(16#3b#)) OR
 					(reg_q813 AND symb_decoder(16#f6#)) OR
 					(reg_q813 AND symb_decoder(16#29#)) OR
 					(reg_q813 AND symb_decoder(16#4e#)) OR
 					(reg_q791 AND symb_decoder(16#95#)) OR
 					(reg_q791 AND symb_decoder(16#33#)) OR
 					(reg_q791 AND symb_decoder(16#74#)) OR
 					(reg_q791 AND symb_decoder(16#59#)) OR
 					(reg_q791 AND symb_decoder(16#91#)) OR
 					(reg_q791 AND symb_decoder(16#f9#)) OR
 					(reg_q791 AND symb_decoder(16#38#)) OR
 					(reg_q791 AND symb_decoder(16#cc#)) OR
 					(reg_q791 AND symb_decoder(16#b9#)) OR
 					(reg_q791 AND symb_decoder(16#e2#)) OR
 					(reg_q791 AND symb_decoder(16#a5#)) OR
 					(reg_q791 AND symb_decoder(16#04#)) OR
 					(reg_q791 AND symb_decoder(16#c0#)) OR
 					(reg_q791 AND symb_decoder(16#55#)) OR
 					(reg_q791 AND symb_decoder(16#cf#)) OR
 					(reg_q791 AND symb_decoder(16#c5#)) OR
 					(reg_q791 AND symb_decoder(16#84#)) OR
 					(reg_q791 AND symb_decoder(16#61#)) OR
 					(reg_q791 AND symb_decoder(16#4b#)) OR
 					(reg_q791 AND symb_decoder(16#a6#)) OR
 					(reg_q791 AND symb_decoder(16#c4#)) OR
 					(reg_q791 AND symb_decoder(16#29#)) OR
 					(reg_q791 AND symb_decoder(16#28#)) OR
 					(reg_q791 AND symb_decoder(16#4e#)) OR
 					(reg_q791 AND symb_decoder(16#a4#)) OR
 					(reg_q791 AND symb_decoder(16#9c#)) OR
 					(reg_q791 AND symb_decoder(16#5e#)) OR
 					(reg_q791 AND symb_decoder(16#e4#)) OR
 					(reg_q791 AND symb_decoder(16#32#)) OR
 					(reg_q791 AND symb_decoder(16#af#)) OR
 					(reg_q791 AND symb_decoder(16#2f#)) OR
 					(reg_q791 AND symb_decoder(16#9d#)) OR
 					(reg_q791 AND symb_decoder(16#26#)) OR
 					(reg_q791 AND symb_decoder(16#e7#)) OR
 					(reg_q791 AND symb_decoder(16#f8#)) OR
 					(reg_q791 AND symb_decoder(16#15#)) OR
 					(reg_q791 AND symb_decoder(16#de#)) OR
 					(reg_q791 AND symb_decoder(16#e1#)) OR
 					(reg_q791 AND symb_decoder(16#ba#)) OR
 					(reg_q791 AND symb_decoder(16#01#)) OR
 					(reg_q791 AND symb_decoder(16#0e#)) OR
 					(reg_q791 AND symb_decoder(16#f1#)) OR
 					(reg_q791 AND symb_decoder(16#6d#)) OR
 					(reg_q791 AND symb_decoder(16#cd#)) OR
 					(reg_q791 AND symb_decoder(16#54#)) OR
 					(reg_q791 AND symb_decoder(16#3a#)) OR
 					(reg_q791 AND symb_decoder(16#ce#)) OR
 					(reg_q791 AND symb_decoder(16#18#)) OR
 					(reg_q791 AND symb_decoder(16#d4#)) OR
 					(reg_q791 AND symb_decoder(16#17#)) OR
 					(reg_q791 AND symb_decoder(16#b4#)) OR
 					(reg_q791 AND symb_decoder(16#da#)) OR
 					(reg_q791 AND symb_decoder(16#89#)) OR
 					(reg_q791 AND symb_decoder(16#51#)) OR
 					(reg_q791 AND symb_decoder(16#5b#)) OR
 					(reg_q791 AND symb_decoder(16#cb#)) OR
 					(reg_q791 AND symb_decoder(16#9f#)) OR
 					(reg_q791 AND symb_decoder(16#98#)) OR
 					(reg_q791 AND symb_decoder(16#75#)) OR
 					(reg_q791 AND symb_decoder(16#a7#)) OR
 					(reg_q791 AND symb_decoder(16#63#)) OR
 					(reg_q791 AND symb_decoder(16#11#)) OR
 					(reg_q791 AND symb_decoder(16#58#)) OR
 					(reg_q791 AND symb_decoder(16#13#)) OR
 					(reg_q791 AND symb_decoder(16#b3#)) OR
 					(reg_q791 AND symb_decoder(16#99#)) OR
 					(reg_q791 AND symb_decoder(16#c2#)) OR
 					(reg_q791 AND symb_decoder(16#8e#)) OR
 					(reg_q791 AND symb_decoder(16#21#)) OR
 					(reg_q791 AND symb_decoder(16#06#)) OR
 					(reg_q791 AND symb_decoder(16#30#)) OR
 					(reg_q791 AND symb_decoder(16#27#)) OR
 					(reg_q791 AND symb_decoder(16#25#)) OR
 					(reg_q791 AND symb_decoder(16#5a#)) OR
 					(reg_q791 AND symb_decoder(16#ef#)) OR
 					(reg_q791 AND symb_decoder(16#87#)) OR
 					(reg_q791 AND symb_decoder(16#85#)) OR
 					(reg_q791 AND symb_decoder(16#d1#)) OR
 					(reg_q791 AND symb_decoder(16#2b#)) OR
 					(reg_q791 AND symb_decoder(16#78#)) OR
 					(reg_q791 AND symb_decoder(16#1a#)) OR
 					(reg_q791 AND symb_decoder(16#19#)) OR
 					(reg_q791 AND symb_decoder(16#93#)) OR
 					(reg_q791 AND symb_decoder(16#ca#)) OR
 					(reg_q791 AND symb_decoder(16#e3#)) OR
 					(reg_q791 AND symb_decoder(16#90#)) OR
 					(reg_q791 AND symb_decoder(16#d0#)) OR
 					(reg_q791 AND symb_decoder(16#ae#)) OR
 					(reg_q791 AND symb_decoder(16#00#)) OR
 					(reg_q791 AND symb_decoder(16#71#)) OR
 					(reg_q791 AND symb_decoder(16#b1#)) OR
 					(reg_q791 AND symb_decoder(16#3c#)) OR
 					(reg_q791 AND symb_decoder(16#02#)) OR
 					(reg_q791 AND symb_decoder(16#62#)) OR
 					(reg_q791 AND symb_decoder(16#d5#)) OR
 					(reg_q791 AND symb_decoder(16#1e#)) OR
 					(reg_q791 AND symb_decoder(16#f7#)) OR
 					(reg_q791 AND symb_decoder(16#83#)) OR
 					(reg_q791 AND symb_decoder(16#8c#)) OR
 					(reg_q791 AND symb_decoder(16#4a#)) OR
 					(reg_q791 AND symb_decoder(16#7b#)) OR
 					(reg_q791 AND symb_decoder(16#5d#)) OR
 					(reg_q791 AND symb_decoder(16#7c#)) OR
 					(reg_q791 AND symb_decoder(16#c1#)) OR
 					(reg_q791 AND symb_decoder(16#6c#)) OR
 					(reg_q791 AND symb_decoder(16#dc#)) OR
 					(reg_q791 AND symb_decoder(16#fa#)) OR
 					(reg_q791 AND symb_decoder(16#88#)) OR
 					(reg_q791 AND symb_decoder(16#2e#)) OR
 					(reg_q791 AND symb_decoder(16#f6#)) OR
 					(reg_q791 AND symb_decoder(16#8d#)) OR
 					(reg_q791 AND symb_decoder(16#72#)) OR
 					(reg_q791 AND symb_decoder(16#bc#)) OR
 					(reg_q791 AND symb_decoder(16#a9#)) OR
 					(reg_q791 AND symb_decoder(16#76#)) OR
 					(reg_q791 AND symb_decoder(16#b0#)) OR
 					(reg_q791 AND symb_decoder(16#d7#)) OR
 					(reg_q791 AND symb_decoder(16#24#)) OR
 					(reg_q791 AND symb_decoder(16#46#)) OR
 					(reg_q791 AND symb_decoder(16#66#)) OR
 					(reg_q791 AND symb_decoder(16#fc#)) OR
 					(reg_q791 AND symb_decoder(16#92#)) OR
 					(reg_q791 AND symb_decoder(16#20#)) OR
 					(reg_q791 AND symb_decoder(16#c3#)) OR
 					(reg_q791 AND symb_decoder(16#0c#)) OR
 					(reg_q791 AND symb_decoder(16#8a#)) OR
 					(reg_q791 AND symb_decoder(16#86#)) OR
 					(reg_q791 AND symb_decoder(16#ac#)) OR
 					(reg_q791 AND symb_decoder(16#a3#)) OR
 					(reg_q791 AND symb_decoder(16#7a#)) OR
 					(reg_q791 AND symb_decoder(16#d6#)) OR
 					(reg_q791 AND symb_decoder(16#6a#)) OR
 					(reg_q791 AND symb_decoder(16#70#)) OR
 					(reg_q791 AND symb_decoder(16#68#)) OR
 					(reg_q791 AND symb_decoder(16#41#)) OR
 					(reg_q791 AND symb_decoder(16#65#)) OR
 					(reg_q791 AND symb_decoder(16#b7#)) OR
 					(reg_q791 AND symb_decoder(16#82#)) OR
 					(reg_q791 AND symb_decoder(16#a2#)) OR
 					(reg_q791 AND symb_decoder(16#aa#)) OR
 					(reg_q791 AND symb_decoder(16#be#)) OR
 					(reg_q791 AND symb_decoder(16#05#)) OR
 					(reg_q791 AND symb_decoder(16#2c#)) OR
 					(reg_q791 AND symb_decoder(16#eb#)) OR
 					(reg_q791 AND symb_decoder(16#34#)) OR
 					(reg_q791 AND symb_decoder(16#40#)) OR
 					(reg_q791 AND symb_decoder(16#e0#)) OR
 					(reg_q791 AND symb_decoder(16#07#)) OR
 					(reg_q791 AND symb_decoder(16#b8#)) OR
 					(reg_q791 AND symb_decoder(16#73#)) OR
 					(reg_q791 AND symb_decoder(16#12#)) OR
 					(reg_q791 AND symb_decoder(16#6e#)) OR
 					(reg_q791 AND symb_decoder(16#80#)) OR
 					(reg_q791 AND symb_decoder(16#79#)) OR
 					(reg_q791 AND symb_decoder(16#2d#)) OR
 					(reg_q791 AND symb_decoder(16#44#)) OR
 					(reg_q791 AND symb_decoder(16#1f#)) OR
 					(reg_q791 AND symb_decoder(16#bd#)) OR
 					(reg_q791 AND symb_decoder(16#47#)) OR
 					(reg_q791 AND symb_decoder(16#42#)) OR
 					(reg_q791 AND symb_decoder(16#b5#)) OR
 					(reg_q791 AND symb_decoder(16#ea#)) OR
 					(reg_q791 AND symb_decoder(16#a1#)) OR
 					(reg_q791 AND symb_decoder(16#f4#)) OR
 					(reg_q791 AND symb_decoder(16#4f#)) OR
 					(reg_q791 AND symb_decoder(16#81#)) OR
 					(reg_q791 AND symb_decoder(16#c7#)) OR
 					(reg_q791 AND symb_decoder(16#77#)) OR
 					(reg_q791 AND symb_decoder(16#22#)) OR
 					(reg_q791 AND symb_decoder(16#3b#)) OR
 					(reg_q791 AND symb_decoder(16#1b#)) OR
 					(reg_q791 AND symb_decoder(16#6f#)) OR
 					(reg_q791 AND symb_decoder(16#bf#)) OR
 					(reg_q791 AND symb_decoder(16#8f#)) OR
 					(reg_q791 AND symb_decoder(16#df#)) OR
 					(reg_q791 AND symb_decoder(16#67#)) OR
 					(reg_q791 AND symb_decoder(16#7f#)) OR
 					(reg_q791 AND symb_decoder(16#3d#)) OR
 					(reg_q791 AND symb_decoder(16#4d#)) OR
 					(reg_q791 AND symb_decoder(16#ff#)) OR
 					(reg_q791 AND symb_decoder(16#9e#)) OR
 					(reg_q791 AND symb_decoder(16#45#)) OR
 					(reg_q791 AND symb_decoder(16#1d#)) OR
 					(reg_q791 AND symb_decoder(16#48#)) OR
 					(reg_q791 AND symb_decoder(16#9a#)) OR
 					(reg_q791 AND symb_decoder(16#0f#)) OR
 					(reg_q791 AND symb_decoder(16#f3#)) OR
 					(reg_q791 AND symb_decoder(16#e8#)) OR
 					(reg_q791 AND symb_decoder(16#dd#)) OR
 					(reg_q791 AND symb_decoder(16#49#)) OR
 					(reg_q791 AND symb_decoder(16#36#)) OR
 					(reg_q791 AND symb_decoder(16#60#)) OR
 					(reg_q791 AND symb_decoder(16#ab#)) OR
 					(reg_q791 AND symb_decoder(16#f0#)) OR
 					(reg_q791 AND symb_decoder(16#97#)) OR
 					(reg_q791 AND symb_decoder(16#e9#)) OR
 					(reg_q791 AND symb_decoder(16#0b#)) OR
 					(reg_q791 AND symb_decoder(16#1c#)) OR
 					(reg_q791 AND symb_decoder(16#c8#)) OR
 					(reg_q791 AND symb_decoder(16#d2#)) OR
 					(reg_q791 AND symb_decoder(16#10#)) OR
 					(reg_q791 AND symb_decoder(16#d3#)) OR
 					(reg_q791 AND symb_decoder(16#8b#)) OR
 					(reg_q791 AND symb_decoder(16#fd#)) OR
 					(reg_q791 AND symb_decoder(16#a8#)) OR
 					(reg_q791 AND symb_decoder(16#14#)) OR
 					(reg_q791 AND symb_decoder(16#e5#)) OR
 					(reg_q791 AND symb_decoder(16#31#)) OR
 					(reg_q791 AND symb_decoder(16#c6#)) OR
 					(reg_q791 AND symb_decoder(16#e6#)) OR
 					(reg_q791 AND symb_decoder(16#16#)) OR
 					(reg_q791 AND symb_decoder(16#53#)) OR
 					(reg_q791 AND symb_decoder(16#9b#)) OR
 					(reg_q791 AND symb_decoder(16#b6#)) OR
 					(reg_q791 AND symb_decoder(16#c9#)) OR
 					(reg_q791 AND symb_decoder(16#2a#)) OR
 					(reg_q791 AND symb_decoder(16#fe#)) OR
 					(reg_q791 AND symb_decoder(16#4c#)) OR
 					(reg_q791 AND symb_decoder(16#94#)) OR
 					(reg_q791 AND symb_decoder(16#6b#)) OR
 					(reg_q791 AND symb_decoder(16#db#)) OR
 					(reg_q791 AND symb_decoder(16#23#)) OR
 					(reg_q791 AND symb_decoder(16#7e#)) OR
 					(reg_q791 AND symb_decoder(16#f5#)) OR
 					(reg_q791 AND symb_decoder(16#56#)) OR
 					(reg_q791 AND symb_decoder(16#3e#)) OR
 					(reg_q791 AND symb_decoder(16#37#)) OR
 					(reg_q791 AND symb_decoder(16#d8#)) OR
 					(reg_q791 AND symb_decoder(16#3f#)) OR
 					(reg_q791 AND symb_decoder(16#52#)) OR
 					(reg_q791 AND symb_decoder(16#03#)) OR
 					(reg_q791 AND symb_decoder(16#35#)) OR
 					(reg_q791 AND symb_decoder(16#08#)) OR
 					(reg_q791 AND symb_decoder(16#5f#)) OR
 					(reg_q791 AND symb_decoder(16#69#)) OR
 					(reg_q791 AND symb_decoder(16#64#)) OR
 					(reg_q791 AND symb_decoder(16#f2#)) OR
 					(reg_q791 AND symb_decoder(16#ec#)) OR
 					(reg_q791 AND symb_decoder(16#09#)) OR
 					(reg_q791 AND symb_decoder(16#bb#)) OR
 					(reg_q791 AND symb_decoder(16#7d#)) OR
 					(reg_q791 AND symb_decoder(16#d9#)) OR
 					(reg_q791 AND symb_decoder(16#ee#)) OR
 					(reg_q791 AND symb_decoder(16#50#)) OR
 					(reg_q791 AND symb_decoder(16#ad#)) OR
 					(reg_q791 AND symb_decoder(16#b2#)) OR
 					(reg_q791 AND symb_decoder(16#fb#)) OR
 					(reg_q791 AND symb_decoder(16#96#)) OR
 					(reg_q791 AND symb_decoder(16#57#)) OR
 					(reg_q791 AND symb_decoder(16#43#)) OR
 					(reg_q791 AND symb_decoder(16#39#)) OR
 					(reg_q791 AND symb_decoder(16#a0#)) OR
 					(reg_q791 AND symb_decoder(16#ed#)) OR
 					(reg_q791 AND symb_decoder(16#5c#));
reg_q1298_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1297 AND symb_decoder(16#0d#)) OR
 					(reg_q1297 AND symb_decoder(16#0a#));
reg_q901_in <= (reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q901 AND symb_decoder(16#31#)) OR
 					(reg_q901 AND symb_decoder(16#30#)) OR
 					(reg_q901 AND symb_decoder(16#35#)) OR
 					(reg_q901 AND symb_decoder(16#38#)) OR
 					(reg_q901 AND symb_decoder(16#37#)) OR
 					(reg_q901 AND symb_decoder(16#36#)) OR
 					(reg_q901 AND symb_decoder(16#39#)) OR
 					(reg_q901 AND symb_decoder(16#33#)) OR
 					(reg_q901 AND symb_decoder(16#32#)) OR
 					(reg_q901 AND symb_decoder(16#34#)) OR
 					(reg_q900 AND symb_decoder(16#34#)) OR
 					(reg_q900 AND symb_decoder(16#36#)) OR
 					(reg_q900 AND symb_decoder(16#32#)) OR
 					(reg_q900 AND symb_decoder(16#33#)) OR
 					(reg_q900 AND symb_decoder(16#38#)) OR
 					(reg_q900 AND symb_decoder(16#39#)) OR
 					(reg_q900 AND symb_decoder(16#35#)) OR
 					(reg_q900 AND symb_decoder(16#31#)) OR
 					(reg_q900 AND symb_decoder(16#37#)) OR
 					(reg_q900 AND symb_decoder(16#30#));
reg_q781_in <= (reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q780 AND symb_decoder(16#44#)) OR
 					(reg_q780 AND symb_decoder(16#64#));
reg_q1052_in <= (reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q1051 AND symb_decoder(16#45#)) OR
 					(reg_q1051 AND symb_decoder(16#65#));
reg_q2126_in <= (reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2125 AND symb_decoder(16#77#)) OR
 					(reg_q2125 AND symb_decoder(16#57#));
reg_q1523_in <= (reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q1522 AND symb_decoder(16#6e#)) OR
 					(reg_q1522 AND symb_decoder(16#4e#));
reg_q2587_in <= (reg_q2585 AND symb_decoder(16#63#)) OR
 					(reg_q2585 AND symb_decoder(16#43#));
reg_q1995_in <= (reg_q1993 AND symb_decoder(16#23#));
reg_fullgraph45_init <= "0000";

reg_fullgraph45_sel <= "0000000" & reg_q1995_in & reg_q2587_in & reg_q1523_in & reg_q2126_in & reg_q1052_in & reg_q781_in & reg_q901_in & reg_q1298_in & reg_q813_in;

	--coder fullgraph45
with reg_fullgraph45_sel select
reg_fullgraph45_in <=
	"0001" when "0000000000000001",
	"0010" when "0000000000000010",
	"0011" when "0000000000000100",
	"0100" when "0000000000001000",
	"0101" when "0000000000010000",
	"0110" when "0000000000100000",
	"0111" when "0000000001000000",
	"1000" when "0000000010000000",
	"1001" when "0000000100000000",
	"0000" when others;
 --end coder

	p_reg_fullgraph45: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph45 <= reg_fullgraph45_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph45 <= reg_fullgraph45_init;
        else
          reg_fullgraph45 <= reg_fullgraph45_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph45

		reg_q813 <= '1' when reg_fullgraph45 = "0001" else '0'; 
		reg_q1298 <= '1' when reg_fullgraph45 = "0010" else '0'; 
		reg_q901 <= '1' when reg_fullgraph45 = "0011" else '0'; 
		reg_q781 <= '1' when reg_fullgraph45 = "0100" else '0'; 
		reg_q1052 <= '1' when reg_fullgraph45 = "0101" else '0'; 
		reg_q2126 <= '1' when reg_fullgraph45 = "0110" else '0'; 
		reg_q1523 <= '1' when reg_fullgraph45 = "0111" else '0'; 
		reg_q2587 <= '1' when reg_fullgraph45 = "1000" else '0'; 
		reg_q1995 <= '1' when reg_fullgraph45 = "1001" else '0'; 
--end decoder 

reg_q714_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q714 AND symb_decoder(16#45#)) OR
 					(reg_q714 AND symb_decoder(16#42#)) OR
 					(reg_q714 AND symb_decoder(16#57#)) OR
 					(reg_q714 AND symb_decoder(16#2c#)) OR
 					(reg_q714 AND symb_decoder(16#e1#)) OR
 					(reg_q714 AND symb_decoder(16#29#)) OR
 					(reg_q714 AND symb_decoder(16#5c#)) OR
 					(reg_q714 AND symb_decoder(16#5f#)) OR
 					(reg_q714 AND symb_decoder(16#fc#)) OR
 					(reg_q714 AND symb_decoder(16#c1#)) OR
 					(reg_q714 AND symb_decoder(16#c4#)) OR
 					(reg_q714 AND symb_decoder(16#44#)) OR
 					(reg_q714 AND symb_decoder(16#f3#)) OR
 					(reg_q714 AND symb_decoder(16#9c#)) OR
 					(reg_q714 AND symb_decoder(16#08#)) OR
 					(reg_q714 AND symb_decoder(16#2e#)) OR
 					(reg_q714 AND symb_decoder(16#b1#)) OR
 					(reg_q714 AND symb_decoder(16#3e#)) OR
 					(reg_q714 AND symb_decoder(16#af#)) OR
 					(reg_q714 AND symb_decoder(16#f9#)) OR
 					(reg_q714 AND symb_decoder(16#ca#)) OR
 					(reg_q714 AND symb_decoder(16#6d#)) OR
 					(reg_q714 AND symb_decoder(16#30#)) OR
 					(reg_q714 AND symb_decoder(16#77#)) OR
 					(reg_q714 AND symb_decoder(16#92#)) OR
 					(reg_q714 AND symb_decoder(16#24#)) OR
 					(reg_q714 AND symb_decoder(16#4a#)) OR
 					(reg_q714 AND symb_decoder(16#48#)) OR
 					(reg_q714 AND symb_decoder(16#d6#)) OR
 					(reg_q714 AND symb_decoder(16#b2#)) OR
 					(reg_q714 AND symb_decoder(16#fb#)) OR
 					(reg_q714 AND symb_decoder(16#90#)) OR
 					(reg_q714 AND symb_decoder(16#50#)) OR
 					(reg_q714 AND symb_decoder(16#88#)) OR
 					(reg_q714 AND symb_decoder(16#5d#)) OR
 					(reg_q714 AND symb_decoder(16#ac#)) OR
 					(reg_q714 AND symb_decoder(16#b8#)) OR
 					(reg_q714 AND symb_decoder(16#55#)) OR
 					(reg_q714 AND symb_decoder(16#84#)) OR
 					(reg_q714 AND symb_decoder(16#2f#)) OR
 					(reg_q714 AND symb_decoder(16#63#)) OR
 					(reg_q714 AND symb_decoder(16#d9#)) OR
 					(reg_q714 AND symb_decoder(16#0a#)) OR
 					(reg_q714 AND symb_decoder(16#3b#)) OR
 					(reg_q714 AND symb_decoder(16#de#)) OR
 					(reg_q714 AND symb_decoder(16#fa#)) OR
 					(reg_q714 AND symb_decoder(16#35#)) OR
 					(reg_q714 AND symb_decoder(16#46#)) OR
 					(reg_q714 AND symb_decoder(16#cf#)) OR
 					(reg_q714 AND symb_decoder(16#54#)) OR
 					(reg_q714 AND symb_decoder(16#cd#)) OR
 					(reg_q714 AND symb_decoder(16#e8#)) OR
 					(reg_q714 AND symb_decoder(16#df#)) OR
 					(reg_q714 AND symb_decoder(16#39#)) OR
 					(reg_q714 AND symb_decoder(16#4e#)) OR
 					(reg_q714 AND symb_decoder(16#9f#)) OR
 					(reg_q714 AND symb_decoder(16#ed#)) OR
 					(reg_q714 AND symb_decoder(16#da#)) OR
 					(reg_q714 AND symb_decoder(16#79#)) OR
 					(reg_q714 AND symb_decoder(16#7e#)) OR
 					(reg_q714 AND symb_decoder(16#cb#)) OR
 					(reg_q714 AND symb_decoder(16#89#)) OR
 					(reg_q714 AND symb_decoder(16#07#)) OR
 					(reg_q714 AND symb_decoder(16#16#)) OR
 					(reg_q714 AND symb_decoder(16#f0#)) OR
 					(reg_q714 AND symb_decoder(16#3d#)) OR
 					(reg_q714 AND symb_decoder(16#a4#)) OR
 					(reg_q714 AND symb_decoder(16#ba#)) OR
 					(reg_q714 AND symb_decoder(16#1c#)) OR
 					(reg_q714 AND symb_decoder(16#d7#)) OR
 					(reg_q714 AND symb_decoder(16#22#)) OR
 					(reg_q714 AND symb_decoder(16#c2#)) OR
 					(reg_q714 AND symb_decoder(16#e6#)) OR
 					(reg_q714 AND symb_decoder(16#bf#)) OR
 					(reg_q714 AND symb_decoder(16#19#)) OR
 					(reg_q714 AND symb_decoder(16#e5#)) OR
 					(reg_q714 AND symb_decoder(16#a3#)) OR
 					(reg_q714 AND symb_decoder(16#ce#)) OR
 					(reg_q714 AND symb_decoder(16#6e#)) OR
 					(reg_q714 AND symb_decoder(16#d2#)) OR
 					(reg_q714 AND symb_decoder(16#a7#)) OR
 					(reg_q714 AND symb_decoder(16#5a#)) OR
 					(reg_q714 AND symb_decoder(16#d3#)) OR
 					(reg_q714 AND symb_decoder(16#17#)) OR
 					(reg_q714 AND symb_decoder(16#47#)) OR
 					(reg_q714 AND symb_decoder(16#c0#)) OR
 					(reg_q714 AND symb_decoder(16#ab#)) OR
 					(reg_q714 AND symb_decoder(16#a9#)) OR
 					(reg_q714 AND symb_decoder(16#7d#)) OR
 					(reg_q714 AND symb_decoder(16#ae#)) OR
 					(reg_q714 AND symb_decoder(16#6b#)) OR
 					(reg_q714 AND symb_decoder(16#72#)) OR
 					(reg_q714 AND symb_decoder(16#7f#)) OR
 					(reg_q714 AND symb_decoder(16#1b#)) OR
 					(reg_q714 AND symb_decoder(16#ef#)) OR
 					(reg_q714 AND symb_decoder(16#c7#)) OR
 					(reg_q714 AND symb_decoder(16#c9#)) OR
 					(reg_q714 AND symb_decoder(16#28#)) OR
 					(reg_q714 AND symb_decoder(16#97#)) OR
 					(reg_q714 AND symb_decoder(16#15#)) OR
 					(reg_q714 AND symb_decoder(16#95#)) OR
 					(reg_q714 AND symb_decoder(16#94#)) OR
 					(reg_q714 AND symb_decoder(16#e3#)) OR
 					(reg_q714 AND symb_decoder(16#a0#)) OR
 					(reg_q714 AND symb_decoder(16#65#)) OR
 					(reg_q714 AND symb_decoder(16#c3#)) OR
 					(reg_q714 AND symb_decoder(16#f2#)) OR
 					(reg_q714 AND symb_decoder(16#d1#)) OR
 					(reg_q714 AND symb_decoder(16#bb#)) OR
 					(reg_q714 AND symb_decoder(16#e4#)) OR
 					(reg_q714 AND symb_decoder(16#87#)) OR
 					(reg_q714 AND symb_decoder(16#59#)) OR
 					(reg_q714 AND symb_decoder(16#9a#)) OR
 					(reg_q714 AND symb_decoder(16#b0#)) OR
 					(reg_q714 AND symb_decoder(16#5b#)) OR
 					(reg_q714 AND symb_decoder(16#bc#)) OR
 					(reg_q714 AND symb_decoder(16#eb#)) OR
 					(reg_q714 AND symb_decoder(16#ad#)) OR
 					(reg_q714 AND symb_decoder(16#dd#)) OR
 					(reg_q714 AND symb_decoder(16#2a#)) OR
 					(reg_q714 AND symb_decoder(16#27#)) OR
 					(reg_q714 AND symb_decoder(16#d5#)) OR
 					(reg_q714 AND symb_decoder(16#86#)) OR
 					(reg_q714 AND symb_decoder(16#3f#)) OR
 					(reg_q714 AND symb_decoder(16#f7#)) OR
 					(reg_q714 AND symb_decoder(16#e0#)) OR
 					(reg_q714 AND symb_decoder(16#fe#)) OR
 					(reg_q714 AND symb_decoder(16#85#)) OR
 					(reg_q714 AND symb_decoder(16#1f#)) OR
 					(reg_q714 AND symb_decoder(16#0d#)) OR
 					(reg_q714 AND symb_decoder(16#dc#)) OR
 					(reg_q714 AND symb_decoder(16#66#)) OR
 					(reg_q714 AND symb_decoder(16#83#)) OR
 					(reg_q714 AND symb_decoder(16#41#)) OR
 					(reg_q714 AND symb_decoder(16#00#)) OR
 					(reg_q714 AND symb_decoder(16#26#)) OR
 					(reg_q714 AND symb_decoder(16#01#)) OR
 					(reg_q714 AND symb_decoder(16#9b#)) OR
 					(reg_q714 AND symb_decoder(16#81#)) OR
 					(reg_q714 AND symb_decoder(16#f5#)) OR
 					(reg_q714 AND symb_decoder(16#b9#)) OR
 					(reg_q714 AND symb_decoder(16#52#)) OR
 					(reg_q714 AND symb_decoder(16#d4#)) OR
 					(reg_q714 AND symb_decoder(16#f4#)) OR
 					(reg_q714 AND symb_decoder(16#53#)) OR
 					(reg_q714 AND symb_decoder(16#4f#)) OR
 					(reg_q714 AND symb_decoder(16#2d#)) OR
 					(reg_q714 AND symb_decoder(16#51#)) OR
 					(reg_q714 AND symb_decoder(16#06#)) OR
 					(reg_q714 AND symb_decoder(16#db#)) OR
 					(reg_q714 AND symb_decoder(16#73#)) OR
 					(reg_q714 AND symb_decoder(16#10#)) OR
 					(reg_q714 AND symb_decoder(16#64#)) OR
 					(reg_q714 AND symb_decoder(16#cc#)) OR
 					(reg_q714 AND symb_decoder(16#71#)) OR
 					(reg_q714 AND symb_decoder(16#5e#)) OR
 					(reg_q714 AND symb_decoder(16#6f#)) OR
 					(reg_q714 AND symb_decoder(16#0c#)) OR
 					(reg_q714 AND symb_decoder(16#ff#)) OR
 					(reg_q714 AND symb_decoder(16#03#)) OR
 					(reg_q714 AND symb_decoder(16#4c#)) OR
 					(reg_q714 AND symb_decoder(16#93#)) OR
 					(reg_q714 AND symb_decoder(16#1a#)) OR
 					(reg_q714 AND symb_decoder(16#7b#)) OR
 					(reg_q714 AND symb_decoder(16#ea#)) OR
 					(reg_q714 AND symb_decoder(16#e9#)) OR
 					(reg_q714 AND symb_decoder(16#0f#)) OR
 					(reg_q714 AND symb_decoder(16#b4#)) OR
 					(reg_q714 AND symb_decoder(16#8a#)) OR
 					(reg_q714 AND symb_decoder(16#b6#)) OR
 					(reg_q714 AND symb_decoder(16#75#)) OR
 					(reg_q714 AND symb_decoder(16#32#)) OR
 					(reg_q714 AND symb_decoder(16#96#)) OR
 					(reg_q714 AND symb_decoder(16#78#)) OR
 					(reg_q714 AND symb_decoder(16#9d#)) OR
 					(reg_q714 AND symb_decoder(16#40#)) OR
 					(reg_q714 AND symb_decoder(16#18#)) OR
 					(reg_q714 AND symb_decoder(16#82#)) OR
 					(reg_q714 AND symb_decoder(16#c5#)) OR
 					(reg_q714 AND symb_decoder(16#69#)) OR
 					(reg_q714 AND symb_decoder(16#f1#)) OR
 					(reg_q714 AND symb_decoder(16#9e#)) OR
 					(reg_q714 AND symb_decoder(16#37#)) OR
 					(reg_q714 AND symb_decoder(16#4b#)) OR
 					(reg_q714 AND symb_decoder(16#0b#)) OR
 					(reg_q714 AND symb_decoder(16#be#)) OR
 					(reg_q714 AND symb_decoder(16#80#)) OR
 					(reg_q714 AND symb_decoder(16#c8#)) OR
 					(reg_q714 AND symb_decoder(16#a2#)) OR
 					(reg_q714 AND symb_decoder(16#3c#)) OR
 					(reg_q714 AND symb_decoder(16#3a#)) OR
 					(reg_q714 AND symb_decoder(16#b7#)) OR
 					(reg_q714 AND symb_decoder(16#8e#)) OR
 					(reg_q714 AND symb_decoder(16#20#)) OR
 					(reg_q714 AND symb_decoder(16#fd#)) OR
 					(reg_q714 AND symb_decoder(16#1d#)) OR
 					(reg_q714 AND symb_decoder(16#99#)) OR
 					(reg_q714 AND symb_decoder(16#58#)) OR
 					(reg_q714 AND symb_decoder(16#49#)) OR
 					(reg_q714 AND symb_decoder(16#a8#)) OR
 					(reg_q714 AND symb_decoder(16#98#)) OR
 					(reg_q714 AND symb_decoder(16#31#)) OR
 					(reg_q714 AND symb_decoder(16#e7#)) OR
 					(reg_q714 AND symb_decoder(16#02#)) OR
 					(reg_q714 AND symb_decoder(16#11#)) OR
 					(reg_q714 AND symb_decoder(16#68#)) OR
 					(reg_q714 AND symb_decoder(16#a1#)) OR
 					(reg_q714 AND symb_decoder(16#7a#)) OR
 					(reg_q714 AND symb_decoder(16#8b#)) OR
 					(reg_q714 AND symb_decoder(16#8d#)) OR
 					(reg_q714 AND symb_decoder(16#bd#)) OR
 					(reg_q714 AND symb_decoder(16#8c#)) OR
 					(reg_q714 AND symb_decoder(16#09#)) OR
 					(reg_q714 AND symb_decoder(16#56#)) OR
 					(reg_q714 AND symb_decoder(16#7c#)) OR
 					(reg_q714 AND symb_decoder(16#a6#)) OR
 					(reg_q714 AND symb_decoder(16#62#)) OR
 					(reg_q714 AND symb_decoder(16#60#)) OR
 					(reg_q714 AND symb_decoder(16#04#)) OR
 					(reg_q714 AND symb_decoder(16#25#)) OR
 					(reg_q714 AND symb_decoder(16#6a#)) OR
 					(reg_q714 AND symb_decoder(16#2b#)) OR
 					(reg_q714 AND symb_decoder(16#d8#)) OR
 					(reg_q714 AND symb_decoder(16#23#)) OR
 					(reg_q714 AND symb_decoder(16#36#)) OR
 					(reg_q714 AND symb_decoder(16#c6#)) OR
 					(reg_q714 AND symb_decoder(16#61#)) OR
 					(reg_q714 AND symb_decoder(16#aa#)) OR
 					(reg_q714 AND symb_decoder(16#05#)) OR
 					(reg_q714 AND symb_decoder(16#0e#)) OR
 					(reg_q714 AND symb_decoder(16#ee#)) OR
 					(reg_q714 AND symb_decoder(16#67#)) OR
 					(reg_q714 AND symb_decoder(16#b5#)) OR
 					(reg_q714 AND symb_decoder(16#14#)) OR
 					(reg_q714 AND symb_decoder(16#74#)) OR
 					(reg_q714 AND symb_decoder(16#12#)) OR
 					(reg_q714 AND symb_decoder(16#f8#)) OR
 					(reg_q714 AND symb_decoder(16#b3#)) OR
 					(reg_q714 AND symb_decoder(16#1e#)) OR
 					(reg_q714 AND symb_decoder(16#4d#)) OR
 					(reg_q714 AND symb_decoder(16#34#)) OR
 					(reg_q714 AND symb_decoder(16#43#)) OR
 					(reg_q714 AND symb_decoder(16#21#)) OR
 					(reg_q714 AND symb_decoder(16#38#)) OR
 					(reg_q714 AND symb_decoder(16#76#)) OR
 					(reg_q714 AND symb_decoder(16#13#)) OR
 					(reg_q714 AND symb_decoder(16#8f#)) OR
 					(reg_q714 AND symb_decoder(16#d0#)) OR
 					(reg_q714 AND symb_decoder(16#70#)) OR
 					(reg_q714 AND symb_decoder(16#33#)) OR
 					(reg_q714 AND symb_decoder(16#91#)) OR
 					(reg_q714 AND symb_decoder(16#f6#)) OR
 					(reg_q714 AND symb_decoder(16#a5#)) OR
 					(reg_q714 AND symb_decoder(16#6c#)) OR
 					(reg_q714 AND symb_decoder(16#ec#)) OR
 					(reg_q714 AND symb_decoder(16#e2#));
reg_q714_init <= '0' ;
	p_reg_q714: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q714 <= reg_q714_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q714 <= reg_q714_init;
        else
          reg_q714 <= reg_q714_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1544_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q1544 AND symb_decoder(16#48#)) OR
 					(reg_q1544 AND symb_decoder(16#d7#)) OR
 					(reg_q1544 AND symb_decoder(16#e2#)) OR
 					(reg_q1544 AND symb_decoder(16#4f#)) OR
 					(reg_q1544 AND symb_decoder(16#ba#)) OR
 					(reg_q1544 AND symb_decoder(16#3b#)) OR
 					(reg_q1544 AND symb_decoder(16#6b#)) OR
 					(reg_q1544 AND symb_decoder(16#27#)) OR
 					(reg_q1544 AND symb_decoder(16#75#)) OR
 					(reg_q1544 AND symb_decoder(16#17#)) OR
 					(reg_q1544 AND symb_decoder(16#94#)) OR
 					(reg_q1544 AND symb_decoder(16#2a#)) OR
 					(reg_q1544 AND symb_decoder(16#0e#)) OR
 					(reg_q1544 AND symb_decoder(16#82#)) OR
 					(reg_q1544 AND symb_decoder(16#6d#)) OR
 					(reg_q1544 AND symb_decoder(16#f9#)) OR
 					(reg_q1544 AND symb_decoder(16#22#)) OR
 					(reg_q1544 AND symb_decoder(16#34#)) OR
 					(reg_q1544 AND symb_decoder(16#64#)) OR
 					(reg_q1544 AND symb_decoder(16#ad#)) OR
 					(reg_q1544 AND symb_decoder(16#ee#)) OR
 					(reg_q1544 AND symb_decoder(16#c3#)) OR
 					(reg_q1544 AND symb_decoder(16#85#)) OR
 					(reg_q1544 AND symb_decoder(16#1d#)) OR
 					(reg_q1544 AND symb_decoder(16#5f#)) OR
 					(reg_q1544 AND symb_decoder(16#63#)) OR
 					(reg_q1544 AND symb_decoder(16#b9#)) OR
 					(reg_q1544 AND symb_decoder(16#29#)) OR
 					(reg_q1544 AND symb_decoder(16#30#)) OR
 					(reg_q1544 AND symb_decoder(16#26#)) OR
 					(reg_q1544 AND symb_decoder(16#c6#)) OR
 					(reg_q1544 AND symb_decoder(16#d8#)) OR
 					(reg_q1544 AND symb_decoder(16#fa#)) OR
 					(reg_q1544 AND symb_decoder(16#c9#)) OR
 					(reg_q1544 AND symb_decoder(16#aa#)) OR
 					(reg_q1544 AND symb_decoder(16#4b#)) OR
 					(reg_q1544 AND symb_decoder(16#f2#)) OR
 					(reg_q1544 AND symb_decoder(16#6a#)) OR
 					(reg_q1544 AND symb_decoder(16#c8#)) OR
 					(reg_q1544 AND symb_decoder(16#51#)) OR
 					(reg_q1544 AND symb_decoder(16#1f#)) OR
 					(reg_q1544 AND symb_decoder(16#a0#)) OR
 					(reg_q1544 AND symb_decoder(16#77#)) OR
 					(reg_q1544 AND symb_decoder(16#08#)) OR
 					(reg_q1544 AND symb_decoder(16#70#)) OR
 					(reg_q1544 AND symb_decoder(16#7c#)) OR
 					(reg_q1544 AND symb_decoder(16#99#)) OR
 					(reg_q1544 AND symb_decoder(16#69#)) OR
 					(reg_q1544 AND symb_decoder(16#c4#)) OR
 					(reg_q1544 AND symb_decoder(16#ea#)) OR
 					(reg_q1544 AND symb_decoder(16#74#)) OR
 					(reg_q1544 AND symb_decoder(16#1a#)) OR
 					(reg_q1544 AND symb_decoder(16#c7#)) OR
 					(reg_q1544 AND symb_decoder(16#d2#)) OR
 					(reg_q1544 AND symb_decoder(16#76#)) OR
 					(reg_q1544 AND symb_decoder(16#7a#)) OR
 					(reg_q1544 AND symb_decoder(16#bc#)) OR
 					(reg_q1544 AND symb_decoder(16#fb#)) OR
 					(reg_q1544 AND symb_decoder(16#4e#)) OR
 					(reg_q1544 AND symb_decoder(16#87#)) OR
 					(reg_q1544 AND symb_decoder(16#61#)) OR
 					(reg_q1544 AND symb_decoder(16#18#)) OR
 					(reg_q1544 AND symb_decoder(16#5e#)) OR
 					(reg_q1544 AND symb_decoder(16#37#)) OR
 					(reg_q1544 AND symb_decoder(16#ff#)) OR
 					(reg_q1544 AND symb_decoder(16#0f#)) OR
 					(reg_q1544 AND symb_decoder(16#36#)) OR
 					(reg_q1544 AND symb_decoder(16#a6#)) OR
 					(reg_q1544 AND symb_decoder(16#67#)) OR
 					(reg_q1544 AND symb_decoder(16#81#)) OR
 					(reg_q1544 AND symb_decoder(16#15#)) OR
 					(reg_q1544 AND symb_decoder(16#43#)) OR
 					(reg_q1544 AND symb_decoder(16#0c#)) OR
 					(reg_q1544 AND symb_decoder(16#80#)) OR
 					(reg_q1544 AND symb_decoder(16#0d#)) OR
 					(reg_q1544 AND symb_decoder(16#0b#)) OR
 					(reg_q1544 AND symb_decoder(16#89#)) OR
 					(reg_q1544 AND symb_decoder(16#b6#)) OR
 					(reg_q1544 AND symb_decoder(16#9c#)) OR
 					(reg_q1544 AND symb_decoder(16#f4#)) OR
 					(reg_q1544 AND symb_decoder(16#91#)) OR
 					(reg_q1544 AND symb_decoder(16#13#)) OR
 					(reg_q1544 AND symb_decoder(16#e7#)) OR
 					(reg_q1544 AND symb_decoder(16#e6#)) OR
 					(reg_q1544 AND symb_decoder(16#02#)) OR
 					(reg_q1544 AND symb_decoder(16#ec#)) OR
 					(reg_q1544 AND symb_decoder(16#7b#)) OR
 					(reg_q1544 AND symb_decoder(16#cf#)) OR
 					(reg_q1544 AND symb_decoder(16#db#)) OR
 					(reg_q1544 AND symb_decoder(16#d9#)) OR
 					(reg_q1544 AND symb_decoder(16#12#)) OR
 					(reg_q1544 AND symb_decoder(16#84#)) OR
 					(reg_q1544 AND symb_decoder(16#2f#)) OR
 					(reg_q1544 AND symb_decoder(16#9f#)) OR
 					(reg_q1544 AND symb_decoder(16#9b#)) OR
 					(reg_q1544 AND symb_decoder(16#eb#)) OR
 					(reg_q1544 AND symb_decoder(16#28#)) OR
 					(reg_q1544 AND symb_decoder(16#cd#)) OR
 					(reg_q1544 AND symb_decoder(16#54#)) OR
 					(reg_q1544 AND symb_decoder(16#fc#)) OR
 					(reg_q1544 AND symb_decoder(16#a7#)) OR
 					(reg_q1544 AND symb_decoder(16#3e#)) OR
 					(reg_q1544 AND symb_decoder(16#b4#)) OR
 					(reg_q1544 AND symb_decoder(16#e5#)) OR
 					(reg_q1544 AND symb_decoder(16#49#)) OR
 					(reg_q1544 AND symb_decoder(16#2e#)) OR
 					(reg_q1544 AND symb_decoder(16#55#)) OR
 					(reg_q1544 AND symb_decoder(16#45#)) OR
 					(reg_q1544 AND symb_decoder(16#6c#)) OR
 					(reg_q1544 AND symb_decoder(16#d6#)) OR
 					(reg_q1544 AND symb_decoder(16#3d#)) OR
 					(reg_q1544 AND symb_decoder(16#1e#)) OR
 					(reg_q1544 AND symb_decoder(16#90#)) OR
 					(reg_q1544 AND symb_decoder(16#c2#)) OR
 					(reg_q1544 AND symb_decoder(16#21#)) OR
 					(reg_q1544 AND symb_decoder(16#42#)) OR
 					(reg_q1544 AND symb_decoder(16#50#)) OR
 					(reg_q1544 AND symb_decoder(16#b0#)) OR
 					(reg_q1544 AND symb_decoder(16#d4#)) OR
 					(reg_q1544 AND symb_decoder(16#b5#)) OR
 					(reg_q1544 AND symb_decoder(16#71#)) OR
 					(reg_q1544 AND symb_decoder(16#9e#)) OR
 					(reg_q1544 AND symb_decoder(16#20#)) OR
 					(reg_q1544 AND symb_decoder(16#7d#)) OR
 					(reg_q1544 AND symb_decoder(16#b7#)) OR
 					(reg_q1544 AND symb_decoder(16#03#)) OR
 					(reg_q1544 AND symb_decoder(16#86#)) OR
 					(reg_q1544 AND symb_decoder(16#24#)) OR
 					(reg_q1544 AND symb_decoder(16#e4#)) OR
 					(reg_q1544 AND symb_decoder(16#e1#)) OR
 					(reg_q1544 AND symb_decoder(16#f8#)) OR
 					(reg_q1544 AND symb_decoder(16#d1#)) OR
 					(reg_q1544 AND symb_decoder(16#e3#)) OR
 					(reg_q1544 AND symb_decoder(16#bd#)) OR
 					(reg_q1544 AND symb_decoder(16#4d#)) OR
 					(reg_q1544 AND symb_decoder(16#a9#)) OR
 					(reg_q1544 AND symb_decoder(16#c0#)) OR
 					(reg_q1544 AND symb_decoder(16#a1#)) OR
 					(reg_q1544 AND symb_decoder(16#33#)) OR
 					(reg_q1544 AND symb_decoder(16#07#)) OR
 					(reg_q1544 AND symb_decoder(16#af#)) OR
 					(reg_q1544 AND symb_decoder(16#f5#)) OR
 					(reg_q1544 AND symb_decoder(16#cb#)) OR
 					(reg_q1544 AND symb_decoder(16#14#)) OR
 					(reg_q1544 AND symb_decoder(16#16#)) OR
 					(reg_q1544 AND symb_decoder(16#a4#)) OR
 					(reg_q1544 AND symb_decoder(16#4c#)) OR
 					(reg_q1544 AND symb_decoder(16#46#)) OR
 					(reg_q1544 AND symb_decoder(16#65#)) OR
 					(reg_q1544 AND symb_decoder(16#d5#)) OR
 					(reg_q1544 AND symb_decoder(16#0a#)) OR
 					(reg_q1544 AND symb_decoder(16#56#)) OR
 					(reg_q1544 AND symb_decoder(16#5c#)) OR
 					(reg_q1544 AND symb_decoder(16#da#)) OR
 					(reg_q1544 AND symb_decoder(16#f0#)) OR
 					(reg_q1544 AND symb_decoder(16#01#)) OR
 					(reg_q1544 AND symb_decoder(16#04#)) OR
 					(reg_q1544 AND symb_decoder(16#6f#)) OR
 					(reg_q1544 AND symb_decoder(16#31#)) OR
 					(reg_q1544 AND symb_decoder(16#5b#)) OR
 					(reg_q1544 AND symb_decoder(16#3a#)) OR
 					(reg_q1544 AND symb_decoder(16#40#)) OR
 					(reg_q1544 AND symb_decoder(16#93#)) OR
 					(reg_q1544 AND symb_decoder(16#ed#)) OR
 					(reg_q1544 AND symb_decoder(16#32#)) OR
 					(reg_q1544 AND symb_decoder(16#be#)) OR
 					(reg_q1544 AND symb_decoder(16#97#)) OR
 					(reg_q1544 AND symb_decoder(16#a3#)) OR
 					(reg_q1544 AND symb_decoder(16#73#)) OR
 					(reg_q1544 AND symb_decoder(16#de#)) OR
 					(reg_q1544 AND symb_decoder(16#ac#)) OR
 					(reg_q1544 AND symb_decoder(16#62#)) OR
 					(reg_q1544 AND symb_decoder(16#52#)) OR
 					(reg_q1544 AND symb_decoder(16#39#)) OR
 					(reg_q1544 AND symb_decoder(16#09#)) OR
 					(reg_q1544 AND symb_decoder(16#fe#)) OR
 					(reg_q1544 AND symb_decoder(16#00#)) OR
 					(reg_q1544 AND symb_decoder(16#5a#)) OR
 					(reg_q1544 AND symb_decoder(16#59#)) OR
 					(reg_q1544 AND symb_decoder(16#05#)) OR
 					(reg_q1544 AND symb_decoder(16#9a#)) OR
 					(reg_q1544 AND symb_decoder(16#e8#)) OR
 					(reg_q1544 AND symb_decoder(16#23#)) OR
 					(reg_q1544 AND symb_decoder(16#57#)) OR
 					(reg_q1544 AND symb_decoder(16#47#)) OR
 					(reg_q1544 AND symb_decoder(16#96#)) OR
 					(reg_q1544 AND symb_decoder(16#8e#)) OR
 					(reg_q1544 AND symb_decoder(16#95#)) OR
 					(reg_q1544 AND symb_decoder(16#ce#)) OR
 					(reg_q1544 AND symb_decoder(16#60#)) OR
 					(reg_q1544 AND symb_decoder(16#f6#)) OR
 					(reg_q1544 AND symb_decoder(16#b8#)) OR
 					(reg_q1544 AND symb_decoder(16#ab#)) OR
 					(reg_q1544 AND symb_decoder(16#a5#)) OR
 					(reg_q1544 AND symb_decoder(16#35#)) OR
 					(reg_q1544 AND symb_decoder(16#7e#)) OR
 					(reg_q1544 AND symb_decoder(16#8f#)) OR
 					(reg_q1544 AND symb_decoder(16#b1#)) OR
 					(reg_q1544 AND symb_decoder(16#92#)) OR
 					(reg_q1544 AND symb_decoder(16#8c#)) OR
 					(reg_q1544 AND symb_decoder(16#6e#)) OR
 					(reg_q1544 AND symb_decoder(16#c5#)) OR
 					(reg_q1544 AND symb_decoder(16#ae#)) OR
 					(reg_q1544 AND symb_decoder(16#72#)) OR
 					(reg_q1544 AND symb_decoder(16#10#)) OR
 					(reg_q1544 AND symb_decoder(16#bf#)) OR
 					(reg_q1544 AND symb_decoder(16#d3#)) OR
 					(reg_q1544 AND symb_decoder(16#ca#)) OR
 					(reg_q1544 AND symb_decoder(16#78#)) OR
 					(reg_q1544 AND symb_decoder(16#8d#)) OR
 					(reg_q1544 AND symb_decoder(16#e9#)) OR
 					(reg_q1544 AND symb_decoder(16#83#)) OR
 					(reg_q1544 AND symb_decoder(16#ef#)) OR
 					(reg_q1544 AND symb_decoder(16#2d#)) OR
 					(reg_q1544 AND symb_decoder(16#19#)) OR
 					(reg_q1544 AND symb_decoder(16#c1#)) OR
 					(reg_q1544 AND symb_decoder(16#44#)) OR
 					(reg_q1544 AND symb_decoder(16#f7#)) OR
 					(reg_q1544 AND symb_decoder(16#88#)) OR
 					(reg_q1544 AND symb_decoder(16#3c#)) OR
 					(reg_q1544 AND symb_decoder(16#d0#)) OR
 					(reg_q1544 AND symb_decoder(16#53#)) OR
 					(reg_q1544 AND symb_decoder(16#f1#)) OR
 					(reg_q1544 AND symb_decoder(16#dc#)) OR
 					(reg_q1544 AND symb_decoder(16#1b#)) OR
 					(reg_q1544 AND symb_decoder(16#25#)) OR
 					(reg_q1544 AND symb_decoder(16#4a#)) OR
 					(reg_q1544 AND symb_decoder(16#b2#)) OR
 					(reg_q1544 AND symb_decoder(16#df#)) OR
 					(reg_q1544 AND symb_decoder(16#58#)) OR
 					(reg_q1544 AND symb_decoder(16#b3#)) OR
 					(reg_q1544 AND symb_decoder(16#fd#)) OR
 					(reg_q1544 AND symb_decoder(16#1c#)) OR
 					(reg_q1544 AND symb_decoder(16#a2#)) OR
 					(reg_q1544 AND symb_decoder(16#8a#)) OR
 					(reg_q1544 AND symb_decoder(16#9d#)) OR
 					(reg_q1544 AND symb_decoder(16#3f#)) OR
 					(reg_q1544 AND symb_decoder(16#8b#)) OR
 					(reg_q1544 AND symb_decoder(16#cc#)) OR
 					(reg_q1544 AND symb_decoder(16#98#)) OR
 					(reg_q1544 AND symb_decoder(16#dd#)) OR
 					(reg_q1544 AND symb_decoder(16#bb#)) OR
 					(reg_q1544 AND symb_decoder(16#2b#)) OR
 					(reg_q1544 AND symb_decoder(16#79#)) OR
 					(reg_q1544 AND symb_decoder(16#41#)) OR
 					(reg_q1544 AND symb_decoder(16#38#)) OR
 					(reg_q1544 AND symb_decoder(16#2c#)) OR
 					(reg_q1544 AND symb_decoder(16#06#)) OR
 					(reg_q1544 AND symb_decoder(16#e0#)) OR
 					(reg_q1544 AND symb_decoder(16#11#)) OR
 					(reg_q1544 AND symb_decoder(16#a8#)) OR
 					(reg_q1544 AND symb_decoder(16#f3#)) OR
 					(reg_q1544 AND symb_decoder(16#66#)) OR
 					(reg_q1544 AND symb_decoder(16#68#)) OR
 					(reg_q1544 AND symb_decoder(16#7f#)) OR
 					(reg_q1544 AND symb_decoder(16#5d#));
reg_q1544_init <= '0' ;
	p_reg_q1544: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1544 <= reg_q1544_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1544 <= reg_q1544_init;
        else
          reg_q1544 <= reg_q1544_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2208_in <= (reg_q2172 AND symb_decoder(16#df#)) OR
 					(reg_q2172 AND symb_decoder(16#b4#)) OR
 					(reg_q2172 AND symb_decoder(16#9d#)) OR
 					(reg_q2172 AND symb_decoder(16#3f#)) OR
 					(reg_q2172 AND symb_decoder(16#64#)) OR
 					(reg_q2172 AND symb_decoder(16#2f#)) OR
 					(reg_q2172 AND symb_decoder(16#0f#)) OR
 					(reg_q2172 AND symb_decoder(16#31#)) OR
 					(reg_q2172 AND symb_decoder(16#8f#)) OR
 					(reg_q2172 AND symb_decoder(16#81#)) OR
 					(reg_q2172 AND symb_decoder(16#8e#)) OR
 					(reg_q2172 AND symb_decoder(16#9e#)) OR
 					(reg_q2172 AND symb_decoder(16#04#)) OR
 					(reg_q2172 AND symb_decoder(16#ff#)) OR
 					(reg_q2172 AND symb_decoder(16#4b#)) OR
 					(reg_q2172 AND symb_decoder(16#46#)) OR
 					(reg_q2172 AND symb_decoder(16#f4#)) OR
 					(reg_q2172 AND symb_decoder(16#0b#)) OR
 					(reg_q2172 AND symb_decoder(16#09#)) OR
 					(reg_q2172 AND symb_decoder(16#e1#)) OR
 					(reg_q2172 AND symb_decoder(16#9f#)) OR
 					(reg_q2172 AND symb_decoder(16#58#)) OR
 					(reg_q2172 AND symb_decoder(16#ae#)) OR
 					(reg_q2172 AND symb_decoder(16#be#)) OR
 					(reg_q2172 AND symb_decoder(16#a0#)) OR
 					(reg_q2172 AND symb_decoder(16#d3#)) OR
 					(reg_q2172 AND symb_decoder(16#84#)) OR
 					(reg_q2172 AND symb_decoder(16#97#)) OR
 					(reg_q2172 AND symb_decoder(16#36#)) OR
 					(reg_q2172 AND symb_decoder(16#e0#)) OR
 					(reg_q2172 AND symb_decoder(16#99#)) OR
 					(reg_q2172 AND symb_decoder(16#96#)) OR
 					(reg_q2172 AND symb_decoder(16#bd#)) OR
 					(reg_q2172 AND symb_decoder(16#63#)) OR
 					(reg_q2172 AND symb_decoder(16#f8#)) OR
 					(reg_q2172 AND symb_decoder(16#c9#)) OR
 					(reg_q2172 AND symb_decoder(16#b2#)) OR
 					(reg_q2172 AND symb_decoder(16#b8#)) OR
 					(reg_q2172 AND symb_decoder(16#af#)) OR
 					(reg_q2172 AND symb_decoder(16#88#)) OR
 					(reg_q2172 AND symb_decoder(16#5c#)) OR
 					(reg_q2172 AND symb_decoder(16#ea#)) OR
 					(reg_q2172 AND symb_decoder(16#56#)) OR
 					(reg_q2172 AND symb_decoder(16#2b#)) OR
 					(reg_q2172 AND symb_decoder(16#5b#)) OR
 					(reg_q2172 AND symb_decoder(16#7d#)) OR
 					(reg_q2172 AND symb_decoder(16#07#)) OR
 					(reg_q2172 AND symb_decoder(16#bf#)) OR
 					(reg_q2172 AND symb_decoder(16#dc#)) OR
 					(reg_q2172 AND symb_decoder(16#c6#)) OR
 					(reg_q2172 AND symb_decoder(16#76#)) OR
 					(reg_q2172 AND symb_decoder(16#23#)) OR
 					(reg_q2172 AND symb_decoder(16#90#)) OR
 					(reg_q2172 AND symb_decoder(16#a8#)) OR
 					(reg_q2172 AND symb_decoder(16#39#)) OR
 					(reg_q2172 AND symb_decoder(16#05#)) OR
 					(reg_q2172 AND symb_decoder(16#ca#)) OR
 					(reg_q2172 AND symb_decoder(16#26#)) OR
 					(reg_q2172 AND symb_decoder(16#c5#)) OR
 					(reg_q2172 AND symb_decoder(16#89#)) OR
 					(reg_q2172 AND symb_decoder(16#e6#)) OR
 					(reg_q2172 AND symb_decoder(16#2d#)) OR
 					(reg_q2172 AND symb_decoder(16#b1#)) OR
 					(reg_q2172 AND symb_decoder(16#74#)) OR
 					(reg_q2172 AND symb_decoder(16#e9#)) OR
 					(reg_q2172 AND symb_decoder(16#37#)) OR
 					(reg_q2172 AND symb_decoder(16#f2#)) OR
 					(reg_q2172 AND symb_decoder(16#b9#)) OR
 					(reg_q2172 AND symb_decoder(16#8c#)) OR
 					(reg_q2172 AND symb_decoder(16#cc#)) OR
 					(reg_q2172 AND symb_decoder(16#ed#)) OR
 					(reg_q2172 AND symb_decoder(16#ba#)) OR
 					(reg_q2172 AND symb_decoder(16#17#)) OR
 					(reg_q2172 AND symb_decoder(16#dd#)) OR
 					(reg_q2172 AND symb_decoder(16#3e#)) OR
 					(reg_q2172 AND symb_decoder(16#19#)) OR
 					(reg_q2172 AND symb_decoder(16#6d#)) OR
 					(reg_q2172 AND symb_decoder(16#5a#)) OR
 					(reg_q2172 AND symb_decoder(16#22#)) OR
 					(reg_q2172 AND symb_decoder(16#68#)) OR
 					(reg_q2172 AND symb_decoder(16#3c#)) OR
 					(reg_q2172 AND symb_decoder(16#f9#)) OR
 					(reg_q2172 AND symb_decoder(16#a4#)) OR
 					(reg_q2172 AND symb_decoder(16#4a#)) OR
 					(reg_q2172 AND symb_decoder(16#eb#)) OR
 					(reg_q2172 AND symb_decoder(16#fd#)) OR
 					(reg_q2172 AND symb_decoder(16#d6#)) OR
 					(reg_q2172 AND symb_decoder(16#86#)) OR
 					(reg_q2172 AND symb_decoder(16#ce#)) OR
 					(reg_q2172 AND symb_decoder(16#03#)) OR
 					(reg_q2172 AND symb_decoder(16#00#)) OR
 					(reg_q2172 AND symb_decoder(16#95#)) OR
 					(reg_q2172 AND symb_decoder(16#d9#)) OR
 					(reg_q2172 AND symb_decoder(16#3a#)) OR
 					(reg_q2172 AND symb_decoder(16#b0#)) OR
 					(reg_q2172 AND symb_decoder(16#35#)) OR
 					(reg_q2172 AND symb_decoder(16#2c#)) OR
 					(reg_q2172 AND symb_decoder(16#45#)) OR
 					(reg_q2172 AND symb_decoder(16#cf#)) OR
 					(reg_q2172 AND symb_decoder(16#59#)) OR
 					(reg_q2172 AND symb_decoder(16#28#)) OR
 					(reg_q2172 AND symb_decoder(16#71#)) OR
 					(reg_q2172 AND symb_decoder(16#0d#)) OR
 					(reg_q2172 AND symb_decoder(16#80#)) OR
 					(reg_q2172 AND symb_decoder(16#d2#)) OR
 					(reg_q2172 AND symb_decoder(16#bc#)) OR
 					(reg_q2172 AND symb_decoder(16#6f#)) OR
 					(reg_q2172 AND symb_decoder(16#8b#)) OR
 					(reg_q2172 AND symb_decoder(16#3b#)) OR
 					(reg_q2172 AND symb_decoder(16#02#)) OR
 					(reg_q2172 AND symb_decoder(16#1f#)) OR
 					(reg_q2172 AND symb_decoder(16#5f#)) OR
 					(reg_q2172 AND symb_decoder(16#3d#)) OR
 					(reg_q2172 AND symb_decoder(16#a7#)) OR
 					(reg_q2172 AND symb_decoder(16#b3#)) OR
 					(reg_q2172 AND symb_decoder(16#a2#)) OR
 					(reg_q2172 AND symb_decoder(16#67#)) OR
 					(reg_q2172 AND symb_decoder(16#25#)) OR
 					(reg_q2172 AND symb_decoder(16#53#)) OR
 					(reg_q2172 AND symb_decoder(16#b6#)) OR
 					(reg_q2172 AND symb_decoder(16#41#)) OR
 					(reg_q2172 AND symb_decoder(16#92#)) OR
 					(reg_q2172 AND symb_decoder(16#54#)) OR
 					(reg_q2172 AND symb_decoder(16#cd#)) OR
 					(reg_q2172 AND symb_decoder(16#f5#)) OR
 					(reg_q2172 AND symb_decoder(16#2e#)) OR
 					(reg_q2172 AND symb_decoder(16#18#)) OR
 					(reg_q2172 AND symb_decoder(16#52#)) OR
 					(reg_q2172 AND symb_decoder(16#ec#)) OR
 					(reg_q2172 AND symb_decoder(16#30#)) OR
 					(reg_q2172 AND symb_decoder(16#f6#)) OR
 					(reg_q2172 AND symb_decoder(16#d8#)) OR
 					(reg_q2172 AND symb_decoder(16#7f#)) OR
 					(reg_q2172 AND symb_decoder(16#91#)) OR
 					(reg_q2172 AND symb_decoder(16#0c#)) OR
 					(reg_q2172 AND symb_decoder(16#20#)) OR
 					(reg_q2172 AND symb_decoder(16#de#)) OR
 					(reg_q2172 AND symb_decoder(16#aa#)) OR
 					(reg_q2172 AND symb_decoder(16#cb#)) OR
 					(reg_q2172 AND symb_decoder(16#87#)) OR
 					(reg_q2172 AND symb_decoder(16#7e#)) OR
 					(reg_q2172 AND symb_decoder(16#d7#)) OR
 					(reg_q2172 AND symb_decoder(16#c4#)) OR
 					(reg_q2172 AND symb_decoder(16#49#)) OR
 					(reg_q2172 AND symb_decoder(16#85#)) OR
 					(reg_q2172 AND symb_decoder(16#da#)) OR
 					(reg_q2172 AND symb_decoder(16#33#)) OR
 					(reg_q2172 AND symb_decoder(16#34#)) OR
 					(reg_q2172 AND symb_decoder(16#47#)) OR
 					(reg_q2172 AND symb_decoder(16#48#)) OR
 					(reg_q2172 AND symb_decoder(16#a1#)) OR
 					(reg_q2172 AND symb_decoder(16#75#)) OR
 					(reg_q2172 AND symb_decoder(16#27#)) OR
 					(reg_q2172 AND symb_decoder(16#12#)) OR
 					(reg_q2172 AND symb_decoder(16#78#)) OR
 					(reg_q2172 AND symb_decoder(16#1b#)) OR
 					(reg_q2172 AND symb_decoder(16#e8#)) OR
 					(reg_q2172 AND symb_decoder(16#d5#)) OR
 					(reg_q2172 AND symb_decoder(16#e7#)) OR
 					(reg_q2172 AND symb_decoder(16#0a#)) OR
 					(reg_q2172 AND symb_decoder(16#5d#)) OR
 					(reg_q2172 AND symb_decoder(16#44#)) OR
 					(reg_q2172 AND symb_decoder(16#06#)) OR
 					(reg_q2172 AND symb_decoder(16#40#)) OR
 					(reg_q2172 AND symb_decoder(16#1c#)) OR
 					(reg_q2172 AND symb_decoder(16#32#)) OR
 					(reg_q2172 AND symb_decoder(16#9a#)) OR
 					(reg_q2172 AND symb_decoder(16#e3#)) OR
 					(reg_q2172 AND symb_decoder(16#e2#)) OR
 					(reg_q2172 AND symb_decoder(16#69#)) OR
 					(reg_q2172 AND symb_decoder(16#6b#)) OR
 					(reg_q2172 AND symb_decoder(16#e4#)) OR
 					(reg_q2172 AND symb_decoder(16#0e#)) OR
 					(reg_q2172 AND symb_decoder(16#8a#)) OR
 					(reg_q2172 AND symb_decoder(16#d4#)) OR
 					(reg_q2172 AND symb_decoder(16#a9#)) OR
 					(reg_q2172 AND symb_decoder(16#b5#)) OR
 					(reg_q2172 AND symb_decoder(16#f3#)) OR
 					(reg_q2172 AND symb_decoder(16#9c#)) OR
 					(reg_q2172 AND symb_decoder(16#77#)) OR
 					(reg_q2172 AND symb_decoder(16#50#)) OR
 					(reg_q2172 AND symb_decoder(16#66#)) OR
 					(reg_q2172 AND symb_decoder(16#fb#)) OR
 					(reg_q2172 AND symb_decoder(16#ee#)) OR
 					(reg_q2172 AND symb_decoder(16#ab#)) OR
 					(reg_q2172 AND symb_decoder(16#bb#)) OR
 					(reg_q2172 AND symb_decoder(16#08#)) OR
 					(reg_q2172 AND symb_decoder(16#6c#)) OR
 					(reg_q2172 AND symb_decoder(16#14#)) OR
 					(reg_q2172 AND symb_decoder(16#c2#)) OR
 					(reg_q2172 AND symb_decoder(16#7c#)) OR
 					(reg_q2172 AND symb_decoder(16#15#)) OR
 					(reg_q2172 AND symb_decoder(16#4f#)) OR
 					(reg_q2172 AND symb_decoder(16#01#)) OR
 					(reg_q2172 AND symb_decoder(16#4e#)) OR
 					(reg_q2172 AND symb_decoder(16#93#)) OR
 					(reg_q2172 AND symb_decoder(16#21#)) OR
 					(reg_q2172 AND symb_decoder(16#c3#)) OR
 					(reg_q2172 AND symb_decoder(16#1e#)) OR
 					(reg_q2172 AND symb_decoder(16#4d#)) OR
 					(reg_q2172 AND symb_decoder(16#ac#)) OR
 					(reg_q2172 AND symb_decoder(16#16#)) OR
 					(reg_q2172 AND symb_decoder(16#a3#)) OR
 					(reg_q2172 AND symb_decoder(16#fe#)) OR
 					(reg_q2172 AND symb_decoder(16#42#)) OR
 					(reg_q2172 AND symb_decoder(16#13#)) OR
 					(reg_q2172 AND symb_decoder(16#ad#)) OR
 					(reg_q2172 AND symb_decoder(16#7b#)) OR
 					(reg_q2172 AND symb_decoder(16#a6#)) OR
 					(reg_q2172 AND symb_decoder(16#d1#)) OR
 					(reg_q2172 AND symb_decoder(16#62#)) OR
 					(reg_q2172 AND symb_decoder(16#9b#)) OR
 					(reg_q2172 AND symb_decoder(16#2a#)) OR
 					(reg_q2172 AND symb_decoder(16#65#)) OR
 					(reg_q2172 AND symb_decoder(16#10#)) OR
 					(reg_q2172 AND symb_decoder(16#a5#)) OR
 					(reg_q2172 AND symb_decoder(16#5e#)) OR
 					(reg_q2172 AND symb_decoder(16#d0#)) OR
 					(reg_q2172 AND symb_decoder(16#6a#)) OR
 					(reg_q2172 AND symb_decoder(16#c7#)) OR
 					(reg_q2172 AND symb_decoder(16#29#)) OR
 					(reg_q2172 AND symb_decoder(16#38#)) OR
 					(reg_q2172 AND symb_decoder(16#f0#)) OR
 					(reg_q2172 AND symb_decoder(16#43#)) OR
 					(reg_q2172 AND symb_decoder(16#94#)) OR
 					(reg_q2172 AND symb_decoder(16#70#)) OR
 					(reg_q2172 AND symb_decoder(16#8d#)) OR
 					(reg_q2172 AND symb_decoder(16#57#)) OR
 					(reg_q2172 AND symb_decoder(16#fc#)) OR
 					(reg_q2172 AND symb_decoder(16#1a#)) OR
 					(reg_q2172 AND symb_decoder(16#72#)) OR
 					(reg_q2172 AND symb_decoder(16#fa#)) OR
 					(reg_q2172 AND symb_decoder(16#4c#)) OR
 					(reg_q2172 AND symb_decoder(16#60#)) OR
 					(reg_q2172 AND symb_decoder(16#c8#)) OR
 					(reg_q2172 AND symb_decoder(16#98#)) OR
 					(reg_q2172 AND symb_decoder(16#f7#)) OR
 					(reg_q2172 AND symb_decoder(16#83#)) OR
 					(reg_q2172 AND symb_decoder(16#6e#)) OR
 					(reg_q2172 AND symb_decoder(16#51#)) OR
 					(reg_q2172 AND symb_decoder(16#55#)) OR
 					(reg_q2172 AND symb_decoder(16#c0#)) OR
 					(reg_q2172 AND symb_decoder(16#11#)) OR
 					(reg_q2172 AND symb_decoder(16#79#)) OR
 					(reg_q2172 AND symb_decoder(16#ef#)) OR
 					(reg_q2172 AND symb_decoder(16#24#)) OR
 					(reg_q2172 AND symb_decoder(16#b7#)) OR
 					(reg_q2172 AND symb_decoder(16#73#)) OR
 					(reg_q2172 AND symb_decoder(16#82#)) OR
 					(reg_q2172 AND symb_decoder(16#e5#)) OR
 					(reg_q2172 AND symb_decoder(16#c1#)) OR
 					(reg_q2172 AND symb_decoder(16#61#)) OR
 					(reg_q2172 AND symb_decoder(16#db#)) OR
 					(reg_q2172 AND symb_decoder(16#7a#)) OR
 					(reg_q2172 AND symb_decoder(16#1d#)) OR
 					(reg_q2172 AND symb_decoder(16#f1#)) OR
 					(reg_q2208 AND symb_decoder(16#db#)) OR
 					(reg_q2208 AND symb_decoder(16#7a#)) OR
 					(reg_q2208 AND symb_decoder(16#2a#)) OR
 					(reg_q2208 AND symb_decoder(16#9a#)) OR
 					(reg_q2208 AND symb_decoder(16#99#)) OR
 					(reg_q2208 AND symb_decoder(16#8d#)) OR
 					(reg_q2208 AND symb_decoder(16#59#)) OR
 					(reg_q2208 AND symb_decoder(16#54#)) OR
 					(reg_q2208 AND symb_decoder(16#cd#)) OR
 					(reg_q2208 AND symb_decoder(16#34#)) OR
 					(reg_q2208 AND symb_decoder(16#41#)) OR
 					(reg_q2208 AND symb_decoder(16#7f#)) OR
 					(reg_q2208 AND symb_decoder(16#d2#)) OR
 					(reg_q2208 AND symb_decoder(16#e9#)) OR
 					(reg_q2208 AND symb_decoder(16#d3#)) OR
 					(reg_q2208 AND symb_decoder(16#21#)) OR
 					(reg_q2208 AND symb_decoder(16#e3#)) OR
 					(reg_q2208 AND symb_decoder(16#16#)) OR
 					(reg_q2208 AND symb_decoder(16#c8#)) OR
 					(reg_q2208 AND symb_decoder(16#56#)) OR
 					(reg_q2208 AND symb_decoder(16#72#)) OR
 					(reg_q2208 AND symb_decoder(16#95#)) OR
 					(reg_q2208 AND symb_decoder(16#2f#)) OR
 					(reg_q2208 AND symb_decoder(16#3c#)) OR
 					(reg_q2208 AND symb_decoder(16#fe#)) OR
 					(reg_q2208 AND symb_decoder(16#6a#)) OR
 					(reg_q2208 AND symb_decoder(16#73#)) OR
 					(reg_q2208 AND symb_decoder(16#61#)) OR
 					(reg_q2208 AND symb_decoder(16#b5#)) OR
 					(reg_q2208 AND symb_decoder(16#7c#)) OR
 					(reg_q2208 AND symb_decoder(16#27#)) OR
 					(reg_q2208 AND symb_decoder(16#44#)) OR
 					(reg_q2208 AND symb_decoder(16#b0#)) OR
 					(reg_q2208 AND symb_decoder(16#04#)) OR
 					(reg_q2208 AND symb_decoder(16#eb#)) OR
 					(reg_q2208 AND symb_decoder(16#6d#)) OR
 					(reg_q2208 AND symb_decoder(16#92#)) OR
 					(reg_q2208 AND symb_decoder(16#7d#)) OR
 					(reg_q2208 AND symb_decoder(16#15#)) OR
 					(reg_q2208 AND symb_decoder(16#12#)) OR
 					(reg_q2208 AND symb_decoder(16#13#)) OR
 					(reg_q2208 AND symb_decoder(16#ed#)) OR
 					(reg_q2208 AND symb_decoder(16#00#)) OR
 					(reg_q2208 AND symb_decoder(16#ca#)) OR
 					(reg_q2208 AND symb_decoder(16#7e#)) OR
 					(reg_q2208 AND symb_decoder(16#2d#)) OR
 					(reg_q2208 AND symb_decoder(16#69#)) OR
 					(reg_q2208 AND symb_decoder(16#e7#)) OR
 					(reg_q2208 AND symb_decoder(16#85#)) OR
 					(reg_q2208 AND symb_decoder(16#f2#)) OR
 					(reg_q2208 AND symb_decoder(16#a9#)) OR
 					(reg_q2208 AND symb_decoder(16#55#)) OR
 					(reg_q2208 AND symb_decoder(16#c0#)) OR
 					(reg_q2208 AND symb_decoder(16#71#)) OR
 					(reg_q2208 AND symb_decoder(16#0a#)) OR
 					(reg_q2208 AND symb_decoder(16#4c#)) OR
 					(reg_q2208 AND symb_decoder(16#bc#)) OR
 					(reg_q2208 AND symb_decoder(16#77#)) OR
 					(reg_q2208 AND symb_decoder(16#45#)) OR
 					(reg_q2208 AND symb_decoder(16#d6#)) OR
 					(reg_q2208 AND symb_decoder(16#10#)) OR
 					(reg_q2208 AND symb_decoder(16#d4#)) OR
 					(reg_q2208 AND symb_decoder(16#b2#)) OR
 					(reg_q2208 AND symb_decoder(16#f6#)) OR
 					(reg_q2208 AND symb_decoder(16#ff#)) OR
 					(reg_q2208 AND symb_decoder(16#93#)) OR
 					(reg_q2208 AND symb_decoder(16#5d#)) OR
 					(reg_q2208 AND symb_decoder(16#d9#)) OR
 					(reg_q2208 AND symb_decoder(16#e8#)) OR
 					(reg_q2208 AND symb_decoder(16#fb#)) OR
 					(reg_q2208 AND symb_decoder(16#ea#)) OR
 					(reg_q2208 AND symb_decoder(16#ba#)) OR
 					(reg_q2208 AND symb_decoder(16#83#)) OR
 					(reg_q2208 AND symb_decoder(16#66#)) OR
 					(reg_q2208 AND symb_decoder(16#82#)) OR
 					(reg_q2208 AND symb_decoder(16#30#)) OR
 					(reg_q2208 AND symb_decoder(16#ee#)) OR
 					(reg_q2208 AND symb_decoder(16#f0#)) OR
 					(reg_q2208 AND symb_decoder(16#18#)) OR
 					(reg_q2208 AND symb_decoder(16#52#)) OR
 					(reg_q2208 AND symb_decoder(16#ec#)) OR
 					(reg_q2208 AND symb_decoder(16#ad#)) OR
 					(reg_q2208 AND symb_decoder(16#0c#)) OR
 					(reg_q2208 AND symb_decoder(16#e1#)) OR
 					(reg_q2208 AND symb_decoder(16#31#)) OR
 					(reg_q2208 AND symb_decoder(16#89#)) OR
 					(reg_q2208 AND symb_decoder(16#a2#)) OR
 					(reg_q2208 AND symb_decoder(16#b7#)) OR
 					(reg_q2208 AND symb_decoder(16#b1#)) OR
 					(reg_q2208 AND symb_decoder(16#a4#)) OR
 					(reg_q2208 AND symb_decoder(16#29#)) OR
 					(reg_q2208 AND symb_decoder(16#74#)) OR
 					(reg_q2208 AND symb_decoder(16#0b#)) OR
 					(reg_q2208 AND symb_decoder(16#4a#)) OR
 					(reg_q2208 AND symb_decoder(16#9d#)) OR
 					(reg_q2208 AND symb_decoder(16#cc#)) OR
 					(reg_q2208 AND symb_decoder(16#bd#)) OR
 					(reg_q2208 AND symb_decoder(16#60#)) OR
 					(reg_q2208 AND symb_decoder(16#51#)) OR
 					(reg_q2208 AND symb_decoder(16#1c#)) OR
 					(reg_q2208 AND symb_decoder(16#1b#)) OR
 					(reg_q2208 AND symb_decoder(16#6c#)) OR
 					(reg_q2208 AND symb_decoder(16#87#)) OR
 					(reg_q2208 AND symb_decoder(16#09#)) OR
 					(reg_q2208 AND symb_decoder(16#67#)) OR
 					(reg_q2208 AND symb_decoder(16#3a#)) OR
 					(reg_q2208 AND symb_decoder(16#1d#)) OR
 					(reg_q2208 AND symb_decoder(16#e5#)) OR
 					(reg_q2208 AND symb_decoder(16#0d#)) OR
 					(reg_q2208 AND symb_decoder(16#6f#)) OR
 					(reg_q2208 AND symb_decoder(16#36#)) OR
 					(reg_q2208 AND symb_decoder(16#96#)) OR
 					(reg_q2208 AND symb_decoder(16#f8#)) OR
 					(reg_q2208 AND symb_decoder(16#8b#)) OR
 					(reg_q2208 AND symb_decoder(16#79#)) OR
 					(reg_q2208 AND symb_decoder(16#06#)) OR
 					(reg_q2208 AND symb_decoder(16#a3#)) OR
 					(reg_q2208 AND symb_decoder(16#ce#)) OR
 					(reg_q2208 AND symb_decoder(16#ab#)) OR
 					(reg_q2208 AND symb_decoder(16#c9#)) OR
 					(reg_q2208 AND symb_decoder(16#8e#)) OR
 					(reg_q2208 AND symb_decoder(16#94#)) OR
 					(reg_q2208 AND symb_decoder(16#a6#)) OR
 					(reg_q2208 AND symb_decoder(16#e4#)) OR
 					(reg_q2208 AND symb_decoder(16#40#)) OR
 					(reg_q2208 AND symb_decoder(16#c2#)) OR
 					(reg_q2208 AND symb_decoder(16#22#)) OR
 					(reg_q2208 AND symb_decoder(16#a7#)) OR
 					(reg_q2208 AND symb_decoder(16#6e#)) OR
 					(reg_q2208 AND symb_decoder(16#17#)) OR
 					(reg_q2208 AND symb_decoder(16#f1#)) OR
 					(reg_q2208 AND symb_decoder(16#ae#)) OR
 					(reg_q2208 AND symb_decoder(16#4b#)) OR
 					(reg_q2208 AND symb_decoder(16#c5#)) OR
 					(reg_q2208 AND symb_decoder(16#f3#)) OR
 					(reg_q2208 AND symb_decoder(16#50#)) OR
 					(reg_q2208 AND symb_decoder(16#05#)) OR
 					(reg_q2208 AND symb_decoder(16#a1#)) OR
 					(reg_q2208 AND symb_decoder(16#80#)) OR
 					(reg_q2208 AND symb_decoder(16#6b#)) OR
 					(reg_q2208 AND symb_decoder(16#14#)) OR
 					(reg_q2208 AND symb_decoder(16#ef#)) OR
 					(reg_q2208 AND symb_decoder(16#49#)) OR
 					(reg_q2208 AND symb_decoder(16#7b#)) OR
 					(reg_q2208 AND symb_decoder(16#58#)) OR
 					(reg_q2208 AND symb_decoder(16#8a#)) OR
 					(reg_q2208 AND symb_decoder(16#b3#)) OR
 					(reg_q2208 AND symb_decoder(16#68#)) OR
 					(reg_q2208 AND symb_decoder(16#4d#)) OR
 					(reg_q2208 AND symb_decoder(16#f4#)) OR
 					(reg_q2208 AND symb_decoder(16#5a#)) OR
 					(reg_q2208 AND symb_decoder(16#76#)) OR
 					(reg_q2208 AND symb_decoder(16#53#)) OR
 					(reg_q2208 AND symb_decoder(16#2c#)) OR
 					(reg_q2208 AND symb_decoder(16#5e#)) OR
 					(reg_q2208 AND symb_decoder(16#01#)) OR
 					(reg_q2208 AND symb_decoder(16#46#)) OR
 					(reg_q2208 AND symb_decoder(16#d8#)) OR
 					(reg_q2208 AND symb_decoder(16#f9#)) OR
 					(reg_q2208 AND symb_decoder(16#2e#)) OR
 					(reg_q2208 AND symb_decoder(16#2b#)) OR
 					(reg_q2208 AND symb_decoder(16#91#)) OR
 					(reg_q2208 AND symb_decoder(16#0e#)) OR
 					(reg_q2208 AND symb_decoder(16#3f#)) OR
 					(reg_q2208 AND symb_decoder(16#1f#)) OR
 					(reg_q2208 AND symb_decoder(16#86#)) OR
 					(reg_q2208 AND symb_decoder(16#dc#)) OR
 					(reg_q2208 AND symb_decoder(16#97#)) OR
 					(reg_q2208 AND symb_decoder(16#37#)) OR
 					(reg_q2208 AND symb_decoder(16#62#)) OR
 					(reg_q2208 AND symb_decoder(16#d1#)) OR
 					(reg_q2208 AND symb_decoder(16#4f#)) OR
 					(reg_q2208 AND symb_decoder(16#28#)) OR
 					(reg_q2208 AND symb_decoder(16#fd#)) OR
 					(reg_q2208 AND symb_decoder(16#33#)) OR
 					(reg_q2208 AND symb_decoder(16#0f#)) OR
 					(reg_q2208 AND symb_decoder(16#3e#)) OR
 					(reg_q2208 AND symb_decoder(16#25#)) OR
 					(reg_q2208 AND symb_decoder(16#fa#)) OR
 					(reg_q2208 AND symb_decoder(16#98#)) OR
 					(reg_q2208 AND symb_decoder(16#a5#)) OR
 					(reg_q2208 AND symb_decoder(16#75#)) OR
 					(reg_q2208 AND symb_decoder(16#e2#)) OR
 					(reg_q2208 AND symb_decoder(16#64#)) OR
 					(reg_q2208 AND symb_decoder(16#23#)) OR
 					(reg_q2208 AND symb_decoder(16#43#)) OR
 					(reg_q2208 AND symb_decoder(16#b4#)) OR
 					(reg_q2208 AND symb_decoder(16#d7#)) OR
 					(reg_q2208 AND symb_decoder(16#02#)) OR
 					(reg_q2208 AND symb_decoder(16#d0#)) OR
 					(reg_q2208 AND symb_decoder(16#78#)) OR
 					(reg_q2208 AND symb_decoder(16#c4#)) OR
 					(reg_q2208 AND symb_decoder(16#24#)) OR
 					(reg_q2208 AND symb_decoder(16#5b#)) OR
 					(reg_q2208 AND symb_decoder(16#32#)) OR
 					(reg_q2208 AND symb_decoder(16#11#)) OR
 					(reg_q2208 AND symb_decoder(16#65#)) OR
 					(reg_q2208 AND symb_decoder(16#b9#)) OR
 					(reg_q2208 AND symb_decoder(16#ac#)) OR
 					(reg_q2208 AND symb_decoder(16#26#)) OR
 					(reg_q2208 AND symb_decoder(16#8f#)) OR
 					(reg_q2208 AND symb_decoder(16#42#)) OR
 					(reg_q2208 AND symb_decoder(16#f5#)) OR
 					(reg_q2208 AND symb_decoder(16#9b#)) OR
 					(reg_q2208 AND symb_decoder(16#f7#)) OR
 					(reg_q2208 AND symb_decoder(16#bb#)) OR
 					(reg_q2208 AND symb_decoder(16#cf#)) OR
 					(reg_q2208 AND symb_decoder(16#aa#)) OR
 					(reg_q2208 AND symb_decoder(16#3b#)) OR
 					(reg_q2208 AND symb_decoder(16#da#)) OR
 					(reg_q2208 AND symb_decoder(16#cb#)) OR
 					(reg_q2208 AND symb_decoder(16#b6#)) OR
 					(reg_q2208 AND symb_decoder(16#07#)) OR
 					(reg_q2208 AND symb_decoder(16#5f#)) OR
 					(reg_q2208 AND symb_decoder(16#63#)) OR
 					(reg_q2208 AND symb_decoder(16#3d#)) OR
 					(reg_q2208 AND symb_decoder(16#9c#)) OR
 					(reg_q2208 AND symb_decoder(16#c6#)) OR
 					(reg_q2208 AND symb_decoder(16#a8#)) OR
 					(reg_q2208 AND symb_decoder(16#bf#)) OR
 					(reg_q2208 AND symb_decoder(16#08#)) OR
 					(reg_q2208 AND symb_decoder(16#df#)) OR
 					(reg_q2208 AND symb_decoder(16#af#)) OR
 					(reg_q2208 AND symb_decoder(16#88#)) OR
 					(reg_q2208 AND symb_decoder(16#be#)) OR
 					(reg_q2208 AND symb_decoder(16#1e#)) OR
 					(reg_q2208 AND symb_decoder(16#c7#)) OR
 					(reg_q2208 AND symb_decoder(16#57#)) OR
 					(reg_q2208 AND symb_decoder(16#e6#)) OR
 					(reg_q2208 AND symb_decoder(16#70#)) OR
 					(reg_q2208 AND symb_decoder(16#fc#)) OR
 					(reg_q2208 AND symb_decoder(16#5c#)) OR
 					(reg_q2208 AND symb_decoder(16#81#)) OR
 					(reg_q2208 AND symb_decoder(16#8c#)) OR
 					(reg_q2208 AND symb_decoder(16#39#)) OR
 					(reg_q2208 AND symb_decoder(16#48#)) OR
 					(reg_q2208 AND symb_decoder(16#03#)) OR
 					(reg_q2208 AND symb_decoder(16#84#)) OR
 					(reg_q2208 AND symb_decoder(16#4e#)) OR
 					(reg_q2208 AND symb_decoder(16#9f#)) OR
 					(reg_q2208 AND symb_decoder(16#1a#)) OR
 					(reg_q2208 AND symb_decoder(16#d5#)) OR
 					(reg_q2208 AND symb_decoder(16#35#)) OR
 					(reg_q2208 AND symb_decoder(16#c1#)) OR
 					(reg_q2208 AND symb_decoder(16#19#)) OR
 					(reg_q2208 AND symb_decoder(16#e0#)) OR
 					(reg_q2208 AND symb_decoder(16#de#)) OR
 					(reg_q2208 AND symb_decoder(16#b8#)) OR
 					(reg_q2208 AND symb_decoder(16#a0#)) OR
 					(reg_q2208 AND symb_decoder(16#dd#)) OR
 					(reg_q2208 AND symb_decoder(16#20#)) OR
 					(reg_q2208 AND symb_decoder(16#47#)) OR
 					(reg_q2208 AND symb_decoder(16#c3#)) OR
 					(reg_q2208 AND symb_decoder(16#90#)) OR
 					(reg_q2208 AND symb_decoder(16#9e#)) OR
 					(reg_q2208 AND symb_decoder(16#38#));
reg_q2208_init <= '0' ;
	p_reg_q2208: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2208 <= reg_q2208_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2208 <= reg_q2208_init;
        else
          reg_q2208 <= reg_q2208_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph49

reg_q1209_in <= (reg_q1209 AND symb_decoder(16#20#)) OR
 					(reg_q1209 AND symb_decoder(16#0a#)) OR
 					(reg_q1209 AND symb_decoder(16#0c#)) OR
 					(reg_q1209 AND symb_decoder(16#09#)) OR
 					(reg_q1209 AND symb_decoder(16#0d#)) OR
 					(reg_q1207 AND symb_decoder(16#0c#)) OR
 					(reg_q1207 AND symb_decoder(16#0d#)) OR
 					(reg_q1207 AND symb_decoder(16#09#)) OR
 					(reg_q1207 AND symb_decoder(16#20#)) OR
 					(reg_q1207 AND symb_decoder(16#0a#));
reg_q832_in <= (reg_q828 AND symb_decoder(16#36#)) OR
 					(reg_q828 AND symb_decoder(16#34#)) OR
 					(reg_q828 AND symb_decoder(16#37#)) OR
 					(reg_q828 AND symb_decoder(16#35#)) OR
 					(reg_q828 AND symb_decoder(16#38#)) OR
 					(reg_q828 AND symb_decoder(16#39#)) OR
 					(reg_q828 AND symb_decoder(16#33#)) OR
 					(reg_q828 AND symb_decoder(16#32#)) OR
 					(reg_q828 AND symb_decoder(16#31#)) OR
 					(reg_q828 AND symb_decoder(16#30#)) OR
 					(reg_q848 AND symb_decoder(16#32#)) OR
 					(reg_q848 AND symb_decoder(16#33#)) OR
 					(reg_q848 AND symb_decoder(16#35#)) OR
 					(reg_q848 AND symb_decoder(16#38#)) OR
 					(reg_q848 AND symb_decoder(16#30#)) OR
 					(reg_q848 AND symb_decoder(16#37#)) OR
 					(reg_q848 AND symb_decoder(16#34#)) OR
 					(reg_q848 AND symb_decoder(16#39#)) OR
 					(reg_q848 AND symb_decoder(16#36#)) OR
 					(reg_q848 AND symb_decoder(16#31#)) OR
 					(reg_q832 AND symb_decoder(16#38#)) OR
 					(reg_q832 AND symb_decoder(16#33#)) OR
 					(reg_q832 AND symb_decoder(16#30#)) OR
 					(reg_q832 AND symb_decoder(16#36#)) OR
 					(reg_q832 AND symb_decoder(16#31#)) OR
 					(reg_q832 AND symb_decoder(16#39#)) OR
 					(reg_q832 AND symb_decoder(16#37#)) OR
 					(reg_q832 AND symb_decoder(16#32#)) OR
 					(reg_q832 AND symb_decoder(16#34#)) OR
 					(reg_q832 AND symb_decoder(16#35#));
reg_q1868_in <= (reg_q1866 AND symb_decoder(16#0d#)) OR
 					(reg_q1866 AND symb_decoder(16#20#)) OR
 					(reg_q1866 AND symb_decoder(16#09#)) OR
 					(reg_q1866 AND symb_decoder(16#0c#)) OR
 					(reg_q1866 AND symb_decoder(16#0a#)) OR
 					(reg_q1868 AND symb_decoder(16#0c#)) OR
 					(reg_q1868 AND symb_decoder(16#0d#)) OR
 					(reg_q1868 AND symb_decoder(16#0a#)) OR
 					(reg_q1868 AND symb_decoder(16#09#)) OR
 					(reg_q1868 AND symb_decoder(16#20#));
reg_q842_in <= (reg_q840 AND symb_decoder(16#2e#));
reg_q1918_in <= (reg_q1918 AND symb_decoder(16#0c#)) OR
 					(reg_q1918 AND symb_decoder(16#09#)) OR
 					(reg_q1918 AND symb_decoder(16#0a#)) OR
 					(reg_q1918 AND symb_decoder(16#0d#)) OR
 					(reg_q1918 AND symb_decoder(16#20#)) OR
 					(reg_q1916 AND symb_decoder(16#09#)) OR
 					(reg_q1916 AND symb_decoder(16#0d#)) OR
 					(reg_q1916 AND symb_decoder(16#0a#)) OR
 					(reg_q1916 AND symb_decoder(16#20#)) OR
 					(reg_q1916 AND symb_decoder(16#0c#));
reg_q2066_in <= (reg_q2064 AND symb_decoder(16#0a#)) OR
 					(reg_q2064 AND symb_decoder(16#0d#)) OR
 					(reg_q2064 AND symb_decoder(16#0c#)) OR
 					(reg_q2064 AND symb_decoder(16#20#)) OR
 					(reg_q2064 AND symb_decoder(16#09#)) OR
 					(reg_q2066 AND symb_decoder(16#0c#)) OR
 					(reg_q2066 AND symb_decoder(16#20#)) OR
 					(reg_q2066 AND symb_decoder(16#09#)) OR
 					(reg_q2066 AND symb_decoder(16#0a#)) OR
 					(reg_q2066 AND symb_decoder(16#0d#));
reg_q10_in <= (reg_q8 AND symb_decoder(16#69#)) OR
 					(reg_q8 AND symb_decoder(16#49#));
reg_q2411_in <= (reg_q2409 AND symb_decoder(16#09#)) OR
 					(reg_q2409 AND symb_decoder(16#0d#)) OR
 					(reg_q2409 AND symb_decoder(16#20#)) OR
 					(reg_q2409 AND symb_decoder(16#0c#)) OR
 					(reg_q2409 AND symb_decoder(16#0a#)) OR
 					(reg_q2411 AND symb_decoder(16#09#)) OR
 					(reg_q2411 AND symb_decoder(16#0a#)) OR
 					(reg_q2411 AND symb_decoder(16#20#)) OR
 					(reg_q2411 AND symb_decoder(16#0c#)) OR
 					(reg_q2411 AND symb_decoder(16#0d#));
reg_q880_in <= (reg_q884 AND symb_decoder(16#00#)) OR
 					(reg_q887 AND symb_decoder(16#00#)) OR
 					(reg_q878 AND symb_decoder(16#00#)) OR
 					(reg_q886 AND symb_decoder(16#00#));
reg_q2417_in <= (reg_q2417 AND symb_decoder(16#0d#)) OR
 					(reg_q2417 AND symb_decoder(16#20#)) OR
 					(reg_q2417 AND symb_decoder(16#0a#)) OR
 					(reg_q2417 AND symb_decoder(16#0c#)) OR
 					(reg_q2417 AND symb_decoder(16#09#)) OR
 					(reg_q2415 AND symb_decoder(16#0d#)) OR
 					(reg_q2415 AND symb_decoder(16#09#)) OR
 					(reg_q2415 AND symb_decoder(16#20#)) OR
 					(reg_q2415 AND symb_decoder(16#0a#)) OR
 					(reg_q2415 AND symb_decoder(16#0c#));
reg_q2427_in <= (reg_q2427 AND symb_decoder(16#20#)) OR
 					(reg_q2427 AND symb_decoder(16#09#)) OR
 					(reg_q2427 AND symb_decoder(16#0a#)) OR
 					(reg_q2427 AND symb_decoder(16#0c#)) OR
 					(reg_q2427 AND symb_decoder(16#0d#)) OR
 					(reg_q2425 AND symb_decoder(16#0a#)) OR
 					(reg_q2425 AND symb_decoder(16#0d#)) OR
 					(reg_q2425 AND symb_decoder(16#0c#)) OR
 					(reg_q2425 AND symb_decoder(16#09#)) OR
 					(reg_q2425 AND symb_decoder(16#20#));
reg_q1373_in <= (reg_q1373 AND symb_decoder(16#0d#)) OR
 					(reg_q1373 AND symb_decoder(16#0a#)) OR
 					(reg_q1373 AND symb_decoder(16#20#)) OR
 					(reg_q1373 AND symb_decoder(16#0c#)) OR
 					(reg_q1373 AND symb_decoder(16#09#)) OR
 					(reg_q1371 AND symb_decoder(16#0d#)) OR
 					(reg_q1371 AND symb_decoder(16#0c#)) OR
 					(reg_q1371 AND symb_decoder(16#20#)) OR
 					(reg_q1371 AND symb_decoder(16#09#)) OR
 					(reg_q1371 AND symb_decoder(16#0a#));
reg_q2074_in <= (reg_q2072 AND symb_decoder(16#0c#)) OR
 					(reg_q2072 AND symb_decoder(16#09#)) OR
 					(reg_q2072 AND symb_decoder(16#0d#)) OR
 					(reg_q2072 AND symb_decoder(16#20#)) OR
 					(reg_q2072 AND symb_decoder(16#0a#)) OR
 					(reg_q2074 AND symb_decoder(16#20#)) OR
 					(reg_q2074 AND symb_decoder(16#0d#)) OR
 					(reg_q2074 AND symb_decoder(16#0c#)) OR
 					(reg_q2074 AND symb_decoder(16#09#)) OR
 					(reg_q2074 AND symb_decoder(16#0a#));
reg_q2194_in <= (reg_q2194 AND symb_decoder(16#20#)) OR
 					(reg_q2194 AND symb_decoder(16#0d#)) OR
 					(reg_q2194 AND symb_decoder(16#0c#)) OR
 					(reg_q2194 AND symb_decoder(16#09#)) OR
 					(reg_q2194 AND symb_decoder(16#0a#)) OR
 					(reg_q2192 AND symb_decoder(16#0d#)) OR
 					(reg_q2192 AND symb_decoder(16#20#)) OR
 					(reg_q2192 AND symb_decoder(16#09#)) OR
 					(reg_q2192 AND symb_decoder(16#0a#)) OR
 					(reg_q2192 AND symb_decoder(16#0c#));
reg_q1802_in <= (reg_q1800 AND symb_decoder(16#0d#)) OR
 					(reg_q1800 AND symb_decoder(16#20#)) OR
 					(reg_q1800 AND symb_decoder(16#0a#)) OR
 					(reg_q1800 AND symb_decoder(16#0c#)) OR
 					(reg_q1800 AND symb_decoder(16#09#)) OR
 					(reg_q1802 AND symb_decoder(16#20#)) OR
 					(reg_q1802 AND symb_decoder(16#0c#)) OR
 					(reg_q1802 AND symb_decoder(16#09#)) OR
 					(reg_q1802 AND symb_decoder(16#0d#)) OR
 					(reg_q1802 AND symb_decoder(16#0a#));
reg_q1395_in <= (reg_q1393 AND symb_decoder(16#0a#)) OR
 					(reg_q1393 AND symb_decoder(16#0d#)) OR
 					(reg_q1393 AND symb_decoder(16#09#)) OR
 					(reg_q1393 AND symb_decoder(16#20#)) OR
 					(reg_q1393 AND symb_decoder(16#0c#)) OR
 					(reg_q1395 AND symb_decoder(16#0d#)) OR
 					(reg_q1395 AND symb_decoder(16#09#)) OR
 					(reg_q1395 AND symb_decoder(16#0c#)) OR
 					(reg_q1395 AND symb_decoder(16#20#)) OR
 					(reg_q1395 AND symb_decoder(16#0a#));
reg_q1926_in <= (reg_q1924 AND symb_decoder(16#09#)) OR
 					(reg_q1924 AND symb_decoder(16#0a#)) OR
 					(reg_q1924 AND symb_decoder(16#0d#)) OR
 					(reg_q1924 AND symb_decoder(16#20#)) OR
 					(reg_q1924 AND symb_decoder(16#0c#)) OR
 					(reg_q1926 AND symb_decoder(16#20#)) OR
 					(reg_q1926 AND symb_decoder(16#0d#)) OR
 					(reg_q1926 AND symb_decoder(16#09#)) OR
 					(reg_q1926 AND symb_decoder(16#0c#)) OR
 					(reg_q1926 AND symb_decoder(16#0a#));
reg_q632_in <= (reg_q630 AND symb_decoder(16#09#)) OR
 					(reg_q630 AND symb_decoder(16#0a#)) OR
 					(reg_q630 AND symb_decoder(16#20#)) OR
 					(reg_q630 AND symb_decoder(16#0d#)) OR
 					(reg_q630 AND symb_decoder(16#0c#)) OR
 					(reg_q632 AND symb_decoder(16#0c#)) OR
 					(reg_q632 AND symb_decoder(16#20#)) OR
 					(reg_q632 AND symb_decoder(16#0d#)) OR
 					(reg_q632 AND symb_decoder(16#0a#)) OR
 					(reg_q632 AND symb_decoder(16#09#));
reg_q887_in <= (reg_q884 AND symb_decoder(16#0d#)) OR
 					(reg_q884 AND symb_decoder(16#09#)) OR
 					(reg_q884 AND symb_decoder(16#0a#)) OR
 					(reg_q884 AND symb_decoder(16#0c#)) OR
 					(reg_q884 AND symb_decoder(16#20#)) OR
 					(reg_q887 AND symb_decoder(16#20#)) OR
 					(reg_q887 AND symb_decoder(16#0c#)) OR
 					(reg_q887 AND symb_decoder(16#09#)) OR
 					(reg_q887 AND symb_decoder(16#0d#)) OR
 					(reg_q887 AND symb_decoder(16#0a#));
reg_q1848_in <= (reg_q1848 AND symb_decoder(16#0a#)) OR
 					(reg_q1848 AND symb_decoder(16#20#)) OR
 					(reg_q1848 AND symb_decoder(16#0d#)) OR
 					(reg_q1848 AND symb_decoder(16#0c#)) OR
 					(reg_q1848 AND symb_decoder(16#09#)) OR
 					(reg_q1846 AND symb_decoder(16#0d#)) OR
 					(reg_q1846 AND symb_decoder(16#0a#)) OR
 					(reg_q1846 AND symb_decoder(16#0c#)) OR
 					(reg_q1846 AND symb_decoder(16#20#)) OR
 					(reg_q1846 AND symb_decoder(16#09#));
reg_q2176_in <= (reg_q2172 AND symb_decoder(16#46#)) OR
 					(reg_q2172 AND symb_decoder(16#66#)) OR
 					(reg_q2208 AND symb_decoder(16#66#)) OR
 					(reg_q2208 AND symb_decoder(16#46#));
reg_q16_in <= (reg_q16 AND symb_decoder(16#0a#)) OR
 					(reg_q16 AND symb_decoder(16#0d#)) OR
 					(reg_q16 AND symb_decoder(16#0c#)) OR
 					(reg_q16 AND symb_decoder(16#09#)) OR
 					(reg_q16 AND symb_decoder(16#20#)) OR
 					(reg_q14 AND symb_decoder(16#20#)) OR
 					(reg_q14 AND symb_decoder(16#0d#)) OR
 					(reg_q14 AND symb_decoder(16#0c#)) OR
 					(reg_q14 AND symb_decoder(16#0a#)) OR
 					(reg_q14 AND symb_decoder(16#09#));
reg_q1361_in <= (reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q1359 AND symb_decoder(16#48#)) OR
 					(reg_q1359 AND symb_decoder(16#68#));
reg_q1938_in <= (reg_q1938 AND symb_decoder(16#0a#)) OR
 					(reg_q1938 AND symb_decoder(16#0d#)) OR
 					(reg_q1938 AND symb_decoder(16#20#)) OR
 					(reg_q1938 AND symb_decoder(16#09#)) OR
 					(reg_q1938 AND symb_decoder(16#0c#)) OR
 					(reg_q1936 AND symb_decoder(16#0c#)) OR
 					(reg_q1936 AND symb_decoder(16#0d#)) OR
 					(reg_q1936 AND symb_decoder(16#20#)) OR
 					(reg_q1936 AND symb_decoder(16#09#)) OR
 					(reg_q1936 AND symb_decoder(16#0a#));
reg_q1383_in <= (reg_q1381 AND symb_decoder(16#09#)) OR
 					(reg_q1381 AND symb_decoder(16#20#)) OR
 					(reg_q1381 AND symb_decoder(16#0a#)) OR
 					(reg_q1381 AND symb_decoder(16#0c#)) OR
 					(reg_q1381 AND symb_decoder(16#0d#)) OR
 					(reg_q1383 AND symb_decoder(16#0c#)) OR
 					(reg_q1383 AND symb_decoder(16#09#)) OR
 					(reg_q1383 AND symb_decoder(16#0d#)) OR
 					(reg_q1383 AND symb_decoder(16#0a#)) OR
 					(reg_q1383 AND symb_decoder(16#20#));
reg_q1880_in <= (reg_q1878 AND symb_decoder(16#20#)) OR
 					(reg_q1878 AND symb_decoder(16#0d#)) OR
 					(reg_q1878 AND symb_decoder(16#0a#)) OR
 					(reg_q1878 AND symb_decoder(16#09#)) OR
 					(reg_q1878 AND symb_decoder(16#0c#)) OR
 					(reg_q1880 AND symb_decoder(16#0a#)) OR
 					(reg_q1880 AND symb_decoder(16#0c#)) OR
 					(reg_q1880 AND symb_decoder(16#09#)) OR
 					(reg_q1880 AND symb_decoder(16#20#)) OR
 					(reg_q1880 AND symb_decoder(16#0d#));
reg_q1886_in <= (reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q1884 AND symb_decoder(16#53#)) OR
 					(reg_q1884 AND symb_decoder(16#73#));
reg_q864_in <= (reg_q864 AND symb_decoder(16#0a#)) OR
 					(reg_q864 AND symb_decoder(16#20#)) OR
 					(reg_q864 AND symb_decoder(16#09#)) OR
 					(reg_q864 AND symb_decoder(16#0d#)) OR
 					(reg_q864 AND symb_decoder(16#0c#)) OR
 					(reg_q862 AND symb_decoder(16#0d#)) OR
 					(reg_q862 AND symb_decoder(16#0a#)) OR
 					(reg_q862 AND symb_decoder(16#09#)) OR
 					(reg_q862 AND symb_decoder(16#0c#)) OR
 					(reg_q862 AND symb_decoder(16#20#));
reg_q1816_in <= (reg_q1814 AND symb_decoder(16#0a#)) OR
 					(reg_q1814 AND symb_decoder(16#0d#)) OR
 					(reg_q1814 AND symb_decoder(16#20#)) OR
 					(reg_q1814 AND symb_decoder(16#09#)) OR
 					(reg_q1814 AND symb_decoder(16#0c#)) OR
 					(reg_q1816 AND symb_decoder(16#0c#)) OR
 					(reg_q1816 AND symb_decoder(16#0a#)) OR
 					(reg_q1816 AND symb_decoder(16#09#)) OR
 					(reg_q1816 AND symb_decoder(16#0d#)) OR
 					(reg_q1816 AND symb_decoder(16#20#));
reg_q893_in <= (reg_q889 AND symb_decoder(16#5c#)) OR
 					(reg_q896 AND symb_decoder(16#5c#));
reg_q604_in <= (reg_q604 AND symb_decoder(16#0c#)) OR
 					(reg_q604 AND symb_decoder(16#09#)) OR
 					(reg_q604 AND symb_decoder(16#0a#)) OR
 					(reg_q604 AND symb_decoder(16#20#)) OR
 					(reg_q604 AND symb_decoder(16#0d#)) OR
 					(reg_q602 AND symb_decoder(16#09#)) OR
 					(reg_q602 AND symb_decoder(16#0a#)) OR
 					(reg_q602 AND symb_decoder(16#20#)) OR
 					(reg_q602 AND symb_decoder(16#0d#)) OR
 					(reg_q602 AND symb_decoder(16#0c#));
reg_q1221_in <= (reg_q1219 AND symb_decoder(16#0d#)) OR
 					(reg_q1219 AND symb_decoder(16#20#)) OR
 					(reg_q1219 AND symb_decoder(16#09#)) OR
 					(reg_q1219 AND symb_decoder(16#0a#)) OR
 					(reg_q1219 AND symb_decoder(16#0c#)) OR
 					(reg_q1221 AND symb_decoder(16#0a#)) OR
 					(reg_q1221 AND symb_decoder(16#20#)) OR
 					(reg_q1221 AND symb_decoder(16#0d#)) OR
 					(reg_q1221 AND symb_decoder(16#09#)) OR
 					(reg_q1221 AND symb_decoder(16#0c#));
reg_q2385_in <= (reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2383 AND symb_decoder(16#23#));
reg_q596_in <= (reg_q594 AND symb_decoder(16#0a#)) OR
 					(reg_q594 AND symb_decoder(16#09#)) OR
 					(reg_q594 AND symb_decoder(16#0c#)) OR
 					(reg_q594 AND symb_decoder(16#0d#)) OR
 					(reg_q594 AND symb_decoder(16#20#)) OR
 					(reg_q596 AND symb_decoder(16#0d#)) OR
 					(reg_q596 AND symb_decoder(16#0c#)) OR
 					(reg_q596 AND symb_decoder(16#20#)) OR
 					(reg_q596 AND symb_decoder(16#0a#)) OR
 					(reg_q596 AND symb_decoder(16#09#));
reg_q716_in <= (reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q715 AND symb_decoder(16#64#)) OR
 					(reg_q715 AND symb_decoder(16#44#));
reg_q1904_in <= (reg_q1904 AND symb_decoder(16#20#)) OR
 					(reg_q1904 AND symb_decoder(16#0c#)) OR
 					(reg_q1904 AND symb_decoder(16#0d#)) OR
 					(reg_q1904 AND symb_decoder(16#09#)) OR
 					(reg_q1904 AND symb_decoder(16#0a#)) OR
 					(reg_q1902 AND symb_decoder(16#20#)) OR
 					(reg_q1902 AND symb_decoder(16#0c#)) OR
 					(reg_q1902 AND symb_decoder(16#09#)) OR
 					(reg_q1902 AND symb_decoder(16#0a#)) OR
 					(reg_q1902 AND symb_decoder(16#0d#));
reg_q458_in <= (reg_q456 AND symb_decoder(16#64#)) OR
 					(reg_q456 AND symb_decoder(16#44#));
reg_q460_in <= (reg_q458 AND symb_decoder(16#79#)) OR
 					(reg_q458 AND symb_decoder(16#59#));
reg_q22_in <= (reg_q20 AND symb_decoder(16#0d#)) OR
 					(reg_q20 AND symb_decoder(16#0a#)) OR
 					(reg_q20 AND symb_decoder(16#20#)) OR
 					(reg_q20 AND symb_decoder(16#0c#)) OR
 					(reg_q20 AND symb_decoder(16#09#)) OR
 					(reg_q22 AND symb_decoder(16#0d#)) OR
 					(reg_q22 AND symb_decoder(16#09#)) OR
 					(reg_q22 AND symb_decoder(16#20#)) OR
 					(reg_q22 AND symb_decoder(16#0c#)) OR
 					(reg_q22 AND symb_decoder(16#0a#));
reg_q558_in <= (reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q556 AND symb_decoder(16#62#)) OR
 					(reg_q556 AND symb_decoder(16#42#));
reg_q811_in <= (reg_q809 AND symb_decoder(16#5e#));
reg_q566_in <= (reg_q564 AND symb_decoder(16#3d#));
reg_q1201_in <= (reg_q1199 AND symb_decoder(16#50#)) OR
 					(reg_q1199 AND symb_decoder(16#70#));
reg_q886_in <= (reg_q893 AND symb_decoder(16#5d#));
reg_q2054_in <= (reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2052 AND symb_decoder(16#54#));
reg_q93_in <= (reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q92 AND symb_decoder(16#30#));
reg_q456_in <= (reg_q454 AND symb_decoder(16#4f#)) OR
 					(reg_q454 AND symb_decoder(16#6f#));
reg_q852_in <= (reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q850 AND symb_decoder(16#5b#));
reg_q95_in <= (reg_q93 AND symb_decoder(16#30#));
reg_fullgraph49_init <= "000000";

reg_fullgraph49_sel <= "000000000000000" & reg_q95_in & reg_q852_in & reg_q456_in & reg_q93_in & reg_q2054_in & reg_q886_in & reg_q1201_in & reg_q566_in & reg_q811_in & reg_q558_in & reg_q22_in & reg_q460_in & reg_q458_in & reg_q1904_in & reg_q716_in & reg_q596_in & reg_q2385_in & reg_q1221_in & reg_q604_in & reg_q893_in & reg_q1816_in & reg_q864_in & reg_q1886_in & reg_q1880_in & reg_q1383_in & reg_q1938_in & reg_q1361_in & reg_q16_in & reg_q2176_in & reg_q1848_in & reg_q887_in & reg_q632_in & reg_q1926_in & reg_q1395_in & reg_q1802_in & reg_q2194_in & reg_q2074_in & reg_q1373_in & reg_q2427_in & reg_q2417_in & reg_q880_in & reg_q2411_in & reg_q10_in & reg_q2066_in & reg_q1918_in & reg_q842_in & reg_q1868_in & reg_q832_in & reg_q1209_in;

	--coder fullgraph49
with reg_fullgraph49_sel select
reg_fullgraph49_in <=
	"000001" when "0000000000000000000000000000000000000000000000000000000000000001",
	"000010" when "0000000000000000000000000000000000000000000000000000000000000010",
	"000011" when "0000000000000000000000000000000000000000000000000000000000000100",
	"000100" when "0000000000000000000000000000000000000000000000000000000000001000",
	"000101" when "0000000000000000000000000000000000000000000000000000000000010000",
	"000110" when "0000000000000000000000000000000000000000000000000000000000100000",
	"000111" when "0000000000000000000000000000000000000000000000000000000001000000",
	"001000" when "0000000000000000000000000000000000000000000000000000000010000000",
	"001001" when "0000000000000000000000000000000000000000000000000000000100000000",
	"001010" when "0000000000000000000000000000000000000000000000000000001000000000",
	"001011" when "0000000000000000000000000000000000000000000000000000010000000000",
	"001100" when "0000000000000000000000000000000000000000000000000000100000000000",
	"001101" when "0000000000000000000000000000000000000000000000000001000000000000",
	"001110" when "0000000000000000000000000000000000000000000000000010000000000000",
	"001111" when "0000000000000000000000000000000000000000000000000100000000000000",
	"010000" when "0000000000000000000000000000000000000000000000001000000000000000",
	"010001" when "0000000000000000000000000000000000000000000000010000000000000000",
	"010010" when "0000000000000000000000000000000000000000000000100000000000000000",
	"010011" when "0000000000000000000000000000000000000000000001000000000000000000",
	"010100" when "0000000000000000000000000000000000000000000010000000000000000000",
	"010101" when "0000000000000000000000000000000000000000000100000000000000000000",
	"010110" when "0000000000000000000000000000000000000000001000000000000000000000",
	"010111" when "0000000000000000000000000000000000000000010000000000000000000000",
	"011000" when "0000000000000000000000000000000000000000100000000000000000000000",
	"011001" when "0000000000000000000000000000000000000001000000000000000000000000",
	"011010" when "0000000000000000000000000000000000000010000000000000000000000000",
	"011011" when "0000000000000000000000000000000000000100000000000000000000000000",
	"011100" when "0000000000000000000000000000000000001000000000000000000000000000",
	"011101" when "0000000000000000000000000000000000010000000000000000000000000000",
	"011110" when "0000000000000000000000000000000000100000000000000000000000000000",
	"011111" when "0000000000000000000000000000000001000000000000000000000000000000",
	"100000" when "0000000000000000000000000000000010000000000000000000000000000000",
	"100001" when "0000000000000000000000000000000100000000000000000000000000000000",
	"100010" when "0000000000000000000000000000001000000000000000000000000000000000",
	"100011" when "0000000000000000000000000000010000000000000000000000000000000000",
	"100100" when "0000000000000000000000000000100000000000000000000000000000000000",
	"100101" when "0000000000000000000000000001000000000000000000000000000000000000",
	"100110" when "0000000000000000000000000010000000000000000000000000000000000000",
	"100111" when "0000000000000000000000000100000000000000000000000000000000000000",
	"101000" when "0000000000000000000000001000000000000000000000000000000000000000",
	"101001" when "0000000000000000000000010000000000000000000000000000000000000000",
	"101010" when "0000000000000000000000100000000000000000000000000000000000000000",
	"101011" when "0000000000000000000001000000000000000000000000000000000000000000",
	"101100" when "0000000000000000000010000000000000000000000000000000000000000000",
	"101101" when "0000000000000000000100000000000000000000000000000000000000000000",
	"101110" when "0000000000000000001000000000000000000000000000000000000000000000",
	"101111" when "0000000000000000010000000000000000000000000000000000000000000000",
	"110000" when "0000000000000000100000000000000000000000000000000000000000000000",
	"110001" when "0000000000000001000000000000000000000000000000000000000000000000",
	"000000" when others;
 --end coder

	p_reg_fullgraph49: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph49 <= reg_fullgraph49_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph49 <= reg_fullgraph49_init;
        else
          reg_fullgraph49 <= reg_fullgraph49_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph49

		reg_q1209 <= '1' when reg_fullgraph49 = "000001" else '0'; 
		reg_q832 <= '1' when reg_fullgraph49 = "000010" else '0'; 
		reg_q1868 <= '1' when reg_fullgraph49 = "000011" else '0'; 
		reg_q842 <= '1' when reg_fullgraph49 = "000100" else '0'; 
		reg_q1918 <= '1' when reg_fullgraph49 = "000101" else '0'; 
		reg_q2066 <= '1' when reg_fullgraph49 = "000110" else '0'; 
		reg_q10 <= '1' when reg_fullgraph49 = "000111" else '0'; 
		reg_q2411 <= '1' when reg_fullgraph49 = "001000" else '0'; 
		reg_q880 <= '1' when reg_fullgraph49 = "001001" else '0'; 
		reg_q2417 <= '1' when reg_fullgraph49 = "001010" else '0'; 
		reg_q2427 <= '1' when reg_fullgraph49 = "001011" else '0'; 
		reg_q1373 <= '1' when reg_fullgraph49 = "001100" else '0'; 
		reg_q2074 <= '1' when reg_fullgraph49 = "001101" else '0'; 
		reg_q2194 <= '1' when reg_fullgraph49 = "001110" else '0'; 
		reg_q1802 <= '1' when reg_fullgraph49 = "001111" else '0'; 
		reg_q1395 <= '1' when reg_fullgraph49 = "010000" else '0'; 
		reg_q1926 <= '1' when reg_fullgraph49 = "010001" else '0'; 
		reg_q632 <= '1' when reg_fullgraph49 = "010010" else '0'; 
		reg_q887 <= '1' when reg_fullgraph49 = "010011" else '0'; 
		reg_q1848 <= '1' when reg_fullgraph49 = "010100" else '0'; 
		reg_q2176 <= '1' when reg_fullgraph49 = "010101" else '0'; 
		reg_q16 <= '1' when reg_fullgraph49 = "010110" else '0'; 
		reg_q1361 <= '1' when reg_fullgraph49 = "010111" else '0'; 
		reg_q1938 <= '1' when reg_fullgraph49 = "011000" else '0'; 
		reg_q1383 <= '1' when reg_fullgraph49 = "011001" else '0'; 
		reg_q1880 <= '1' when reg_fullgraph49 = "011010" else '0'; 
		reg_q1886 <= '1' when reg_fullgraph49 = "011011" else '0'; 
		reg_q864 <= '1' when reg_fullgraph49 = "011100" else '0'; 
		reg_q1816 <= '1' when reg_fullgraph49 = "011101" else '0'; 
		reg_q893 <= '1' when reg_fullgraph49 = "011110" else '0'; 
		reg_q604 <= '1' when reg_fullgraph49 = "011111" else '0'; 
		reg_q1221 <= '1' when reg_fullgraph49 = "100000" else '0'; 
		reg_q2385 <= '1' when reg_fullgraph49 = "100001" else '0'; 
		reg_q596 <= '1' when reg_fullgraph49 = "100010" else '0'; 
		reg_q716 <= '1' when reg_fullgraph49 = "100011" else '0'; 
		reg_q1904 <= '1' when reg_fullgraph49 = "100100" else '0'; 
		reg_q458 <= '1' when reg_fullgraph49 = "100101" else '0'; 
		reg_q460 <= '1' when reg_fullgraph49 = "100110" else '0'; 
		reg_q22 <= '1' when reg_fullgraph49 = "100111" else '0'; 
		reg_q558 <= '1' when reg_fullgraph49 = "101000" else '0'; 
		reg_q811 <= '1' when reg_fullgraph49 = "101001" else '0'; 
		reg_q566 <= '1' when reg_fullgraph49 = "101010" else '0'; 
		reg_q1201 <= '1' when reg_fullgraph49 = "101011" else '0'; 
		reg_q886 <= '1' when reg_fullgraph49 = "101100" else '0'; 
		reg_q2054 <= '1' when reg_fullgraph49 = "101101" else '0'; 
		reg_q93 <= '1' when reg_fullgraph49 = "101110" else '0'; 
		reg_q456 <= '1' when reg_fullgraph49 = "101111" else '0'; 
		reg_q852 <= '1' when reg_fullgraph49 = "110000" else '0'; 
		reg_q95 <= '1' when reg_fullgraph49 = "110001" else '0'; 
--end decoder 

reg_q2518_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2518 AND symb_decoder(16#60#)) OR
 					(reg_q2518 AND symb_decoder(16#6e#)) OR
 					(reg_q2518 AND symb_decoder(16#a6#)) OR
 					(reg_q2518 AND symb_decoder(16#c7#)) OR
 					(reg_q2518 AND symb_decoder(16#24#)) OR
 					(reg_q2518 AND symb_decoder(16#b4#)) OR
 					(reg_q2518 AND symb_decoder(16#6a#)) OR
 					(reg_q2518 AND symb_decoder(16#77#)) OR
 					(reg_q2518 AND symb_decoder(16#db#)) OR
 					(reg_q2518 AND symb_decoder(16#d5#)) OR
 					(reg_q2518 AND symb_decoder(16#f8#)) OR
 					(reg_q2518 AND symb_decoder(16#d3#)) OR
 					(reg_q2518 AND symb_decoder(16#fa#)) OR
 					(reg_q2518 AND symb_decoder(16#0c#)) OR
 					(reg_q2518 AND symb_decoder(16#19#)) OR
 					(reg_q2518 AND symb_decoder(16#31#)) OR
 					(reg_q2518 AND symb_decoder(16#a7#)) OR
 					(reg_q2518 AND symb_decoder(16#21#)) OR
 					(reg_q2518 AND symb_decoder(16#9d#)) OR
 					(reg_q2518 AND symb_decoder(16#dc#)) OR
 					(reg_q2518 AND symb_decoder(16#ca#)) OR
 					(reg_q2518 AND symb_decoder(16#3b#)) OR
 					(reg_q2518 AND symb_decoder(16#ea#)) OR
 					(reg_q2518 AND symb_decoder(16#92#)) OR
 					(reg_q2518 AND symb_decoder(16#53#)) OR
 					(reg_q2518 AND symb_decoder(16#98#)) OR
 					(reg_q2518 AND symb_decoder(16#56#)) OR
 					(reg_q2518 AND symb_decoder(16#b6#)) OR
 					(reg_q2518 AND symb_decoder(16#f6#)) OR
 					(reg_q2518 AND symb_decoder(16#3c#)) OR
 					(reg_q2518 AND symb_decoder(16#4f#)) OR
 					(reg_q2518 AND symb_decoder(16#90#)) OR
 					(reg_q2518 AND symb_decoder(16#3f#)) OR
 					(reg_q2518 AND symb_decoder(16#09#)) OR
 					(reg_q2518 AND symb_decoder(16#36#)) OR
 					(reg_q2518 AND symb_decoder(16#ec#)) OR
 					(reg_q2518 AND symb_decoder(16#fc#)) OR
 					(reg_q2518 AND symb_decoder(16#1b#)) OR
 					(reg_q2518 AND symb_decoder(16#0b#)) OR
 					(reg_q2518 AND symb_decoder(16#22#)) OR
 					(reg_q2518 AND symb_decoder(16#c5#)) OR
 					(reg_q2518 AND symb_decoder(16#0a#)) OR
 					(reg_q2518 AND symb_decoder(16#ff#)) OR
 					(reg_q2518 AND symb_decoder(16#84#)) OR
 					(reg_q2518 AND symb_decoder(16#cb#)) OR
 					(reg_q2518 AND symb_decoder(16#06#)) OR
 					(reg_q2518 AND symb_decoder(16#7b#)) OR
 					(reg_q2518 AND symb_decoder(16#bd#)) OR
 					(reg_q2518 AND symb_decoder(16#b3#)) OR
 					(reg_q2518 AND symb_decoder(16#58#)) OR
 					(reg_q2518 AND symb_decoder(16#9a#)) OR
 					(reg_q2518 AND symb_decoder(16#b8#)) OR
 					(reg_q2518 AND symb_decoder(16#ef#)) OR
 					(reg_q2518 AND symb_decoder(16#df#)) OR
 					(reg_q2518 AND symb_decoder(16#bb#)) OR
 					(reg_q2518 AND symb_decoder(16#85#)) OR
 					(reg_q2518 AND symb_decoder(16#57#)) OR
 					(reg_q2518 AND symb_decoder(16#62#)) OR
 					(reg_q2518 AND symb_decoder(16#9c#)) OR
 					(reg_q2518 AND symb_decoder(16#6d#)) OR
 					(reg_q2518 AND symb_decoder(16#8f#)) OR
 					(reg_q2518 AND symb_decoder(16#8b#)) OR
 					(reg_q2518 AND symb_decoder(16#63#)) OR
 					(reg_q2518 AND symb_decoder(16#28#)) OR
 					(reg_q2518 AND symb_decoder(16#1d#)) OR
 					(reg_q2518 AND symb_decoder(16#10#)) OR
 					(reg_q2518 AND symb_decoder(16#3a#)) OR
 					(reg_q2518 AND symb_decoder(16#95#)) OR
 					(reg_q2518 AND symb_decoder(16#33#)) OR
 					(reg_q2518 AND symb_decoder(16#81#)) OR
 					(reg_q2518 AND symb_decoder(16#49#)) OR
 					(reg_q2518 AND symb_decoder(16#8a#)) OR
 					(reg_q2518 AND symb_decoder(16#89#)) OR
 					(reg_q2518 AND symb_decoder(16#e4#)) OR
 					(reg_q2518 AND symb_decoder(16#25#)) OR
 					(reg_q2518 AND symb_decoder(16#13#)) OR
 					(reg_q2518 AND symb_decoder(16#15#)) OR
 					(reg_q2518 AND symb_decoder(16#48#)) OR
 					(reg_q2518 AND symb_decoder(16#45#)) OR
 					(reg_q2518 AND symb_decoder(16#61#)) OR
 					(reg_q2518 AND symb_decoder(16#f1#)) OR
 					(reg_q2518 AND symb_decoder(16#c0#)) OR
 					(reg_q2518 AND symb_decoder(16#e9#)) OR
 					(reg_q2518 AND symb_decoder(16#44#)) OR
 					(reg_q2518 AND symb_decoder(16#76#)) OR
 					(reg_q2518 AND symb_decoder(16#5c#)) OR
 					(reg_q2518 AND symb_decoder(16#42#)) OR
 					(reg_q2518 AND symb_decoder(16#7c#)) OR
 					(reg_q2518 AND symb_decoder(16#d1#)) OR
 					(reg_q2518 AND symb_decoder(16#4a#)) OR
 					(reg_q2518 AND symb_decoder(16#47#)) OR
 					(reg_q2518 AND symb_decoder(16#a2#)) OR
 					(reg_q2518 AND symb_decoder(16#4d#)) OR
 					(reg_q2518 AND symb_decoder(16#1e#)) OR
 					(reg_q2518 AND symb_decoder(16#79#)) OR
 					(reg_q2518 AND symb_decoder(16#1c#)) OR
 					(reg_q2518 AND symb_decoder(16#41#)) OR
 					(reg_q2518 AND symb_decoder(16#ab#)) OR
 					(reg_q2518 AND symb_decoder(16#32#)) OR
 					(reg_q2518 AND symb_decoder(16#b1#)) OR
 					(reg_q2518 AND symb_decoder(16#7a#)) OR
 					(reg_q2518 AND symb_decoder(16#b0#)) OR
 					(reg_q2518 AND symb_decoder(16#26#)) OR
 					(reg_q2518 AND symb_decoder(16#34#)) OR
 					(reg_q2518 AND symb_decoder(16#e1#)) OR
 					(reg_q2518 AND symb_decoder(16#a1#)) OR
 					(reg_q2518 AND symb_decoder(16#8e#)) OR
 					(reg_q2518 AND symb_decoder(16#71#)) OR
 					(reg_q2518 AND symb_decoder(16#af#)) OR
 					(reg_q2518 AND symb_decoder(16#de#)) OR
 					(reg_q2518 AND symb_decoder(16#82#)) OR
 					(reg_q2518 AND symb_decoder(16#d8#)) OR
 					(reg_q2518 AND symb_decoder(16#ba#)) OR
 					(reg_q2518 AND symb_decoder(16#2e#)) OR
 					(reg_q2518 AND symb_decoder(16#35#)) OR
 					(reg_q2518 AND symb_decoder(16#c1#)) OR
 					(reg_q2518 AND symb_decoder(16#97#)) OR
 					(reg_q2518 AND symb_decoder(16#12#)) OR
 					(reg_q2518 AND symb_decoder(16#d4#)) OR
 					(reg_q2518 AND symb_decoder(16#0e#)) OR
 					(reg_q2518 AND symb_decoder(16#05#)) OR
 					(reg_q2518 AND symb_decoder(16#67#)) OR
 					(reg_q2518 AND symb_decoder(16#c4#)) OR
 					(reg_q2518 AND symb_decoder(16#20#)) OR
 					(reg_q2518 AND symb_decoder(16#70#)) OR
 					(reg_q2518 AND symb_decoder(16#2f#)) OR
 					(reg_q2518 AND symb_decoder(16#a9#)) OR
 					(reg_q2518 AND symb_decoder(16#73#)) OR
 					(reg_q2518 AND symb_decoder(16#a4#)) OR
 					(reg_q2518 AND symb_decoder(16#38#)) OR
 					(reg_q2518 AND symb_decoder(16#fd#)) OR
 					(reg_q2518 AND symb_decoder(16#96#)) OR
 					(reg_q2518 AND symb_decoder(16#11#)) OR
 					(reg_q2518 AND symb_decoder(16#9b#)) OR
 					(reg_q2518 AND symb_decoder(16#5e#)) OR
 					(reg_q2518 AND symb_decoder(16#55#)) OR
 					(reg_q2518 AND symb_decoder(16#75#)) OR
 					(reg_q2518 AND symb_decoder(16#ed#)) OR
 					(reg_q2518 AND symb_decoder(16#ad#)) OR
 					(reg_q2518 AND symb_decoder(16#23#)) OR
 					(reg_q2518 AND symb_decoder(16#27#)) OR
 					(reg_q2518 AND symb_decoder(16#29#)) OR
 					(reg_q2518 AND symb_decoder(16#c9#)) OR
 					(reg_q2518 AND symb_decoder(16#0d#)) OR
 					(reg_q2518 AND symb_decoder(16#59#)) OR
 					(reg_q2518 AND symb_decoder(16#d7#)) OR
 					(reg_q2518 AND symb_decoder(16#3d#)) OR
 					(reg_q2518 AND symb_decoder(16#9f#)) OR
 					(reg_q2518 AND symb_decoder(16#5b#)) OR
 					(reg_q2518 AND symb_decoder(16#01#)) OR
 					(reg_q2518 AND symb_decoder(16#d2#)) OR
 					(reg_q2518 AND symb_decoder(16#aa#)) OR
 					(reg_q2518 AND symb_decoder(16#04#)) OR
 					(reg_q2518 AND symb_decoder(16#52#)) OR
 					(reg_q2518 AND symb_decoder(16#c2#)) OR
 					(reg_q2518 AND symb_decoder(16#a8#)) OR
 					(reg_q2518 AND symb_decoder(16#2a#)) OR
 					(reg_q2518 AND symb_decoder(16#16#)) OR
 					(reg_q2518 AND symb_decoder(16#07#)) OR
 					(reg_q2518 AND symb_decoder(16#50#)) OR
 					(reg_q2518 AND symb_decoder(16#a0#)) OR
 					(reg_q2518 AND symb_decoder(16#fb#)) OR
 					(reg_q2518 AND symb_decoder(16#51#)) OR
 					(reg_q2518 AND symb_decoder(16#87#)) OR
 					(reg_q2518 AND symb_decoder(16#9e#)) OR
 					(reg_q2518 AND symb_decoder(16#1f#)) OR
 					(reg_q2518 AND symb_decoder(16#bc#)) OR
 					(reg_q2518 AND symb_decoder(16#b5#)) OR
 					(reg_q2518 AND symb_decoder(16#94#)) OR
 					(reg_q2518 AND symb_decoder(16#69#)) OR
 					(reg_q2518 AND symb_decoder(16#2c#)) OR
 					(reg_q2518 AND symb_decoder(16#40#)) OR
 					(reg_q2518 AND symb_decoder(16#f3#)) OR
 					(reg_q2518 AND symb_decoder(16#fe#)) OR
 					(reg_q2518 AND symb_decoder(16#f2#)) OR
 					(reg_q2518 AND symb_decoder(16#e3#)) OR
 					(reg_q2518 AND symb_decoder(16#2b#)) OR
 					(reg_q2518 AND symb_decoder(16#37#)) OR
 					(reg_q2518 AND symb_decoder(16#83#)) OR
 					(reg_q2518 AND symb_decoder(16#bf#)) OR
 					(reg_q2518 AND symb_decoder(16#e5#)) OR
 					(reg_q2518 AND symb_decoder(16#91#)) OR
 					(reg_q2518 AND symb_decoder(16#6b#)) OR
 					(reg_q2518 AND symb_decoder(16#c8#)) OR
 					(reg_q2518 AND symb_decoder(16#e2#)) OR
 					(reg_q2518 AND symb_decoder(16#ac#)) OR
 					(reg_q2518 AND symb_decoder(16#cf#)) OR
 					(reg_q2518 AND symb_decoder(16#65#)) OR
 					(reg_q2518 AND symb_decoder(16#66#)) OR
 					(reg_q2518 AND symb_decoder(16#f4#)) OR
 					(reg_q2518 AND symb_decoder(16#7d#)) OR
 					(reg_q2518 AND symb_decoder(16#da#)) OR
 					(reg_q2518 AND symb_decoder(16#5f#)) OR
 					(reg_q2518 AND symb_decoder(16#8d#)) OR
 					(reg_q2518 AND symb_decoder(16#7f#)) OR
 					(reg_q2518 AND symb_decoder(16#be#)) OR
 					(reg_q2518 AND symb_decoder(16#d6#)) OR
 					(reg_q2518 AND symb_decoder(16#39#)) OR
 					(reg_q2518 AND symb_decoder(16#0f#)) OR
 					(reg_q2518 AND symb_decoder(16#80#)) OR
 					(reg_q2518 AND symb_decoder(16#d0#)) OR
 					(reg_q2518 AND symb_decoder(16#a3#)) OR
 					(reg_q2518 AND symb_decoder(16#99#)) OR
 					(reg_q2518 AND symb_decoder(16#c6#)) OR
 					(reg_q2518 AND symb_decoder(16#8c#)) OR
 					(reg_q2518 AND symb_decoder(16#5a#)) OR
 					(reg_q2518 AND symb_decoder(16#d9#)) OR
 					(reg_q2518 AND symb_decoder(16#c3#)) OR
 					(reg_q2518 AND symb_decoder(16#b9#)) OR
 					(reg_q2518 AND symb_decoder(16#00#)) OR
 					(reg_q2518 AND symb_decoder(16#43#)) OR
 					(reg_q2518 AND symb_decoder(16#03#)) OR
 					(reg_q2518 AND symb_decoder(16#cc#)) OR
 					(reg_q2518 AND symb_decoder(16#88#)) OR
 					(reg_q2518 AND symb_decoder(16#78#)) OR
 					(reg_q2518 AND symb_decoder(16#eb#)) OR
 					(reg_q2518 AND symb_decoder(16#dd#)) OR
 					(reg_q2518 AND symb_decoder(16#3e#)) OR
 					(reg_q2518 AND symb_decoder(16#f9#)) OR
 					(reg_q2518 AND symb_decoder(16#b7#)) OR
 					(reg_q2518 AND symb_decoder(16#4c#)) OR
 					(reg_q2518 AND symb_decoder(16#ee#)) OR
 					(reg_q2518 AND symb_decoder(16#30#)) OR
 					(reg_q2518 AND symb_decoder(16#cd#)) OR
 					(reg_q2518 AND symb_decoder(16#54#)) OR
 					(reg_q2518 AND symb_decoder(16#68#)) OR
 					(reg_q2518 AND symb_decoder(16#1a#)) OR
 					(reg_q2518 AND symb_decoder(16#4e#)) OR
 					(reg_q2518 AND symb_decoder(16#46#)) OR
 					(reg_q2518 AND symb_decoder(16#74#)) OR
 					(reg_q2518 AND symb_decoder(16#64#)) OR
 					(reg_q2518 AND symb_decoder(16#7e#)) OR
 					(reg_q2518 AND symb_decoder(16#14#)) OR
 					(reg_q2518 AND symb_decoder(16#f7#)) OR
 					(reg_q2518 AND symb_decoder(16#ae#)) OR
 					(reg_q2518 AND symb_decoder(16#17#)) OR
 					(reg_q2518 AND symb_decoder(16#b2#)) OR
 					(reg_q2518 AND symb_decoder(16#86#)) OR
 					(reg_q2518 AND symb_decoder(16#f0#)) OR
 					(reg_q2518 AND symb_decoder(16#72#)) OR
 					(reg_q2518 AND symb_decoder(16#02#)) OR
 					(reg_q2518 AND symb_decoder(16#93#)) OR
 					(reg_q2518 AND symb_decoder(16#e0#)) OR
 					(reg_q2518 AND symb_decoder(16#08#)) OR
 					(reg_q2518 AND symb_decoder(16#f5#)) OR
 					(reg_q2518 AND symb_decoder(16#2d#)) OR
 					(reg_q2518 AND symb_decoder(16#18#)) OR
 					(reg_q2518 AND symb_decoder(16#a5#)) OR
 					(reg_q2518 AND symb_decoder(16#4b#)) OR
 					(reg_q2518 AND symb_decoder(16#6c#)) OR
 					(reg_q2518 AND symb_decoder(16#5d#)) OR
 					(reg_q2518 AND symb_decoder(16#e6#)) OR
 					(reg_q2518 AND symb_decoder(16#e7#)) OR
 					(reg_q2518 AND symb_decoder(16#6f#)) OR
 					(reg_q2518 AND symb_decoder(16#e8#)) OR
 					(reg_q2518 AND symb_decoder(16#ce#));
reg_q2518_init <= '0' ;
	p_reg_q2518: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2518 <= reg_q2518_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2518 <= reg_q2518_init;
        else
          reg_q2518 <= reg_q2518_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2052_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q2052 AND symb_decoder(16#2a#)) OR
 					(reg_q2052 AND symb_decoder(16#67#)) OR
 					(reg_q2052 AND symb_decoder(16#06#)) OR
 					(reg_q2052 AND symb_decoder(16#bf#)) OR
 					(reg_q2052 AND symb_decoder(16#92#)) OR
 					(reg_q2052 AND symb_decoder(16#ff#)) OR
 					(reg_q2052 AND symb_decoder(16#56#)) OR
 					(reg_q2052 AND symb_decoder(16#c8#)) OR
 					(reg_q2052 AND symb_decoder(16#b4#)) OR
 					(reg_q2052 AND symb_decoder(16#d8#)) OR
 					(reg_q2052 AND symb_decoder(16#4d#)) OR
 					(reg_q2052 AND symb_decoder(16#fb#)) OR
 					(reg_q2052 AND symb_decoder(16#a3#)) OR
 					(reg_q2052 AND symb_decoder(16#5a#)) OR
 					(reg_q2052 AND symb_decoder(16#3f#)) OR
 					(reg_q2052 AND symb_decoder(16#f8#)) OR
 					(reg_q2052 AND symb_decoder(16#8b#)) OR
 					(reg_q2052 AND symb_decoder(16#ac#)) OR
 					(reg_q2052 AND symb_decoder(16#f9#)) OR
 					(reg_q2052 AND symb_decoder(16#90#)) OR
 					(reg_q2052 AND symb_decoder(16#ad#)) OR
 					(reg_q2052 AND symb_decoder(16#93#)) OR
 					(reg_q2052 AND symb_decoder(16#0e#)) OR
 					(reg_q2052 AND symb_decoder(16#55#)) OR
 					(reg_q2052 AND symb_decoder(16#cb#)) OR
 					(reg_q2052 AND symb_decoder(16#42#)) OR
 					(reg_q2052 AND symb_decoder(16#09#)) OR
 					(reg_q2052 AND symb_decoder(16#8d#)) OR
 					(reg_q2052 AND symb_decoder(16#3e#)) OR
 					(reg_q2052 AND symb_decoder(16#66#)) OR
 					(reg_q2052 AND symb_decoder(16#f2#)) OR
 					(reg_q2052 AND symb_decoder(16#63#)) OR
 					(reg_q2052 AND symb_decoder(16#76#)) OR
 					(reg_q2052 AND symb_decoder(16#5f#)) OR
 					(reg_q2052 AND symb_decoder(16#95#)) OR
 					(reg_q2052 AND symb_decoder(16#05#)) OR
 					(reg_q2052 AND symb_decoder(16#0d#)) OR
 					(reg_q2052 AND symb_decoder(16#f0#)) OR
 					(reg_q2052 AND symb_decoder(16#c9#)) OR
 					(reg_q2052 AND symb_decoder(16#e5#)) OR
 					(reg_q2052 AND symb_decoder(16#f7#)) OR
 					(reg_q2052 AND symb_decoder(16#3a#)) OR
 					(reg_q2052 AND symb_decoder(16#fa#)) OR
 					(reg_q2052 AND symb_decoder(16#45#)) OR
 					(reg_q2052 AND symb_decoder(16#71#)) OR
 					(reg_q2052 AND symb_decoder(16#be#)) OR
 					(reg_q2052 AND symb_decoder(16#5d#)) OR
 					(reg_q2052 AND symb_decoder(16#5c#)) OR
 					(reg_q2052 AND symb_decoder(16#f6#)) OR
 					(reg_q2052 AND symb_decoder(16#12#)) OR
 					(reg_q2052 AND symb_decoder(16#59#)) OR
 					(reg_q2052 AND symb_decoder(16#b6#)) OR
 					(reg_q2052 AND symb_decoder(16#ca#)) OR
 					(reg_q2052 AND symb_decoder(16#a4#)) OR
 					(reg_q2052 AND symb_decoder(16#d1#)) OR
 					(reg_q2052 AND symb_decoder(16#c5#)) OR
 					(reg_q2052 AND symb_decoder(16#89#)) OR
 					(reg_q2052 AND symb_decoder(16#c6#)) OR
 					(reg_q2052 AND symb_decoder(16#8a#)) OR
 					(reg_q2052 AND symb_decoder(16#de#)) OR
 					(reg_q2052 AND symb_decoder(16#d9#)) OR
 					(reg_q2052 AND symb_decoder(16#a1#)) OR
 					(reg_q2052 AND symb_decoder(16#ee#)) OR
 					(reg_q2052 AND symb_decoder(16#da#)) OR
 					(reg_q2052 AND symb_decoder(16#b5#)) OR
 					(reg_q2052 AND symb_decoder(16#fe#)) OR
 					(reg_q2052 AND symb_decoder(16#1d#)) OR
 					(reg_q2052 AND symb_decoder(16#23#)) OR
 					(reg_q2052 AND symb_decoder(16#39#)) OR
 					(reg_q2052 AND symb_decoder(16#0f#)) OR
 					(reg_q2052 AND symb_decoder(16#15#)) OR
 					(reg_q2052 AND symb_decoder(16#86#)) OR
 					(reg_q2052 AND symb_decoder(16#e3#)) OR
 					(reg_q2052 AND symb_decoder(16#c3#)) OR
 					(reg_q2052 AND symb_decoder(16#df#)) OR
 					(reg_q2052 AND symb_decoder(16#d2#)) OR
 					(reg_q2052 AND symb_decoder(16#e4#)) OR
 					(reg_q2052 AND symb_decoder(16#57#)) OR
 					(reg_q2052 AND symb_decoder(16#e2#)) OR
 					(reg_q2052 AND symb_decoder(16#54#)) OR
 					(reg_q2052 AND symb_decoder(16#69#)) OR
 					(reg_q2052 AND symb_decoder(16#73#)) OR
 					(reg_q2052 AND symb_decoder(16#ce#)) OR
 					(reg_q2052 AND symb_decoder(16#a9#)) OR
 					(reg_q2052 AND symb_decoder(16#87#)) OR
 					(reg_q2052 AND symb_decoder(16#1a#)) OR
 					(reg_q2052 AND symb_decoder(16#9a#)) OR
 					(reg_q2052 AND symb_decoder(16#3c#)) OR
 					(reg_q2052 AND symb_decoder(16#2d#)) OR
 					(reg_q2052 AND symb_decoder(16#4f#)) OR
 					(reg_q2052 AND symb_decoder(16#e6#)) OR
 					(reg_q2052 AND symb_decoder(16#30#)) OR
 					(reg_q2052 AND symb_decoder(16#fc#)) OR
 					(reg_q2052 AND symb_decoder(16#25#)) OR
 					(reg_q2052 AND symb_decoder(16#ba#)) OR
 					(reg_q2052 AND symb_decoder(16#47#)) OR
 					(reg_q2052 AND symb_decoder(16#11#)) OR
 					(reg_q2052 AND symb_decoder(16#41#)) OR
 					(reg_q2052 AND symb_decoder(16#83#)) OR
 					(reg_q2052 AND symb_decoder(16#03#)) OR
 					(reg_q2052 AND symb_decoder(16#7c#)) OR
 					(reg_q2052 AND symb_decoder(16#26#)) OR
 					(reg_q2052 AND symb_decoder(16#d5#)) OR
 					(reg_q2052 AND symb_decoder(16#ab#)) OR
 					(reg_q2052 AND symb_decoder(16#cc#)) OR
 					(reg_q2052 AND symb_decoder(16#7f#)) OR
 					(reg_q2052 AND symb_decoder(16#9b#)) OR
 					(reg_q2052 AND symb_decoder(16#62#)) OR
 					(reg_q2052 AND symb_decoder(16#a8#)) OR
 					(reg_q2052 AND symb_decoder(16#6e#)) OR
 					(reg_q2052 AND symb_decoder(16#e8#)) OR
 					(reg_q2052 AND symb_decoder(16#20#)) OR
 					(reg_q2052 AND symb_decoder(16#cd#)) OR
 					(reg_q2052 AND symb_decoder(16#1c#)) OR
 					(reg_q2052 AND symb_decoder(16#91#)) OR
 					(reg_q2052 AND symb_decoder(16#2e#)) OR
 					(reg_q2052 AND symb_decoder(16#84#)) OR
 					(reg_q2052 AND symb_decoder(16#28#)) OR
 					(reg_q2052 AND symb_decoder(16#e1#)) OR
 					(reg_q2052 AND symb_decoder(16#04#)) OR
 					(reg_q2052 AND symb_decoder(16#9f#)) OR
 					(reg_q2052 AND symb_decoder(16#a6#)) OR
 					(reg_q2052 AND symb_decoder(16#ed#)) OR
 					(reg_q2052 AND symb_decoder(16#c2#)) OR
 					(reg_q2052 AND symb_decoder(16#18#)) OR
 					(reg_q2052 AND symb_decoder(16#bc#)) OR
 					(reg_q2052 AND symb_decoder(16#1b#)) OR
 					(reg_q2052 AND symb_decoder(16#82#)) OR
 					(reg_q2052 AND symb_decoder(16#bd#)) OR
 					(reg_q2052 AND symb_decoder(16#65#)) OR
 					(reg_q2052 AND symb_decoder(16#c7#)) OR
 					(reg_q2052 AND symb_decoder(16#0a#)) OR
 					(reg_q2052 AND symb_decoder(16#31#)) OR
 					(reg_q2052 AND symb_decoder(16#60#)) OR
 					(reg_q2052 AND symb_decoder(16#7a#)) OR
 					(reg_q2052 AND symb_decoder(16#77#)) OR
 					(reg_q2052 AND symb_decoder(16#24#)) OR
 					(reg_q2052 AND symb_decoder(16#7b#)) OR
 					(reg_q2052 AND symb_decoder(16#00#)) OR
 					(reg_q2052 AND symb_decoder(16#a2#)) OR
 					(reg_q2052 AND symb_decoder(16#b8#)) OR
 					(reg_q2052 AND symb_decoder(16#96#)) OR
 					(reg_q2052 AND symb_decoder(16#38#)) OR
 					(reg_q2052 AND symb_decoder(16#70#)) OR
 					(reg_q2052 AND symb_decoder(16#48#)) OR
 					(reg_q2052 AND symb_decoder(16#b0#)) OR
 					(reg_q2052 AND symb_decoder(16#10#)) OR
 					(reg_q2052 AND symb_decoder(16#61#)) OR
 					(reg_q2052 AND symb_decoder(16#b7#)) OR
 					(reg_q2052 AND symb_decoder(16#53#)) OR
 					(reg_q2052 AND symb_decoder(16#34#)) OR
 					(reg_q2052 AND symb_decoder(16#bb#)) OR
 					(reg_q2052 AND symb_decoder(16#6f#)) OR
 					(reg_q2052 AND symb_decoder(16#a0#)) OR
 					(reg_q2052 AND symb_decoder(16#19#)) OR
 					(reg_q2052 AND symb_decoder(16#2f#)) OR
 					(reg_q2052 AND symb_decoder(16#4a#)) OR
 					(reg_q2052 AND symb_decoder(16#44#)) OR
 					(reg_q2052 AND symb_decoder(16#13#)) OR
 					(reg_q2052 AND symb_decoder(16#97#)) OR
 					(reg_q2052 AND symb_decoder(16#75#)) OR
 					(reg_q2052 AND symb_decoder(16#af#)) OR
 					(reg_q2052 AND symb_decoder(16#72#)) OR
 					(reg_q2052 AND symb_decoder(16#74#)) OR
 					(reg_q2052 AND symb_decoder(16#98#)) OR
 					(reg_q2052 AND symb_decoder(16#40#)) OR
 					(reg_q2052 AND symb_decoder(16#88#)) OR
 					(reg_q2052 AND symb_decoder(16#79#)) OR
 					(reg_q2052 AND symb_decoder(16#e7#)) OR
 					(reg_q2052 AND symb_decoder(16#80#)) OR
 					(reg_q2052 AND symb_decoder(16#7d#)) OR
 					(reg_q2052 AND symb_decoder(16#78#)) OR
 					(reg_q2052 AND symb_decoder(16#d7#)) OR
 					(reg_q2052 AND symb_decoder(16#d3#)) OR
 					(reg_q2052 AND symb_decoder(16#f3#)) OR
 					(reg_q2052 AND symb_decoder(16#c0#)) OR
 					(reg_q2052 AND symb_decoder(16#eb#)) OR
 					(reg_q2052 AND symb_decoder(16#dc#)) OR
 					(reg_q2052 AND symb_decoder(16#f4#)) OR
 					(reg_q2052 AND symb_decoder(16#58#)) OR
 					(reg_q2052 AND symb_decoder(16#ec#)) OR
 					(reg_q2052 AND symb_decoder(16#0c#)) OR
 					(reg_q2052 AND symb_decoder(16#33#)) OR
 					(reg_q2052 AND symb_decoder(16#64#)) OR
 					(reg_q2052 AND symb_decoder(16#5b#)) OR
 					(reg_q2052 AND symb_decoder(16#1e#)) OR
 					(reg_q2052 AND symb_decoder(16#d0#)) OR
 					(reg_q2052 AND symb_decoder(16#aa#)) OR
 					(reg_q2052 AND symb_decoder(16#1f#)) OR
 					(reg_q2052 AND symb_decoder(16#29#)) OR
 					(reg_q2052 AND symb_decoder(16#9e#)) OR
 					(reg_q2052 AND symb_decoder(16#cf#)) OR
 					(reg_q2052 AND symb_decoder(16#14#)) OR
 					(reg_q2052 AND symb_decoder(16#2b#)) OR
 					(reg_q2052 AND symb_decoder(16#ea#)) OR
 					(reg_q2052 AND symb_decoder(16#5e#)) OR
 					(reg_q2052 AND symb_decoder(16#17#)) OR
 					(reg_q2052 AND symb_decoder(16#c4#)) OR
 					(reg_q2052 AND symb_decoder(16#3b#)) OR
 					(reg_q2052 AND symb_decoder(16#8c#)) OR
 					(reg_q2052 AND symb_decoder(16#08#)) OR
 					(reg_q2052 AND symb_decoder(16#99#)) OR
 					(reg_q2052 AND symb_decoder(16#37#)) OR
 					(reg_q2052 AND symb_decoder(16#4b#)) OR
 					(reg_q2052 AND symb_decoder(16#22#)) OR
 					(reg_q2052 AND symb_decoder(16#b2#)) OR
 					(reg_q2052 AND symb_decoder(16#7e#)) OR
 					(reg_q2052 AND symb_decoder(16#0b#)) OR
 					(reg_q2052 AND symb_decoder(16#c1#)) OR
 					(reg_q2052 AND symb_decoder(16#b3#)) OR
 					(reg_q2052 AND symb_decoder(16#4e#)) OR
 					(reg_q2052 AND symb_decoder(16#8e#)) OR
 					(reg_q2052 AND symb_decoder(16#16#)) OR
 					(reg_q2052 AND symb_decoder(16#dd#)) OR
 					(reg_q2052 AND symb_decoder(16#a7#)) OR
 					(reg_q2052 AND symb_decoder(16#32#)) OR
 					(reg_q2052 AND symb_decoder(16#f1#)) OR
 					(reg_q2052 AND symb_decoder(16#46#)) OR
 					(reg_q2052 AND symb_decoder(16#3d#)) OR
 					(reg_q2052 AND symb_decoder(16#6d#)) OR
 					(reg_q2052 AND symb_decoder(16#49#)) OR
 					(reg_q2052 AND symb_decoder(16#35#)) OR
 					(reg_q2052 AND symb_decoder(16#ef#)) OR
 					(reg_q2052 AND symb_decoder(16#50#)) OR
 					(reg_q2052 AND symb_decoder(16#b9#)) OR
 					(reg_q2052 AND symb_decoder(16#85#)) OR
 					(reg_q2052 AND symb_decoder(16#d6#)) OR
 					(reg_q2052 AND symb_decoder(16#21#)) OR
 					(reg_q2052 AND symb_decoder(16#8f#)) OR
 					(reg_q2052 AND symb_decoder(16#4c#)) OR
 					(reg_q2052 AND symb_decoder(16#b1#)) OR
 					(reg_q2052 AND symb_decoder(16#01#)) OR
 					(reg_q2052 AND symb_decoder(16#9d#)) OR
 					(reg_q2052 AND symb_decoder(16#6c#)) OR
 					(reg_q2052 AND symb_decoder(16#36#)) OR
 					(reg_q2052 AND symb_decoder(16#a5#)) OR
 					(reg_q2052 AND symb_decoder(16#f5#)) OR
 					(reg_q2052 AND symb_decoder(16#51#)) OR
 					(reg_q2052 AND symb_decoder(16#07#)) OR
 					(reg_q2052 AND symb_decoder(16#db#)) OR
 					(reg_q2052 AND symb_decoder(16#6a#)) OR
 					(reg_q2052 AND symb_decoder(16#fd#)) OR
 					(reg_q2052 AND symb_decoder(16#27#)) OR
 					(reg_q2052 AND symb_decoder(16#e9#)) OR
 					(reg_q2052 AND symb_decoder(16#2c#)) OR
 					(reg_q2052 AND symb_decoder(16#d4#)) OR
 					(reg_q2052 AND symb_decoder(16#43#)) OR
 					(reg_q2052 AND symb_decoder(16#ae#)) OR
 					(reg_q2052 AND symb_decoder(16#68#)) OR
 					(reg_q2052 AND symb_decoder(16#02#)) OR
 					(reg_q2052 AND symb_decoder(16#52#)) OR
 					(reg_q2052 AND symb_decoder(16#e0#)) OR
 					(reg_q2052 AND symb_decoder(16#6b#)) OR
 					(reg_q2052 AND symb_decoder(16#9c#)) OR
 					(reg_q2052 AND symb_decoder(16#81#)) OR
 					(reg_q2052 AND symb_decoder(16#94#));
reg_q2052_init <= '0' ;
	p_reg_q2052: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2052 <= reg_q2052_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2052 <= reg_q2052_init;
        else
          reg_q2052 <= reg_q2052_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q779_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q779 AND symb_decoder(16#5a#)) OR
 					(reg_q779 AND symb_decoder(16#df#)) OR
 					(reg_q779 AND symb_decoder(16#c5#)) OR
 					(reg_q779 AND symb_decoder(16#20#)) OR
 					(reg_q779 AND symb_decoder(16#74#)) OR
 					(reg_q779 AND symb_decoder(16#4a#)) OR
 					(reg_q779 AND symb_decoder(16#12#)) OR
 					(reg_q779 AND symb_decoder(16#5d#)) OR
 					(reg_q779 AND symb_decoder(16#bd#)) OR
 					(reg_q779 AND symb_decoder(16#41#)) OR
 					(reg_q779 AND symb_decoder(16#93#)) OR
 					(reg_q779 AND symb_decoder(16#a6#)) OR
 					(reg_q779 AND symb_decoder(16#92#)) OR
 					(reg_q779 AND symb_decoder(16#d1#)) OR
 					(reg_q779 AND symb_decoder(16#61#)) OR
 					(reg_q779 AND symb_decoder(16#3e#)) OR
 					(reg_q779 AND symb_decoder(16#ee#)) OR
 					(reg_q779 AND symb_decoder(16#bb#)) OR
 					(reg_q779 AND symb_decoder(16#6a#)) OR
 					(reg_q779 AND symb_decoder(16#84#)) OR
 					(reg_q779 AND symb_decoder(16#f7#)) OR
 					(reg_q779 AND symb_decoder(16#e2#)) OR
 					(reg_q779 AND symb_decoder(16#3a#)) OR
 					(reg_q779 AND symb_decoder(16#2f#)) OR
 					(reg_q779 AND symb_decoder(16#58#)) OR
 					(reg_q779 AND symb_decoder(16#9f#)) OR
 					(reg_q779 AND symb_decoder(16#75#)) OR
 					(reg_q779 AND symb_decoder(16#05#)) OR
 					(reg_q779 AND symb_decoder(16#7f#)) OR
 					(reg_q779 AND symb_decoder(16#fe#)) OR
 					(reg_q779 AND symb_decoder(16#85#)) OR
 					(reg_q779 AND symb_decoder(16#23#)) OR
 					(reg_q779 AND symb_decoder(16#ac#)) OR
 					(reg_q779 AND symb_decoder(16#9e#)) OR
 					(reg_q779 AND symb_decoder(16#45#)) OR
 					(reg_q779 AND symb_decoder(16#83#)) OR
 					(reg_q779 AND symb_decoder(16#97#)) OR
 					(reg_q779 AND symb_decoder(16#53#)) OR
 					(reg_q779 AND symb_decoder(16#f4#)) OR
 					(reg_q779 AND symb_decoder(16#70#)) OR
 					(reg_q779 AND symb_decoder(16#f9#)) OR
 					(reg_q779 AND symb_decoder(16#26#)) OR
 					(reg_q779 AND symb_decoder(16#d8#)) OR
 					(reg_q779 AND symb_decoder(16#24#)) OR
 					(reg_q779 AND symb_decoder(16#02#)) OR
 					(reg_q779 AND symb_decoder(16#0d#)) OR
 					(reg_q779 AND symb_decoder(16#aa#)) OR
 					(reg_q779 AND symb_decoder(16#d3#)) OR
 					(reg_q779 AND symb_decoder(16#48#)) OR
 					(reg_q779 AND symb_decoder(16#1d#)) OR
 					(reg_q779 AND symb_decoder(16#ef#)) OR
 					(reg_q779 AND symb_decoder(16#73#)) OR
 					(reg_q779 AND symb_decoder(16#a8#)) OR
 					(reg_q779 AND symb_decoder(16#30#)) OR
 					(reg_q779 AND symb_decoder(16#b8#)) OR
 					(reg_q779 AND symb_decoder(16#ce#)) OR
 					(reg_q779 AND symb_decoder(16#43#)) OR
 					(reg_q779 AND symb_decoder(16#44#)) OR
 					(reg_q779 AND symb_decoder(16#47#)) OR
 					(reg_q779 AND symb_decoder(16#c7#)) OR
 					(reg_q779 AND symb_decoder(16#c4#)) OR
 					(reg_q779 AND symb_decoder(16#b7#)) OR
 					(reg_q779 AND symb_decoder(16#bf#)) OR
 					(reg_q779 AND symb_decoder(16#56#)) OR
 					(reg_q779 AND symb_decoder(16#2a#)) OR
 					(reg_q779 AND symb_decoder(16#00#)) OR
 					(reg_q779 AND symb_decoder(16#a4#)) OR
 					(reg_q779 AND symb_decoder(16#cf#)) OR
 					(reg_q779 AND symb_decoder(16#7b#)) OR
 					(reg_q779 AND symb_decoder(16#0e#)) OR
 					(reg_q779 AND symb_decoder(16#38#)) OR
 					(reg_q779 AND symb_decoder(16#da#)) OR
 					(reg_q779 AND symb_decoder(16#77#)) OR
 					(reg_q779 AND symb_decoder(16#f5#)) OR
 					(reg_q779 AND symb_decoder(16#27#)) OR
 					(reg_q779 AND symb_decoder(16#4b#)) OR
 					(reg_q779 AND symb_decoder(16#76#)) OR
 					(reg_q779 AND symb_decoder(16#dd#)) OR
 					(reg_q779 AND symb_decoder(16#fb#)) OR
 					(reg_q779 AND symb_decoder(16#c6#)) OR
 					(reg_q779 AND symb_decoder(16#9b#)) OR
 					(reg_q779 AND symb_decoder(16#d2#)) OR
 					(reg_q779 AND symb_decoder(16#e1#)) OR
 					(reg_q779 AND symb_decoder(16#5c#)) OR
 					(reg_q779 AND symb_decoder(16#60#)) OR
 					(reg_q779 AND symb_decoder(16#29#)) OR
 					(reg_q779 AND symb_decoder(16#04#)) OR
 					(reg_q779 AND symb_decoder(16#dc#)) OR
 					(reg_q779 AND symb_decoder(16#49#)) OR
 					(reg_q779 AND symb_decoder(16#51#)) OR
 					(reg_q779 AND symb_decoder(16#36#)) OR
 					(reg_q779 AND symb_decoder(16#f8#)) OR
 					(reg_q779 AND symb_decoder(16#2b#)) OR
 					(reg_q779 AND symb_decoder(16#40#)) OR
 					(reg_q779 AND symb_decoder(16#c8#)) OR
 					(reg_q779 AND symb_decoder(16#17#)) OR
 					(reg_q779 AND symb_decoder(16#72#)) OR
 					(reg_q779 AND symb_decoder(16#b1#)) OR
 					(reg_q779 AND symb_decoder(16#f1#)) OR
 					(reg_q779 AND symb_decoder(16#f3#)) OR
 					(reg_q779 AND symb_decoder(16#79#)) OR
 					(reg_q779 AND symb_decoder(16#a7#)) OR
 					(reg_q779 AND symb_decoder(16#4e#)) OR
 					(reg_q779 AND symb_decoder(16#57#)) OR
 					(reg_q779 AND symb_decoder(16#5f#)) OR
 					(reg_q779 AND symb_decoder(16#80#)) OR
 					(reg_q779 AND symb_decoder(16#31#)) OR
 					(reg_q779 AND symb_decoder(16#3f#)) OR
 					(reg_q779 AND symb_decoder(16#d6#)) OR
 					(reg_q779 AND symb_decoder(16#d9#)) OR
 					(reg_q779 AND symb_decoder(16#65#)) OR
 					(reg_q779 AND symb_decoder(16#22#)) OR
 					(reg_q779 AND symb_decoder(16#9c#)) OR
 					(reg_q779 AND symb_decoder(16#71#)) OR
 					(reg_q779 AND symb_decoder(16#a2#)) OR
 					(reg_q779 AND symb_decoder(16#ab#)) OR
 					(reg_q779 AND symb_decoder(16#28#)) OR
 					(reg_q779 AND symb_decoder(16#86#)) OR
 					(reg_q779 AND symb_decoder(16#5e#)) OR
 					(reg_q779 AND symb_decoder(16#b3#)) OR
 					(reg_q779 AND symb_decoder(16#18#)) OR
 					(reg_q779 AND symb_decoder(16#39#)) OR
 					(reg_q779 AND symb_decoder(16#54#)) OR
 					(reg_q779 AND symb_decoder(16#cd#)) OR
 					(reg_q779 AND symb_decoder(16#b2#)) OR
 					(reg_q779 AND symb_decoder(16#1c#)) OR
 					(reg_q779 AND symb_decoder(16#e6#)) OR
 					(reg_q779 AND symb_decoder(16#ba#)) OR
 					(reg_q779 AND symb_decoder(16#78#)) OR
 					(reg_q779 AND symb_decoder(16#01#)) OR
 					(reg_q779 AND symb_decoder(16#e8#)) OR
 					(reg_q779 AND symb_decoder(16#90#)) OR
 					(reg_q779 AND symb_decoder(16#1a#)) OR
 					(reg_q779 AND symb_decoder(16#19#)) OR
 					(reg_q779 AND symb_decoder(16#16#)) OR
 					(reg_q779 AND symb_decoder(16#87#)) OR
 					(reg_q779 AND symb_decoder(16#a9#)) OR
 					(reg_q779 AND symb_decoder(16#c3#)) OR
 					(reg_q779 AND symb_decoder(16#34#)) OR
 					(reg_q779 AND symb_decoder(16#3d#)) OR
 					(reg_q779 AND symb_decoder(16#de#)) OR
 					(reg_q779 AND symb_decoder(16#ff#)) OR
 					(reg_q779 AND symb_decoder(16#11#)) OR
 					(reg_q779 AND symb_decoder(16#b6#)) OR
 					(reg_q779 AND symb_decoder(16#0a#)) OR
 					(reg_q779 AND symb_decoder(16#bc#)) OR
 					(reg_q779 AND symb_decoder(16#15#)) OR
 					(reg_q779 AND symb_decoder(16#68#)) OR
 					(reg_q779 AND symb_decoder(16#21#)) OR
 					(reg_q779 AND symb_decoder(16#8e#)) OR
 					(reg_q779 AND symb_decoder(16#a1#)) OR
 					(reg_q779 AND symb_decoder(16#2e#)) OR
 					(reg_q779 AND symb_decoder(16#5b#)) OR
 					(reg_q779 AND symb_decoder(16#4d#)) OR
 					(reg_q779 AND symb_decoder(16#8d#)) OR
 					(reg_q779 AND symb_decoder(16#8c#)) OR
 					(reg_q779 AND symb_decoder(16#f2#)) OR
 					(reg_q779 AND symb_decoder(16#91#)) OR
 					(reg_q779 AND symb_decoder(16#08#)) OR
 					(reg_q779 AND symb_decoder(16#cb#)) OR
 					(reg_q779 AND symb_decoder(16#8b#)) OR
 					(reg_q779 AND symb_decoder(16#55#)) OR
 					(reg_q779 AND symb_decoder(16#4f#)) OR
 					(reg_q779 AND symb_decoder(16#e4#)) OR
 					(reg_q779 AND symb_decoder(16#9d#)) OR
 					(reg_q779 AND symb_decoder(16#32#)) OR
 					(reg_q779 AND symb_decoder(16#63#)) OR
 					(reg_q779 AND symb_decoder(16#e3#)) OR
 					(reg_q779 AND symb_decoder(16#ed#)) OR
 					(reg_q779 AND symb_decoder(16#98#)) OR
 					(reg_q779 AND symb_decoder(16#64#)) OR
 					(reg_q779 AND symb_decoder(16#fd#)) OR
 					(reg_q779 AND symb_decoder(16#37#)) OR
 					(reg_q779 AND symb_decoder(16#d7#)) OR
 					(reg_q779 AND symb_decoder(16#e9#)) OR
 					(reg_q779 AND symb_decoder(16#52#)) OR
 					(reg_q779 AND symb_decoder(16#06#)) OR
 					(reg_q779 AND symb_decoder(16#96#)) OR
 					(reg_q779 AND symb_decoder(16#9a#)) OR
 					(reg_q779 AND symb_decoder(16#94#)) OR
 					(reg_q779 AND symb_decoder(16#88#)) OR
 					(reg_q779 AND symb_decoder(16#c2#)) OR
 					(reg_q779 AND symb_decoder(16#14#)) OR
 					(reg_q779 AND symb_decoder(16#d5#)) OR
 					(reg_q779 AND symb_decoder(16#69#)) OR
 					(reg_q779 AND symb_decoder(16#f0#)) OR
 					(reg_q779 AND symb_decoder(16#13#)) OR
 					(reg_q779 AND symb_decoder(16#a5#)) OR
 					(reg_q779 AND symb_decoder(16#ca#)) OR
 					(reg_q779 AND symb_decoder(16#35#)) OR
 					(reg_q779 AND symb_decoder(16#1e#)) OR
 					(reg_q779 AND symb_decoder(16#8f#)) OR
 					(reg_q779 AND symb_decoder(16#6f#)) OR
 					(reg_q779 AND symb_decoder(16#0c#)) OR
 					(reg_q779 AND symb_decoder(16#8a#)) OR
 					(reg_q779 AND symb_decoder(16#25#)) OR
 					(reg_q779 AND symb_decoder(16#a0#)) OR
 					(reg_q779 AND symb_decoder(16#2c#)) OR
 					(reg_q779 AND symb_decoder(16#ad#)) OR
 					(reg_q779 AND symb_decoder(16#b9#)) OR
 					(reg_q779 AND symb_decoder(16#6b#)) OR
 					(reg_q779 AND symb_decoder(16#ec#)) OR
 					(reg_q779 AND symb_decoder(16#81#)) OR
 					(reg_q779 AND symb_decoder(16#eb#)) OR
 					(reg_q779 AND symb_decoder(16#59#)) OR
 					(reg_q779 AND symb_decoder(16#99#)) OR
 					(reg_q779 AND symb_decoder(16#33#)) OR
 					(reg_q779 AND symb_decoder(16#89#)) OR
 					(reg_q779 AND symb_decoder(16#0b#)) OR
 					(reg_q779 AND symb_decoder(16#09#)) OR
 					(reg_q779 AND symb_decoder(16#fa#)) OR
 					(reg_q779 AND symb_decoder(16#ea#)) OR
 					(reg_q779 AND symb_decoder(16#3b#)) OR
 					(reg_q779 AND symb_decoder(16#46#)) OR
 					(reg_q779 AND symb_decoder(16#7c#)) OR
 					(reg_q779 AND symb_decoder(16#1b#)) OR
 					(reg_q779 AND symb_decoder(16#0f#)) OR
 					(reg_q779 AND symb_decoder(16#7e#)) OR
 					(reg_q779 AND symb_decoder(16#3c#)) OR
 					(reg_q779 AND symb_decoder(16#03#)) OR
 					(reg_q779 AND symb_decoder(16#fc#)) OR
 					(reg_q779 AND symb_decoder(16#c0#)) OR
 					(reg_q779 AND symb_decoder(16#b5#)) OR
 					(reg_q779 AND symb_decoder(16#95#)) OR
 					(reg_q779 AND symb_decoder(16#1f#)) OR
 					(reg_q779 AND symb_decoder(16#2d#)) OR
 					(reg_q779 AND symb_decoder(16#66#)) OR
 					(reg_q779 AND symb_decoder(16#4c#)) OR
 					(reg_q779 AND symb_decoder(16#10#)) OR
 					(reg_q779 AND symb_decoder(16#d0#)) OR
 					(reg_q779 AND symb_decoder(16#e0#)) OR
 					(reg_q779 AND symb_decoder(16#42#)) OR
 					(reg_q779 AND symb_decoder(16#7d#)) OR
 					(reg_q779 AND symb_decoder(16#f6#)) OR
 					(reg_q779 AND symb_decoder(16#50#)) OR
 					(reg_q779 AND symb_decoder(16#e5#)) OR
 					(reg_q779 AND symb_decoder(16#cc#)) OR
 					(reg_q779 AND symb_decoder(16#82#)) OR
 					(reg_q779 AND symb_decoder(16#07#)) OR
 					(reg_q779 AND symb_decoder(16#d4#)) OR
 					(reg_q779 AND symb_decoder(16#af#)) OR
 					(reg_q779 AND symb_decoder(16#62#)) OR
 					(reg_q779 AND symb_decoder(16#c9#)) OR
 					(reg_q779 AND symb_decoder(16#6c#)) OR
 					(reg_q779 AND symb_decoder(16#e7#)) OR
 					(reg_q779 AND symb_decoder(16#c1#)) OR
 					(reg_q779 AND symb_decoder(16#db#)) OR
 					(reg_q779 AND symb_decoder(16#a3#)) OR
 					(reg_q779 AND symb_decoder(16#6e#)) OR
 					(reg_q779 AND symb_decoder(16#ae#)) OR
 					(reg_q779 AND symb_decoder(16#67#)) OR
 					(reg_q779 AND symb_decoder(16#be#)) OR
 					(reg_q779 AND symb_decoder(16#6d#)) OR
 					(reg_q779 AND symb_decoder(16#b4#)) OR
 					(reg_q779 AND symb_decoder(16#b0#)) OR
 					(reg_q779 AND symb_decoder(16#7a#));
reg_q779_init <= '0' ;
	p_reg_q779: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q779 <= reg_q779_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q779 <= reg_q779_init;
        else
          reg_q779 <= reg_q779_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q91_in <= (reg_q2695 AND symb_decoder(16#f5#)) OR
 					(reg_q2695 AND symb_decoder(16#b3#)) OR
 					(reg_q2695 AND symb_decoder(16#ea#)) OR
 					(reg_q2695 AND symb_decoder(16#d7#)) OR
 					(reg_q2695 AND symb_decoder(16#d5#)) OR
 					(reg_q2695 AND symb_decoder(16#a4#)) OR
 					(reg_q2695 AND symb_decoder(16#49#)) OR
 					(reg_q2695 AND symb_decoder(16#85#)) OR
 					(reg_q2695 AND symb_decoder(16#3a#)) OR
 					(reg_q2695 AND symb_decoder(16#2c#)) OR
 					(reg_q2695 AND symb_decoder(16#c1#)) OR
 					(reg_q2695 AND symb_decoder(16#ba#)) OR
 					(reg_q2695 AND symb_decoder(16#0f#)) OR
 					(reg_q2695 AND symb_decoder(16#df#)) OR
 					(reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#e8#)) OR
 					(reg_q2695 AND symb_decoder(16#2d#)) OR
 					(reg_q2695 AND symb_decoder(16#bf#)) OR
 					(reg_q2695 AND symb_decoder(16#7a#)) OR
 					(reg_q2695 AND symb_decoder(16#31#)) OR
 					(reg_q2695 AND symb_decoder(16#97#)) OR
 					(reg_q2695 AND symb_decoder(16#93#)) OR
 					(reg_q2695 AND symb_decoder(16#11#)) OR
 					(reg_q2695 AND symb_decoder(16#1d#)) OR
 					(reg_q2695 AND symb_decoder(16#6f#)) OR
 					(reg_q2695 AND symb_decoder(16#f6#)) OR
 					(reg_q2695 AND symb_decoder(16#50#)) OR
 					(reg_q2695 AND symb_decoder(16#de#)) OR
 					(reg_q2695 AND symb_decoder(16#1f#)) OR
 					(reg_q2695 AND symb_decoder(16#6c#)) OR
 					(reg_q2695 AND symb_decoder(16#59#)) OR
 					(reg_q2695 AND symb_decoder(16#39#)) OR
 					(reg_q2695 AND symb_decoder(16#7d#)) OR
 					(reg_q2695 AND symb_decoder(16#d2#)) OR
 					(reg_q2695 AND symb_decoder(16#27#)) OR
 					(reg_q2695 AND symb_decoder(16#2f#)) OR
 					(reg_q2695 AND symb_decoder(16#8d#)) OR
 					(reg_q2695 AND symb_decoder(16#a7#)) OR
 					(reg_q2695 AND symb_decoder(16#e2#)) OR
 					(reg_q2695 AND symb_decoder(16#c3#)) OR
 					(reg_q2695 AND symb_decoder(16#67#)) OR
 					(reg_q2695 AND symb_decoder(16#38#)) OR
 					(reg_q2695 AND symb_decoder(16#ad#)) OR
 					(reg_q2695 AND symb_decoder(16#cc#)) OR
 					(reg_q2695 AND symb_decoder(16#01#)) OR
 					(reg_q2695 AND symb_decoder(16#ec#)) OR
 					(reg_q2695 AND symb_decoder(16#15#)) OR
 					(reg_q2695 AND symb_decoder(16#c5#)) OR
 					(reg_q2695 AND symb_decoder(16#ef#)) OR
 					(reg_q2695 AND symb_decoder(16#e5#)) OR
 					(reg_q2695 AND symb_decoder(16#a9#)) OR
 					(reg_q2695 AND symb_decoder(16#6e#)) OR
 					(reg_q2695 AND symb_decoder(16#4a#)) OR
 					(reg_q2695 AND symb_decoder(16#9c#)) OR
 					(reg_q2695 AND symb_decoder(16#9f#)) OR
 					(reg_q2695 AND symb_decoder(16#54#)) OR
 					(reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#cd#)) OR
 					(reg_q2695 AND symb_decoder(16#63#)) OR
 					(reg_q2695 AND symb_decoder(16#dd#)) OR
 					(reg_q2695 AND symb_decoder(16#19#)) OR
 					(reg_q2695 AND symb_decoder(16#d1#)) OR
 					(reg_q2695 AND symb_decoder(16#72#)) OR
 					(reg_q2695 AND symb_decoder(16#7f#)) OR
 					(reg_q2695 AND symb_decoder(16#75#)) OR
 					(reg_q2695 AND symb_decoder(16#08#)) OR
 					(reg_q2695 AND symb_decoder(16#1c#)) OR
 					(reg_q2695 AND symb_decoder(16#6d#)) OR
 					(reg_q2695 AND symb_decoder(16#f8#)) OR
 					(reg_q2695 AND symb_decoder(16#16#)) OR
 					(reg_q2695 AND symb_decoder(16#35#)) OR
 					(reg_q2695 AND symb_decoder(16#e7#)) OR
 					(reg_q2695 AND symb_decoder(16#ce#)) OR
 					(reg_q2695 AND symb_decoder(16#b2#)) OR
 					(reg_q2695 AND symb_decoder(16#14#)) OR
 					(reg_q2695 AND symb_decoder(16#6b#)) OR
 					(reg_q2695 AND symb_decoder(16#7c#)) OR
 					(reg_q2695 AND symb_decoder(16#e9#)) OR
 					(reg_q2695 AND symb_decoder(16#2b#)) OR
 					(reg_q2695 AND symb_decoder(16#d4#)) OR
 					(reg_q2695 AND symb_decoder(16#ab#)) OR
 					(reg_q2695 AND symb_decoder(16#5a#)) OR
 					(reg_q2695 AND symb_decoder(16#82#)) OR
 					(reg_q2695 AND symb_decoder(16#5f#)) OR
 					(reg_q2695 AND symb_decoder(16#a5#)) OR
 					(reg_q2695 AND symb_decoder(16#83#)) OR
 					(reg_q2695 AND symb_decoder(16#37#)) OR
 					(reg_q2695 AND symb_decoder(16#84#)) OR
 					(reg_q2695 AND symb_decoder(16#87#)) OR
 					(reg_q2695 AND symb_decoder(16#fa#)) OR
 					(reg_q2695 AND symb_decoder(16#04#)) OR
 					(reg_q2695 AND symb_decoder(16#9b#)) OR
 					(reg_q2695 AND symb_decoder(16#55#)) OR
 					(reg_q2695 AND symb_decoder(16#1a#)) OR
 					(reg_q2695 AND symb_decoder(16#c8#)) OR
 					(reg_q2695 AND symb_decoder(16#58#)) OR
 					(reg_q2695 AND symb_decoder(16#b9#)) OR
 					(reg_q2695 AND symb_decoder(16#db#)) OR
 					(reg_q2695 AND symb_decoder(16#cf#)) OR
 					(reg_q2695 AND symb_decoder(16#0e#)) OR
 					(reg_q2695 AND symb_decoder(16#76#)) OR
 					(reg_q2695 AND symb_decoder(16#06#)) OR
 					(reg_q2695 AND symb_decoder(16#9e#)) OR
 					(reg_q2695 AND symb_decoder(16#9a#)) OR
 					(reg_q2695 AND symb_decoder(16#d6#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q2695 AND symb_decoder(16#23#)) OR
 					(reg_q2695 AND symb_decoder(16#43#)) OR
 					(reg_q2695 AND symb_decoder(16#bd#)) OR
 					(reg_q2695 AND symb_decoder(16#8f#)) OR
 					(reg_q2695 AND symb_decoder(16#1e#)) OR
 					(reg_q2695 AND symb_decoder(16#61#)) OR
 					(reg_q2695 AND symb_decoder(16#f2#)) OR
 					(reg_q2695 AND symb_decoder(16#5e#)) OR
 					(reg_q2695 AND symb_decoder(16#86#)) OR
 					(reg_q2695 AND symb_decoder(16#a3#)) OR
 					(reg_q2695 AND symb_decoder(16#fd#)) OR
 					(reg_q2695 AND symb_decoder(16#ff#)) OR
 					(reg_q2695 AND symb_decoder(16#17#)) OR
 					(reg_q2695 AND symb_decoder(16#2a#)) OR
 					(reg_q2695 AND symb_decoder(16#5b#)) OR
 					(reg_q2695 AND symb_decoder(16#28#)) OR
 					(reg_q2695 AND symb_decoder(16#3f#)) OR
 					(reg_q2695 AND symb_decoder(16#89#)) OR
 					(reg_q2695 AND symb_decoder(16#6a#)) OR
 					(reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#00#)) OR
 					(reg_q2695 AND symb_decoder(16#c7#)) OR
 					(reg_q2695 AND symb_decoder(16#4c#)) OR
 					(reg_q2695 AND symb_decoder(16#03#)) OR
 					(reg_q2695 AND symb_decoder(16#57#)) OR
 					(reg_q2695 AND symb_decoder(16#d8#)) OR
 					(reg_q2695 AND symb_decoder(16#eb#)) OR
 					(reg_q2695 AND symb_decoder(16#a2#)) OR
 					(reg_q2695 AND symb_decoder(16#1b#)) OR
 					(reg_q2695 AND symb_decoder(16#b1#)) OR
 					(reg_q2695 AND symb_decoder(16#b0#)) OR
 					(reg_q2695 AND symb_decoder(16#12#)) OR
 					(reg_q2695 AND symb_decoder(16#05#)) OR
 					(reg_q2695 AND symb_decoder(16#7b#)) OR
 					(reg_q2695 AND symb_decoder(16#c6#)) OR
 					(reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#45#)) OR
 					(reg_q2695 AND symb_decoder(16#91#)) OR
 					(reg_q2695 AND symb_decoder(16#21#)) OR
 					(reg_q2695 AND symb_decoder(16#7e#)) OR
 					(reg_q2695 AND symb_decoder(16#a1#)) OR
 					(reg_q2695 AND symb_decoder(16#c0#)) OR
 					(reg_q2695 AND symb_decoder(16#4f#)) OR
 					(reg_q2695 AND symb_decoder(16#48#)) OR
 					(reg_q2695 AND symb_decoder(16#fc#)) OR
 					(reg_q2695 AND symb_decoder(16#44#)) OR
 					(reg_q2695 AND symb_decoder(16#4b#)) OR
 					(reg_q2695 AND symb_decoder(16#d0#)) OR
 					(reg_q2695 AND symb_decoder(16#40#)) OR
 					(reg_q2695 AND symb_decoder(16#34#)) OR
 					(reg_q2695 AND symb_decoder(16#ca#)) OR
 					(reg_q2695 AND symb_decoder(16#81#)) OR
 					(reg_q2695 AND symb_decoder(16#70#)) OR
 					(reg_q2695 AND symb_decoder(16#b8#)) OR
 					(reg_q2695 AND symb_decoder(16#bb#)) OR
 					(reg_q2695 AND symb_decoder(16#a0#)) OR
 					(reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q2695 AND symb_decoder(16#60#)) OR
 					(reg_q2695 AND symb_decoder(16#13#)) OR
 					(reg_q2695 AND symb_decoder(16#e0#)) OR
 					(reg_q2695 AND symb_decoder(16#94#)) OR
 					(reg_q2695 AND symb_decoder(16#e1#)) OR
 					(reg_q2695 AND symb_decoder(16#ed#)) OR
 					(reg_q2695 AND symb_decoder(16#41#)) OR
 					(reg_q2695 AND symb_decoder(16#b4#)) OR
 					(reg_q2695 AND symb_decoder(16#be#)) OR
 					(reg_q2695 AND symb_decoder(16#e3#)) OR
 					(reg_q2695 AND symb_decoder(16#25#)) OR
 					(reg_q2695 AND symb_decoder(16#02#)) OR
 					(reg_q2695 AND symb_decoder(16#22#)) OR
 					(reg_q2695 AND symb_decoder(16#36#)) OR
 					(reg_q2695 AND symb_decoder(16#52#)) OR
 					(reg_q2695 AND symb_decoder(16#ae#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#c2#)) OR
 					(reg_q2695 AND symb_decoder(16#26#)) OR
 					(reg_q2695 AND symb_decoder(16#c9#)) OR
 					(reg_q2695 AND symb_decoder(16#f9#)) OR
 					(reg_q2695 AND symb_decoder(16#8a#)) OR
 					(reg_q2695 AND symb_decoder(16#4d#)) OR
 					(reg_q2695 AND symb_decoder(16#3d#)) OR
 					(reg_q2695 AND symb_decoder(16#bc#)) OR
 					(reg_q2695 AND symb_decoder(16#dc#)) OR
 					(reg_q2695 AND symb_decoder(16#f7#)) OR
 					(reg_q2695 AND symb_decoder(16#8c#)) OR
 					(reg_q2695 AND symb_decoder(16#aa#)) OR
 					(reg_q2695 AND symb_decoder(16#f3#)) OR
 					(reg_q2695 AND symb_decoder(16#77#)) OR
 					(reg_q2695 AND symb_decoder(16#ac#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#95#)) OR
 					(reg_q2695 AND symb_decoder(16#98#)) OR
 					(reg_q2695 AND symb_decoder(16#b7#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q2695 AND symb_decoder(16#51#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q2695 AND symb_decoder(16#e6#)) OR
 					(reg_q2695 AND symb_decoder(16#4e#)) OR
 					(reg_q2695 AND symb_decoder(16#e4#)) OR
 					(reg_q2695 AND symb_decoder(16#74#)) OR
 					(reg_q2695 AND symb_decoder(16#71#)) OR
 					(reg_q2695 AND symb_decoder(16#a6#)) OR
 					(reg_q2695 AND symb_decoder(16#f4#)) OR
 					(reg_q2695 AND symb_decoder(16#2e#)) OR
 					(reg_q2695 AND symb_decoder(16#5d#)) OR
 					(reg_q2695 AND symb_decoder(16#64#)) OR
 					(reg_q2695 AND symb_decoder(16#78#)) OR
 					(reg_q2695 AND symb_decoder(16#80#)) OR
 					(reg_q2695 AND symb_decoder(16#fb#)) OR
 					(reg_q2695 AND symb_decoder(16#29#)) OR
 					(reg_q2695 AND symb_decoder(16#b5#)) OR
 					(reg_q2695 AND symb_decoder(16#24#)) OR
 					(reg_q2695 AND symb_decoder(16#88#)) OR
 					(reg_q2695 AND symb_decoder(16#f1#)) OR
 					(reg_q2695 AND symb_decoder(16#fe#)) OR
 					(reg_q2695 AND symb_decoder(16#92#)) OR
 					(reg_q2695 AND symb_decoder(16#68#)) OR
 					(reg_q2695 AND symb_decoder(16#ee#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q2695 AND symb_decoder(16#af#)) OR
 					(reg_q2695 AND symb_decoder(16#33#)) OR
 					(reg_q2695 AND symb_decoder(16#8e#)) OR
 					(reg_q2695 AND symb_decoder(16#8b#)) OR
 					(reg_q2695 AND symb_decoder(16#79#)) OR
 					(reg_q2695 AND symb_decoder(16#07#)) OR
 					(reg_q2695 AND symb_decoder(16#32#)) OR
 					(reg_q2695 AND symb_decoder(16#5c#)) OR
 					(reg_q2695 AND symb_decoder(16#a8#)) OR
 					(reg_q2695 AND symb_decoder(16#56#)) OR
 					(reg_q2695 AND symb_decoder(16#10#)) OR
 					(reg_q2695 AND symb_decoder(16#3e#)) OR
 					(reg_q2695 AND symb_decoder(16#cb#)) OR
 					(reg_q2695 AND symb_decoder(16#b6#)) OR
 					(reg_q2695 AND symb_decoder(16#3c#)) OR
 					(reg_q2695 AND symb_decoder(16#90#)) OR
 					(reg_q2695 AND symb_decoder(16#9d#)) OR
 					(reg_q2695 AND symb_decoder(16#3b#)) OR
 					(reg_q2695 AND symb_decoder(16#65#)) OR
 					(reg_q2695 AND symb_decoder(16#99#)) OR
 					(reg_q2695 AND symb_decoder(16#d9#)) OR
 					(reg_q2695 AND symb_decoder(16#0b#)) OR
 					(reg_q2695 AND symb_decoder(16#f0#)) OR
 					(reg_q2695 AND symb_decoder(16#18#)) OR
 					(reg_q2695 AND symb_decoder(16#c4#)) OR
 					(reg_q2695 AND symb_decoder(16#69#)) OR
 					(reg_q2695 AND symb_decoder(16#96#)) OR
 					(reg_q2695 AND symb_decoder(16#d3#)) OR
 					(reg_q2695 AND symb_decoder(16#da#)) OR
 					(reg_q2695 AND symb_decoder(16#47#)) OR
 					(reg_q91 AND symb_decoder(16#af#)) OR
 					(reg_q91 AND symb_decoder(16#2f#)) OR
 					(reg_q91 AND symb_decoder(16#46#)) OR
 					(reg_q91 AND symb_decoder(16#ac#)) OR
 					(reg_q91 AND symb_decoder(16#05#)) OR
 					(reg_q91 AND symb_decoder(16#e5#)) OR
 					(reg_q91 AND symb_decoder(16#c6#)) OR
 					(reg_q91 AND symb_decoder(16#d6#)) OR
 					(reg_q91 AND symb_decoder(16#6b#)) OR
 					(reg_q91 AND symb_decoder(16#35#)) OR
 					(reg_q91 AND symb_decoder(16#94#)) OR
 					(reg_q91 AND symb_decoder(16#d5#)) OR
 					(reg_q91 AND symb_decoder(16#12#)) OR
 					(reg_q91 AND symb_decoder(16#68#)) OR
 					(reg_q91 AND symb_decoder(16#ce#)) OR
 					(reg_q91 AND symb_decoder(16#fc#)) OR
 					(reg_q91 AND symb_decoder(16#01#)) OR
 					(reg_q91 AND symb_decoder(16#8e#)) OR
 					(reg_q91 AND symb_decoder(16#73#)) OR
 					(reg_q91 AND symb_decoder(16#b4#)) OR
 					(reg_q91 AND symb_decoder(16#1d#)) OR
 					(reg_q91 AND symb_decoder(16#b3#)) OR
 					(reg_q91 AND symb_decoder(16#a8#)) OR
 					(reg_q91 AND symb_decoder(16#d1#)) OR
 					(reg_q91 AND symb_decoder(16#a4#)) OR
 					(reg_q91 AND symb_decoder(16#25#)) OR
 					(reg_q91 AND symb_decoder(16#5e#)) OR
 					(reg_q91 AND symb_decoder(16#5f#)) OR
 					(reg_q91 AND symb_decoder(16#56#)) OR
 					(reg_q91 AND symb_decoder(16#17#)) OR
 					(reg_q91 AND symb_decoder(16#76#)) OR
 					(reg_q91 AND symb_decoder(16#f5#)) OR
 					(reg_q91 AND symb_decoder(16#0b#)) OR
 					(reg_q91 AND symb_decoder(16#39#)) OR
 					(reg_q91 AND symb_decoder(16#8f#)) OR
 					(reg_q91 AND symb_decoder(16#6a#)) OR
 					(reg_q91 AND symb_decoder(16#3e#)) OR
 					(reg_q91 AND symb_decoder(16#a2#)) OR
 					(reg_q91 AND symb_decoder(16#78#)) OR
 					(reg_q91 AND symb_decoder(16#a0#)) OR
 					(reg_q91 AND symb_decoder(16#5a#)) OR
 					(reg_q91 AND symb_decoder(16#58#)) OR
 					(reg_q91 AND symb_decoder(16#7d#)) OR
 					(reg_q91 AND symb_decoder(16#47#)) OR
 					(reg_q91 AND symb_decoder(16#3a#)) OR
 					(reg_q91 AND symb_decoder(16#2c#)) OR
 					(reg_q91 AND symb_decoder(16#96#)) OR
 					(reg_q91 AND symb_decoder(16#45#)) OR
 					(reg_q91 AND symb_decoder(16#9f#)) OR
 					(reg_q91 AND symb_decoder(16#6e#)) OR
 					(reg_q91 AND symb_decoder(16#93#)) OR
 					(reg_q91 AND symb_decoder(16#c1#)) OR
 					(reg_q91 AND symb_decoder(16#d7#)) OR
 					(reg_q91 AND symb_decoder(16#3c#)) OR
 					(reg_q91 AND symb_decoder(16#71#)) OR
 					(reg_q91 AND symb_decoder(16#53#)) OR
 					(reg_q91 AND symb_decoder(16#1e#)) OR
 					(reg_q91 AND symb_decoder(16#cb#)) OR
 					(reg_q91 AND symb_decoder(16#4a#)) OR
 					(reg_q91 AND symb_decoder(16#f1#)) OR
 					(reg_q91 AND symb_decoder(16#36#)) OR
 					(reg_q91 AND symb_decoder(16#20#)) OR
 					(reg_q91 AND symb_decoder(16#04#)) OR
 					(reg_q91 AND symb_decoder(16#0f#)) OR
 					(reg_q91 AND symb_decoder(16#c7#)) OR
 					(reg_q91 AND symb_decoder(16#21#)) OR
 					(reg_q91 AND symb_decoder(16#99#)) OR
 					(reg_q91 AND symb_decoder(16#cc#)) OR
 					(reg_q91 AND symb_decoder(16#d3#)) OR
 					(reg_q91 AND symb_decoder(16#87#)) OR
 					(reg_q91 AND symb_decoder(16#ba#)) OR
 					(reg_q91 AND symb_decoder(16#6d#)) OR
 					(reg_q91 AND symb_decoder(16#bc#)) OR
 					(reg_q91 AND symb_decoder(16#24#)) OR
 					(reg_q91 AND symb_decoder(16#b0#)) OR
 					(reg_q91 AND symb_decoder(16#f3#)) OR
 					(reg_q91 AND symb_decoder(16#c2#)) OR
 					(reg_q91 AND symb_decoder(16#d8#)) OR
 					(reg_q91 AND symb_decoder(16#c5#)) OR
 					(reg_q91 AND symb_decoder(16#db#)) OR
 					(reg_q91 AND symb_decoder(16#0e#)) OR
 					(reg_q91 AND symb_decoder(16#2d#)) OR
 					(reg_q91 AND symb_decoder(16#07#)) OR
 					(reg_q91 AND symb_decoder(16#79#)) OR
 					(reg_q91 AND symb_decoder(16#03#)) OR
 					(reg_q91 AND symb_decoder(16#65#)) OR
 					(reg_q91 AND symb_decoder(16#d4#)) OR
 					(reg_q91 AND symb_decoder(16#ec#)) OR
 					(reg_q91 AND symb_decoder(16#9d#)) OR
 					(reg_q91 AND symb_decoder(16#55#)) OR
 					(reg_q91 AND symb_decoder(16#9b#)) OR
 					(reg_q91 AND symb_decoder(16#19#)) OR
 					(reg_q91 AND symb_decoder(16#83#)) OR
 					(reg_q91 AND symb_decoder(16#2b#)) OR
 					(reg_q91 AND symb_decoder(16#2e#)) OR
 					(reg_q91 AND symb_decoder(16#ef#)) OR
 					(reg_q91 AND symb_decoder(16#cf#)) OR
 					(reg_q91 AND symb_decoder(16#0c#)) OR
 					(reg_q91 AND symb_decoder(16#ea#)) OR
 					(reg_q91 AND symb_decoder(16#e9#)) OR
 					(reg_q91 AND symb_decoder(16#c4#)) OR
 					(reg_q91 AND symb_decoder(16#5c#)) OR
 					(reg_q91 AND symb_decoder(16#22#)) OR
 					(reg_q91 AND symb_decoder(16#3d#)) OR
 					(reg_q91 AND symb_decoder(16#a9#)) OR
 					(reg_q91 AND symb_decoder(16#0a#)) OR
 					(reg_q91 AND symb_decoder(16#66#)) OR
 					(reg_q91 AND symb_decoder(16#54#)) OR
 					(reg_q91 AND symb_decoder(16#cd#)) OR
 					(reg_q91 AND symb_decoder(16#dd#)) OR
 					(reg_q91 AND symb_decoder(16#1f#)) OR
 					(reg_q91 AND symb_decoder(16#0d#)) OR
 					(reg_q91 AND symb_decoder(16#1a#)) OR
 					(reg_q91 AND symb_decoder(16#f2#)) OR
 					(reg_q91 AND symb_decoder(16#13#)) OR
 					(reg_q91 AND symb_decoder(16#3b#)) OR
 					(reg_q91 AND symb_decoder(16#9a#)) OR
 					(reg_q91 AND symb_decoder(16#eb#)) OR
 					(reg_q91 AND symb_decoder(16#b8#)) OR
 					(reg_q91 AND symb_decoder(16#08#)) OR
 					(reg_q91 AND symb_decoder(16#02#)) OR
 					(reg_q91 AND symb_decoder(16#52#)) OR
 					(reg_q91 AND symb_decoder(16#89#)) OR
 					(reg_q91 AND symb_decoder(16#49#)) OR
 					(reg_q91 AND symb_decoder(16#63#)) OR
 					(reg_q91 AND symb_decoder(16#50#)) OR
 					(reg_q91 AND symb_decoder(16#1b#)) OR
 					(reg_q91 AND symb_decoder(16#b1#)) OR
 					(reg_q91 AND symb_decoder(16#48#)) OR
 					(reg_q91 AND symb_decoder(16#4f#)) OR
 					(reg_q91 AND symb_decoder(16#14#)) OR
 					(reg_q91 AND symb_decoder(16#e7#)) OR
 					(reg_q91 AND symb_decoder(16#c8#)) OR
 					(reg_q91 AND symb_decoder(16#ab#)) OR
 					(reg_q91 AND symb_decoder(16#bd#)) OR
 					(reg_q91 AND symb_decoder(16#4e#)) OR
 					(reg_q91 AND symb_decoder(16#1c#)) OR
 					(reg_q91 AND symb_decoder(16#23#)) OR
 					(reg_q91 AND symb_decoder(16#92#)) OR
 					(reg_q91 AND symb_decoder(16#6c#)) OR
 					(reg_q91 AND symb_decoder(16#7b#)) OR
 					(reg_q91 AND symb_decoder(16#29#)) OR
 					(reg_q91 AND symb_decoder(16#a3#)) OR
 					(reg_q91 AND symb_decoder(16#75#)) OR
 					(reg_q91 AND symb_decoder(16#e1#)) OR
 					(reg_q91 AND symb_decoder(16#7f#)) OR
 					(reg_q91 AND symb_decoder(16#34#)) OR
 					(reg_q91 AND symb_decoder(16#df#)) OR
 					(reg_q91 AND symb_decoder(16#38#)) OR
 					(reg_q91 AND symb_decoder(16#90#)) OR
 					(reg_q91 AND symb_decoder(16#41#)) OR
 					(reg_q91 AND symb_decoder(16#43#)) OR
 					(reg_q91 AND symb_decoder(16#72#)) OR
 					(reg_q91 AND symb_decoder(16#a7#)) OR
 					(reg_q91 AND symb_decoder(16#be#)) OR
 					(reg_q91 AND symb_decoder(16#b2#)) OR
 					(reg_q91 AND symb_decoder(16#95#)) OR
 					(reg_q91 AND symb_decoder(16#e8#)) OR
 					(reg_q91 AND symb_decoder(16#7a#)) OR
 					(reg_q91 AND symb_decoder(16#b6#)) OR
 					(reg_q91 AND symb_decoder(16#97#)) OR
 					(reg_q91 AND symb_decoder(16#18#)) OR
 					(reg_q91 AND symb_decoder(16#f8#)) OR
 					(reg_q91 AND symb_decoder(16#5d#)) OR
 					(reg_q91 AND symb_decoder(16#ff#)) OR
 					(reg_q91 AND symb_decoder(16#bf#)) OR
 					(reg_q91 AND symb_decoder(16#10#)) OR
 					(reg_q91 AND symb_decoder(16#11#)) OR
 					(reg_q91 AND symb_decoder(16#7c#)) OR
 					(reg_q91 AND symb_decoder(16#d9#)) OR
 					(reg_q91 AND symb_decoder(16#fa#)) OR
 					(reg_q91 AND symb_decoder(16#e6#)) OR
 					(reg_q91 AND symb_decoder(16#86#)) OR
 					(reg_q91 AND symb_decoder(16#b9#)) OR
 					(reg_q91 AND symb_decoder(16#8d#)) OR
 					(reg_q91 AND symb_decoder(16#37#)) OR
 					(reg_q91 AND symb_decoder(16#64#)) OR
 					(reg_q91 AND symb_decoder(16#33#)) OR
 					(reg_q91 AND symb_decoder(16#f6#)) OR
 					(reg_q91 AND symb_decoder(16#7e#)) OR
 					(reg_q91 AND symb_decoder(16#44#)) OR
 					(reg_q91 AND symb_decoder(16#00#)) OR
 					(reg_q91 AND symb_decoder(16#f7#)) OR
 					(reg_q91 AND symb_decoder(16#57#)) OR
 					(reg_q91 AND symb_decoder(16#06#)) OR
 					(reg_q91 AND symb_decoder(16#a1#)) OR
 					(reg_q91 AND symb_decoder(16#27#)) OR
 					(reg_q91 AND symb_decoder(16#f9#)) OR
 					(reg_q91 AND symb_decoder(16#9e#)) OR
 					(reg_q91 AND symb_decoder(16#ee#)) OR
 					(reg_q91 AND symb_decoder(16#5b#)) OR
 					(reg_q91 AND symb_decoder(16#84#)) OR
 					(reg_q91 AND symb_decoder(16#a6#)) OR
 					(reg_q91 AND symb_decoder(16#81#)) OR
 					(reg_q91 AND symb_decoder(16#8c#)) OR
 					(reg_q91 AND symb_decoder(16#88#)) OR
 					(reg_q91 AND symb_decoder(16#67#)) OR
 					(reg_q91 AND symb_decoder(16#32#)) OR
 					(reg_q91 AND symb_decoder(16#aa#)) OR
 					(reg_q91 AND symb_decoder(16#09#)) OR
 					(reg_q91 AND symb_decoder(16#15#)) OR
 					(reg_q91 AND symb_decoder(16#4c#)) OR
 					(reg_q91 AND symb_decoder(16#d0#)) OR
 					(reg_q91 AND symb_decoder(16#dc#)) OR
 					(reg_q91 AND symb_decoder(16#ad#)) OR
 					(reg_q91 AND symb_decoder(16#ca#)) OR
 					(reg_q91 AND symb_decoder(16#60#)) OR
 					(reg_q91 AND symb_decoder(16#26#)) OR
 					(reg_q91 AND symb_decoder(16#e0#)) OR
 					(reg_q91 AND symb_decoder(16#ed#)) OR
 					(reg_q91 AND symb_decoder(16#40#)) OR
 					(reg_q91 AND symb_decoder(16#a5#)) OR
 					(reg_q91 AND symb_decoder(16#de#)) OR
 					(reg_q91 AND symb_decoder(16#d2#)) OR
 					(reg_q91 AND symb_decoder(16#c3#)) OR
 					(reg_q91 AND symb_decoder(16#3f#)) OR
 					(reg_q91 AND symb_decoder(16#fb#)) OR
 					(reg_q91 AND symb_decoder(16#fe#)) OR
 					(reg_q91 AND symb_decoder(16#f0#)) OR
 					(reg_q91 AND symb_decoder(16#e2#)) OR
 					(reg_q91 AND symb_decoder(16#51#)) OR
 					(reg_q91 AND symb_decoder(16#2a#)) OR
 					(reg_q91 AND symb_decoder(16#61#)) OR
 					(reg_q91 AND symb_decoder(16#e3#)) OR
 					(reg_q91 AND symb_decoder(16#fd#)) OR
 					(reg_q91 AND symb_decoder(16#28#)) OR
 					(reg_q91 AND symb_decoder(16#80#)) OR
 					(reg_q91 AND symb_decoder(16#82#)) OR
 					(reg_q91 AND symb_decoder(16#8a#)) OR
 					(reg_q91 AND symb_decoder(16#ae#)) OR
 					(reg_q91 AND symb_decoder(16#e4#)) OR
 					(reg_q91 AND symb_decoder(16#4b#)) OR
 					(reg_q91 AND symb_decoder(16#59#)) OR
 					(reg_q91 AND symb_decoder(16#70#)) OR
 					(reg_q91 AND symb_decoder(16#9c#)) OR
 					(reg_q91 AND symb_decoder(16#69#)) OR
 					(reg_q91 AND symb_decoder(16#da#)) OR
 					(reg_q91 AND symb_decoder(16#8b#)) OR
 					(reg_q91 AND symb_decoder(16#31#)) OR
 					(reg_q91 AND symb_decoder(16#91#)) OR
 					(reg_q91 AND symb_decoder(16#98#)) OR
 					(reg_q91 AND symb_decoder(16#16#)) OR
 					(reg_q91 AND symb_decoder(16#42#)) OR
 					(reg_q91 AND symb_decoder(16#bb#)) OR
 					(reg_q91 AND symb_decoder(16#c0#)) OR
 					(reg_q91 AND symb_decoder(16#62#)) OR
 					(reg_q91 AND symb_decoder(16#c9#)) OR
 					(reg_q91 AND symb_decoder(16#b5#)) OR
 					(reg_q91 AND symb_decoder(16#74#)) OR
 					(reg_q91 AND symb_decoder(16#4d#)) OR
 					(reg_q91 AND symb_decoder(16#f4#)) OR
 					(reg_q91 AND symb_decoder(16#b7#)) OR
 					(reg_q91 AND symb_decoder(16#85#)) OR
 					(reg_q91 AND symb_decoder(16#30#)) OR
 					(reg_q91 AND symb_decoder(16#6f#)) OR
 					(reg_q91 AND symb_decoder(16#77#));
reg_q91_init <= '0' ;
	p_reg_q91: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q91 <= reg_q91_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q91 <= reg_q91_init;
        else
          reg_q91 <= reg_q91_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph54

reg_q844_in <= (reg_q842 AND symb_decoder(16#32#)) OR
 					(reg_q842 AND symb_decoder(16#34#)) OR
 					(reg_q842 AND symb_decoder(16#36#)) OR
 					(reg_q842 AND symb_decoder(16#37#)) OR
 					(reg_q842 AND symb_decoder(16#38#)) OR
 					(reg_q842 AND symb_decoder(16#35#)) OR
 					(reg_q842 AND symb_decoder(16#39#)) OR
 					(reg_q842 AND symb_decoder(16#33#)) OR
 					(reg_q842 AND symb_decoder(16#30#)) OR
 					(reg_q842 AND symb_decoder(16#31#)) OR
 					(reg_q844 AND symb_decoder(16#37#)) OR
 					(reg_q844 AND symb_decoder(16#35#)) OR
 					(reg_q844 AND symb_decoder(16#39#)) OR
 					(reg_q844 AND symb_decoder(16#33#)) OR
 					(reg_q844 AND symb_decoder(16#32#)) OR
 					(reg_q844 AND symb_decoder(16#36#)) OR
 					(reg_q844 AND symb_decoder(16#38#)) OR
 					(reg_q844 AND symb_decoder(16#34#)) OR
 					(reg_q844 AND symb_decoder(16#30#)) OR
 					(reg_q844 AND symb_decoder(16#31#));
reg_q1645_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1644 AND symb_decoder(16#0a#)) OR
 					(reg_q1644 AND symb_decoder(16#0d#));
reg_q834_in <= (reg_q832 AND symb_decoder(16#2e#));
reg_q1882_in <= (reg_q1880 AND symb_decoder(16#35#)) OR
 					(reg_q1880 AND symb_decoder(16#39#)) OR
 					(reg_q1880 AND symb_decoder(16#30#)) OR
 					(reg_q1880 AND symb_decoder(16#36#)) OR
 					(reg_q1880 AND symb_decoder(16#37#)) OR
 					(reg_q1880 AND symb_decoder(16#31#)) OR
 					(reg_q1880 AND symb_decoder(16#33#)) OR
 					(reg_q1880 AND symb_decoder(16#32#)) OR
 					(reg_q1880 AND symb_decoder(16#38#)) OR
 					(reg_q1880 AND symb_decoder(16#34#)) OR
 					(reg_q1882 AND symb_decoder(16#30#)) OR
 					(reg_q1882 AND symb_decoder(16#38#)) OR
 					(reg_q1882 AND symb_decoder(16#34#)) OR
 					(reg_q1882 AND symb_decoder(16#39#)) OR
 					(reg_q1882 AND symb_decoder(16#36#)) OR
 					(reg_q1882 AND symb_decoder(16#33#)) OR
 					(reg_q1882 AND symb_decoder(16#35#)) OR
 					(reg_q1882 AND symb_decoder(16#37#)) OR
 					(reg_q1882 AND symb_decoder(16#31#)) OR
 					(reg_q1882 AND symb_decoder(16#32#));
reg_q620_in <= (reg_q618 AND symb_decoder(16#73#)) OR
 					(reg_q618 AND symb_decoder(16#53#));
reg_q2387_in <= (reg_q2385 AND symb_decoder(16#31#));
reg_q454_in <= (reg_q2695 AND symb_decoder(16#42#)) OR
 					(reg_q2695 AND symb_decoder(16#62#)) OR
 					(reg_q452 AND symb_decoder(16#62#)) OR
 					(reg_q452 AND symb_decoder(16#42#));
reg_q1197_in <= (reg_q2695 AND symb_decoder(16#66#)) OR
 					(reg_q2695 AND symb_decoder(16#46#)) OR
 					(reg_q1195 AND symb_decoder(16#46#)) OR
 					(reg_q1195 AND symb_decoder(16#66#));
reg_q846_in <= (reg_q844 AND symb_decoder(16#5e#));
reg_q2389_in <= (reg_q2387 AND symb_decoder(16#23#));
reg_fullgraph54_init <= "0000";

reg_fullgraph54_sel <= "000000" & reg_q2389_in & reg_q846_in & reg_q1197_in & reg_q454_in & reg_q2387_in & reg_q620_in & reg_q1882_in & reg_q834_in & reg_q1645_in & reg_q844_in;

	--coder fullgraph54
with reg_fullgraph54_sel select
reg_fullgraph54_in <=
	"0001" when "0000000000000001",
	"0010" when "0000000000000010",
	"0011" when "0000000000000100",
	"0100" when "0000000000001000",
	"0101" when "0000000000010000",
	"0110" when "0000000000100000",
	"0111" when "0000000001000000",
	"1000" when "0000000010000000",
	"1001" when "0000000100000000",
	"1010" when "0000001000000000",
	"0000" when others;
 --end coder

	p_reg_fullgraph54: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph54 <= reg_fullgraph54_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph54 <= reg_fullgraph54_init;
        else
          reg_fullgraph54 <= reg_fullgraph54_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph54

		reg_q844 <= '1' when reg_fullgraph54 = "0001" else '0'; 
		reg_q1645 <= '1' when reg_fullgraph54 = "0010" else '0'; 
		reg_q834 <= '1' when reg_fullgraph54 = "0011" else '0'; 
		reg_q1882 <= '1' when reg_fullgraph54 = "0100" else '0'; 
		reg_q620 <= '1' when reg_fullgraph54 = "0101" else '0'; 
		reg_q2387 <= '1' when reg_fullgraph54 = "0110" else '0'; 
		reg_q454 <= '1' when reg_fullgraph54 = "0111" else '0'; 
		reg_q1197 <= '1' when reg_fullgraph54 = "1000" else '0'; 
		reg_q846 <= '1' when reg_fullgraph54 = "1001" else '0'; 
		reg_q2389 <= '1' when reg_fullgraph54 = "1010" else '0'; 
--end decoder 
--######################################################
--fullgraph55

reg_q1768_in <= (reg_q1766 AND symb_decoder(16#0a#)) OR
 					(reg_q1766 AND symb_decoder(16#0c#)) OR
 					(reg_q1766 AND symb_decoder(16#0d#)) OR
 					(reg_q1766 AND symb_decoder(16#20#)) OR
 					(reg_q1766 AND symb_decoder(16#09#));
reg_q836_in <= (reg_q834 AND symb_decoder(16#37#)) OR
 					(reg_q834 AND symb_decoder(16#35#)) OR
 					(reg_q834 AND symb_decoder(16#32#)) OR
 					(reg_q834 AND symb_decoder(16#39#)) OR
 					(reg_q834 AND symb_decoder(16#33#)) OR
 					(reg_q834 AND symb_decoder(16#36#)) OR
 					(reg_q834 AND symb_decoder(16#30#)) OR
 					(reg_q834 AND symb_decoder(16#38#)) OR
 					(reg_q834 AND symb_decoder(16#31#)) OR
 					(reg_q834 AND symb_decoder(16#34#)) OR
 					(reg_q836 AND symb_decoder(16#33#)) OR
 					(reg_q836 AND symb_decoder(16#36#)) OR
 					(reg_q836 AND symb_decoder(16#37#)) OR
 					(reg_q836 AND symb_decoder(16#30#)) OR
 					(reg_q836 AND symb_decoder(16#39#)) OR
 					(reg_q836 AND symb_decoder(16#34#)) OR
 					(reg_q836 AND symb_decoder(16#35#)) OR
 					(reg_q836 AND symb_decoder(16#32#)) OR
 					(reg_q836 AND symb_decoder(16#31#)) OR
 					(reg_q836 AND symb_decoder(16#38#));
reg_q838_in <= (reg_q836 AND symb_decoder(16#2e#));
reg_q1828_in <= (reg_q2695 AND symb_decoder(16#53#)) OR
 					(reg_q2695 AND symb_decoder(16#73#)) OR
 					(reg_q1826 AND symb_decoder(16#53#)) OR
 					(reg_q1826 AND symb_decoder(16#73#));
reg_fullgraph55_init <= "000";

reg_fullgraph55_sel <= "0000" & reg_q1828_in & reg_q838_in & reg_q836_in & reg_q1768_in;

	--coder fullgraph55
with reg_fullgraph55_sel select
reg_fullgraph55_in <=
	"001" when "00000001",
	"010" when "00000010",
	"011" when "00000100",
	"100" when "00001000",
	"000" when others;
 --end coder

	p_reg_fullgraph55: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph55 <= reg_fullgraph55_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph55 <= reg_fullgraph55_init;
        else
          reg_fullgraph55 <= reg_fullgraph55_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph55

		reg_q1768 <= '1' when reg_fullgraph55 = "001" else '0'; 
		reg_q836 <= '1' when reg_fullgraph55 = "010" else '0'; 
		reg_q838 <= '1' when reg_fullgraph55 = "011" else '0'; 
		reg_q1828 <= '1' when reg_fullgraph55 = "100" else '0'; 
--end decoder 
--######################################################
--fullgraph56

reg_q817_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q816 AND symb_decoder(16#0a#)) OR
 					(reg_q816 AND symb_decoder(16#0d#));
reg_q840_in <= (reg_q838 AND symb_decoder(16#33#)) OR
 					(reg_q838 AND symb_decoder(16#36#)) OR
 					(reg_q838 AND symb_decoder(16#35#)) OR
 					(reg_q838 AND symb_decoder(16#31#)) OR
 					(reg_q838 AND symb_decoder(16#39#)) OR
 					(reg_q838 AND symb_decoder(16#34#)) OR
 					(reg_q838 AND symb_decoder(16#32#)) OR
 					(reg_q838 AND symb_decoder(16#38#)) OR
 					(reg_q838 AND symb_decoder(16#37#)) OR
 					(reg_q838 AND symb_decoder(16#30#)) OR
 					(reg_q840 AND symb_decoder(16#35#)) OR
 					(reg_q840 AND symb_decoder(16#32#)) OR
 					(reg_q840 AND symb_decoder(16#33#)) OR
 					(reg_q840 AND symb_decoder(16#34#)) OR
 					(reg_q840 AND symb_decoder(16#38#)) OR
 					(reg_q840 AND symb_decoder(16#37#)) OR
 					(reg_q840 AND symb_decoder(16#31#)) OR
 					(reg_q840 AND symb_decoder(16#36#)) OR
 					(reg_q840 AND symb_decoder(16#39#)) OR
 					(reg_q840 AND symb_decoder(16#30#));
reg_fullgraph56_init <= "00";

reg_fullgraph56_sel <= "00" & reg_q840_in & reg_q817_in;

	--coder fullgraph56
with reg_fullgraph56_sel select
reg_fullgraph56_in <=
	"01" when "0001",
	"10" when "0010",
	"00" when others;
 --end coder

	p_reg_fullgraph56: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph56 <= reg_fullgraph56_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph56 <= reg_fullgraph56_init;
        else
          reg_fullgraph56 <= reg_fullgraph56_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph56

		reg_q817 <= '1' when reg_fullgraph56 = "01" else '0'; 
		reg_q840 <= '1' when reg_fullgraph56 = "10" else '0'; 
--end decoder 
--######################################################
--fullgraph57

reg_q1782_in <= (reg_q1780 AND symb_decoder(16#20#)) OR
 					(reg_q1780 AND symb_decoder(16#09#)) OR
 					(reg_q1780 AND symb_decoder(16#0a#)) OR
 					(reg_q1780 AND symb_decoder(16#0c#)) OR
 					(reg_q1780 AND symb_decoder(16#0d#));
reg_q2_in <= (reg_q2695 AND symb_decoder(16#30#)) OR
 					(reg_q0 AND symb_decoder(16#30#));
reg_fullgraph57_init <= "00";

reg_fullgraph57_sel <= "00" & reg_q2_in & reg_q1782_in;

	--coder fullgraph57
with reg_fullgraph57_sel select
reg_fullgraph57_in <=
	"01" when "0001",
	"10" when "0010",
	"00" when others;
 --end coder

	p_reg_fullgraph57: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph57 <= reg_fullgraph57_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph57 <= reg_fullgraph57_init;
        else
          reg_fullgraph57 <= reg_fullgraph57_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph57

		reg_q1782 <= '1' when reg_fullgraph57 = "01" else '0'; 
		reg_q2 <= '1' when reg_fullgraph57 = "10" else '0'; 
--end decoder 
--######################################################
--fullgraph58

reg_q1784_in <= (reg_q1782 AND symb_decoder(16#0c#)) OR
 					(reg_q1782 AND symb_decoder(16#0a#)) OR
 					(reg_q1782 AND symb_decoder(16#20#)) OR
 					(reg_q1782 AND symb_decoder(16#09#)) OR
 					(reg_q1782 AND symb_decoder(16#0d#));
reg_q4_in <= (reg_q2 AND symb_decoder(16#30#));
reg_fullgraph58_init <= "00";

reg_fullgraph58_sel <= "00" & reg_q4_in & reg_q1784_in;

	--coder fullgraph58
with reg_fullgraph58_sel select
reg_fullgraph58_in <=
	"01" when "0001",
	"10" when "0010",
	"00" when others;
 --end coder

	p_reg_fullgraph58: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph58 <= reg_fullgraph58_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph58 <= reg_fullgraph58_init;
        else
          reg_fullgraph58 <= reg_fullgraph58_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph58

		reg_q1784 <= '1' when reg_fullgraph58 = "01" else '0'; 
		reg_q4 <= '1' when reg_fullgraph58 = "10" else '0'; 
--end decoder 
--######################################################
--fullgraph59

reg_q2092_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2091 AND symb_decoder(16#0a#)) OR
 					(reg_q2091 AND symb_decoder(16#0d#));
reg_q6_in <= (reg_q4 AND symb_decoder(16#30#));
reg_fullgraph59_init <= "00";

reg_fullgraph59_sel <= "00" & reg_q6_in & reg_q2092_in;

	--coder fullgraph59
with reg_fullgraph59_sel select
reg_fullgraph59_in <=
	"01" when "0001",
	"10" when "0010",
	"00" when others;
 --end coder

	p_reg_fullgraph59: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph59 <= reg_fullgraph59_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph59 <= reg_fullgraph59_init;
        else
          reg_fullgraph59 <= reg_fullgraph59_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph59

		reg_q2092 <= '1' when reg_fullgraph59 = "01" else '0'; 
		reg_q6 <= '1' when reg_fullgraph59 = "10" else '0'; 
--end decoder 

reg_q1225_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1224 AND symb_decoder(16#0a#)) OR
 					(reg_q1224 AND symb_decoder(16#0d#));
reg_q1225_init <= '0' ;
	p_reg_q1225: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1225 <= reg_q1225_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1225 <= reg_q1225_init;
        else
          reg_q1225 <= reg_q1225_in;
        end if;
      end if;
    end if;
  end process;

	--######################################################
--fullgraph61

reg_q2583_in <= (reg_q2579 AND symb_decoder(16#0d#)) OR
 					(reg_q2615 AND symb_decoder(16#0d#));
reg_q2585_in <= (reg_q2583 AND symb_decoder(16#0a#));
reg_fullgraph61_init <= "00";

reg_fullgraph61_sel <= "00" & reg_q2585_in & reg_q2583_in;

	--coder fullgraph61
with reg_fullgraph61_sel select
reg_fullgraph61_in <=
	"01" when "0001",
	"10" when "0010",
	"00" when others;
 --end coder

	p_reg_fullgraph61: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_fullgraph61 <= reg_fullgraph61_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_fullgraph61 <= reg_fullgraph61_init;
        else
          reg_fullgraph61 <= reg_fullgraph61_in;
        end if;
      end if;
    end if;
  end process;

	-- docoder fullgraph61

		reg_q2583 <= '1' when reg_fullgraph61 = "01" else '0'; 
		reg_q2585 <= '1' when reg_fullgraph61 = "10" else '0'; 
--end decoder 

reg_q2001_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2000 AND symb_decoder(16#0a#)) OR
 					(reg_q2000 AND symb_decoder(16#0d#));
reg_q2001_init <= '0' ;
	p_reg_q2001: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2001 <= reg_q2001_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2001 <= reg_q2001_init;
        else
          reg_q2001 <= reg_q2001_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q681_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q680 AND symb_decoder(16#0d#)) OR
 					(reg_q680 AND symb_decoder(16#0a#));
reg_q681_init <= '0' ;
	p_reg_q681: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q681 <= reg_q681_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q681 <= reg_q681_init;
        else
          reg_q681 <= reg_q681_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1754_in <= (reg_q1752 AND symb_decoder(16#0d#)) OR
 					(reg_q1752 AND symb_decoder(16#20#)) OR
 					(reg_q1752 AND symb_decoder(16#0c#)) OR
 					(reg_q1752 AND symb_decoder(16#09#)) OR
 					(reg_q1752 AND symb_decoder(16#0a#));
reg_q1754_init <= '0' ;
	p_reg_q1754: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1754 <= reg_q1754_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1754 <= reg_q1754_init;
        else
          reg_q1754 <= reg_q1754_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1756_in <= (reg_q1754 AND symb_decoder(16#0a#)) OR
 					(reg_q1754 AND symb_decoder(16#20#)) OR
 					(reg_q1754 AND symb_decoder(16#09#)) OR
 					(reg_q1754 AND symb_decoder(16#0c#)) OR
 					(reg_q1754 AND symb_decoder(16#0d#));
reg_q1756_init <= '0' ;
	p_reg_q1756: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1756 <= reg_q1756_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1756 <= reg_q1756_init;
        else
          reg_q1756 <= reg_q1756_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q959_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q958 AND symb_decoder(16#0a#)) OR
 					(reg_q958 AND symb_decoder(16#0d#));
reg_q959_init <= '0' ;
	p_reg_q959: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q959 <= reg_q959_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q959 <= reg_q959_init;
        else
          reg_q959 <= reg_q959_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q900_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q899 AND symb_decoder(16#0d#)) OR
 					(reg_q899 AND symb_decoder(16#0a#));
reg_q900_init <= '0' ;
	p_reg_q900: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q900 <= reg_q900_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q900 <= reg_q900_init;
        else
          reg_q900 <= reg_q900_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q304_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q303 AND symb_decoder(16#0a#)) OR
 					(reg_q303 AND symb_decoder(16#0d#));
reg_q304_init <= '0' ;
	p_reg_q304: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q304 <= reg_q304_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q304 <= reg_q304_init;
        else
          reg_q304 <= reg_q304_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1786_in <= (reg_q1784 AND symb_decoder(16#09#)) OR
 					(reg_q1784 AND symb_decoder(16#20#)) OR
 					(reg_q1784 AND symb_decoder(16#0a#)) OR
 					(reg_q1784 AND symb_decoder(16#0c#)) OR
 					(reg_q1784 AND symb_decoder(16#0d#));
reg_q1786_init <= '0' ;
	p_reg_q1786: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1786 <= reg_q1786_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1786 <= reg_q1786_init;
        else
          reg_q1786 <= reg_q1786_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1788_in <= (reg_q1786 AND symb_decoder(16#0a#)) OR
 					(reg_q1786 AND symb_decoder(16#0c#)) OR
 					(reg_q1786 AND symb_decoder(16#09#)) OR
 					(reg_q1786 AND symb_decoder(16#0d#)) OR
 					(reg_q1786 AND symb_decoder(16#20#));
reg_q1788_init <= '0' ;
	p_reg_q1788: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1788 <= reg_q1788_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1788 <= reg_q1788_init;
        else
          reg_q1788 <= reg_q1788_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1746_in <= (reg_q1744 AND symb_decoder(16#0d#)) OR
 					(reg_q1744 AND symb_decoder(16#20#)) OR
 					(reg_q1744 AND symb_decoder(16#0c#)) OR
 					(reg_q1744 AND symb_decoder(16#09#)) OR
 					(reg_q1744 AND symb_decoder(16#0a#));
reg_q1746_init <= '0' ;
	p_reg_q1746: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1746 <= reg_q1746_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1746 <= reg_q1746_init;
        else
          reg_q1746 <= reg_q1746_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1748_in <= (reg_q1746 AND symb_decoder(16#0a#)) OR
 					(reg_q1746 AND symb_decoder(16#0d#)) OR
 					(reg_q1746 AND symb_decoder(16#20#)) OR
 					(reg_q1746 AND symb_decoder(16#0c#)) OR
 					(reg_q1746 AND symb_decoder(16#09#));
reg_q1748_init <= '0' ;
	p_reg_q1748: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1748 <= reg_q1748_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1748 <= reg_q1748_init;
        else
          reg_q1748 <= reg_q1748_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1051_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1050 AND symb_decoder(16#0d#)) OR
 					(reg_q1050 AND symb_decoder(16#0a#));
reg_q1051_init <= '0' ;
	p_reg_q1051: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1051 <= reg_q1051_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1051 <= reg_q1051_init;
        else
          reg_q1051 <= reg_q1051_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1764_in <= (reg_q1762 AND symb_decoder(16#0c#)) OR
 					(reg_q1762 AND symb_decoder(16#0a#)) OR
 					(reg_q1762 AND symb_decoder(16#20#)) OR
 					(reg_q1762 AND symb_decoder(16#09#)) OR
 					(reg_q1762 AND symb_decoder(16#0d#));
reg_q1764_init <= '0' ;
	p_reg_q1764: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1764 <= reg_q1764_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1764 <= reg_q1764_init;
        else
          reg_q1764 <= reg_q1764_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1766_in <= (reg_q1764 AND symb_decoder(16#0a#)) OR
 					(reg_q1764 AND symb_decoder(16#09#)) OR
 					(reg_q1764 AND symb_decoder(16#0d#)) OR
 					(reg_q1764 AND symb_decoder(16#20#)) OR
 					(reg_q1764 AND symb_decoder(16#0c#));
reg_q1766_init <= '0' ;
	p_reg_q1766: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1766 <= reg_q1766_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1766 <= reg_q1766_init;
        else
          reg_q1766 <= reg_q1766_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1453_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1452 AND symb_decoder(16#0a#)) OR
 					(reg_q1452 AND symb_decoder(16#0d#));
reg_q1453_init <= '0' ;
	p_reg_q1453: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1453 <= reg_q1453_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1453 <= reg_q1453_init;
        else
          reg_q1453 <= reg_q1453_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1744_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#09#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2695 AND symb_decoder(16#0c#)) OR
 					(reg_q2695 AND symb_decoder(16#20#)) OR
 					(reg_q1742 AND symb_decoder(16#0a#)) OR
 					(reg_q1742 AND symb_decoder(16#0d#)) OR
 					(reg_q1742 AND symb_decoder(16#0c#)) OR
 					(reg_q1742 AND symb_decoder(16#09#)) OR
 					(reg_q1742 AND symb_decoder(16#20#));
reg_q1744_init <= '0' ;
	p_reg_q1744: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1744 <= reg_q1744_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1744 <= reg_q1744_init;
        else
          reg_q1744 <= reg_q1744_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1774_in <= (reg_q1772 AND symb_decoder(16#09#)) OR
 					(reg_q1772 AND symb_decoder(16#20#)) OR
 					(reg_q1772 AND symb_decoder(16#0c#)) OR
 					(reg_q1772 AND symb_decoder(16#0d#)) OR
 					(reg_q1772 AND symb_decoder(16#0a#));
reg_q1774_init <= '0' ;
	p_reg_q1774: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1774 <= reg_q1774_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1774 <= reg_q1774_init;
        else
          reg_q1774 <= reg_q1774_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1776_in <= (reg_q1774 AND symb_decoder(16#0a#)) OR
 					(reg_q1774 AND symb_decoder(16#0d#)) OR
 					(reg_q1774 AND symb_decoder(16#20#)) OR
 					(reg_q1774 AND symb_decoder(16#0c#)) OR
 					(reg_q1774 AND symb_decoder(16#09#));
reg_q1776_init <= '0' ;
	p_reg_q1776: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1776 <= reg_q1776_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1776 <= reg_q1776_init;
        else
          reg_q1776 <= reg_q1776_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1014_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1013 AND symb_decoder(16#0a#)) OR
 					(reg_q1013 AND symb_decoder(16#0d#));
reg_q1014_init <= '0' ;
	p_reg_q1014: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1014 <= reg_q1014_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1014 <= reg_q1014_init;
        else
          reg_q1014 <= reg_q1014_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1545_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1544 AND symb_decoder(16#0d#)) OR
 					(reg_q1544 AND symb_decoder(16#0a#));
reg_q1545_init <= '0' ;
	p_reg_q1545: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1545 <= reg_q1545_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1545 <= reg_q1545_init;
        else
          reg_q1545 <= reg_q1545_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1780_in <= (reg_q1778 AND symb_decoder(16#20#)) OR
 					(reg_q1778 AND symb_decoder(16#09#)) OR
 					(reg_q1778 AND symb_decoder(16#0a#)) OR
 					(reg_q1778 AND symb_decoder(16#0d#)) OR
 					(reg_q1778 AND symb_decoder(16#0c#));
reg_q1780_init <= '0' ;
	p_reg_q1780: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1780 <= reg_q1780_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1780 <= reg_q1780_init;
        else
          reg_q1780 <= reg_q1780_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2619_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2618 AND symb_decoder(16#0a#)) OR
 					(reg_q2618 AND symb_decoder(16#0d#));
reg_q2619_init <= '0' ;
	p_reg_q2619: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2619 <= reg_q2619_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2619 <= reg_q2619_init;
        else
          reg_q2619 <= reg_q2619_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q666_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q665 AND symb_decoder(16#0d#)) OR
 					(reg_q665 AND symb_decoder(16#0a#));
reg_q666_init <= '0' ;
	p_reg_q666: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q666 <= reg_q666_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q666 <= reg_q666_init;
        else
          reg_q666 <= reg_q666_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2324_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2323 AND symb_decoder(16#0a#)) OR
 					(reg_q2323 AND symb_decoder(16#0d#));
reg_q2324_init <= '0' ;
	p_reg_q2324: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2324 <= reg_q2324_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2324 <= reg_q2324_init;
        else
          reg_q2324 <= reg_q2324_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1752_in <= (reg_q1750 AND symb_decoder(16#0c#)) OR
 					(reg_q1750 AND symb_decoder(16#0d#)) OR
 					(reg_q1750 AND symb_decoder(16#09#)) OR
 					(reg_q1750 AND symb_decoder(16#20#)) OR
 					(reg_q1750 AND symb_decoder(16#0a#));
reg_q1752_init <= '0' ;
	p_reg_q1752: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1752 <= reg_q1752_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1752 <= reg_q1752_init;
        else
          reg_q1752 <= reg_q1752_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q704_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q703 AND symb_decoder(16#0d#)) OR
 					(reg_q703 AND symb_decoder(16#0a#));
reg_q704_init <= '0' ;
	p_reg_q704: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q704 <= reg_q704_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q704 <= reg_q704_init;
        else
          reg_q704 <= reg_q704_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1522_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1521 AND symb_decoder(16#0d#)) OR
 					(reg_q1521 AND symb_decoder(16#0a#));
reg_q1522_init <= '0' ;
	p_reg_q1522: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1522 <= reg_q1522_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1522 <= reg_q1522_init;
        else
          reg_q1522 <= reg_q1522_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1956_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1955 AND symb_decoder(16#0a#)) OR
 					(reg_q1955 AND symb_decoder(16#0d#));
reg_q1956_init <= '0' ;
	p_reg_q1956: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1956 <= reg_q1956_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1956 <= reg_q1956_init;
        else
          reg_q1956 <= reg_q1956_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2534_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2533 AND symb_decoder(16#0d#)) OR
 					(reg_q2533 AND symb_decoder(16#0a#));
reg_q2534_init <= '0' ;
	p_reg_q2534: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2534 <= reg_q2534_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2534 <= reg_q2534_init;
        else
          reg_q2534 <= reg_q2534_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q780_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q779 AND symb_decoder(16#0d#)) OR
 					(reg_q779 AND symb_decoder(16#0a#));
reg_q780_init <= '0' ;
	p_reg_q780: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q780 <= reg_q780_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q780 <= reg_q780_init;
        else
          reg_q780 <= reg_q780_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q715_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q714 AND symb_decoder(16#0a#)) OR
 					(reg_q714 AND symb_decoder(16#0d#));
reg_q715_init <= '0' ;
	p_reg_q715: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q715 <= reg_q715_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q715 <= reg_q715_init;
        else
          reg_q715 <= reg_q715_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1778_in <= (reg_q1776 AND symb_decoder(16#09#)) OR
 					(reg_q1776 AND symb_decoder(16#0d#)) OR
 					(reg_q1776 AND symb_decoder(16#0a#)) OR
 					(reg_q1776 AND symb_decoder(16#0c#)) OR
 					(reg_q1776 AND symb_decoder(16#20#));
reg_q1778_init <= '0' ;
	p_reg_q1778: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1778 <= reg_q1778_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1778 <= reg_q1778_init;
        else
          reg_q1778 <= reg_q1778_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1604_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q1603 AND symb_decoder(16#0d#)) OR
 					(reg_q1603 AND symb_decoder(16#0a#));
reg_q1604_init <= '0' ;
	p_reg_q1604: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1604 <= reg_q1604_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1604 <= reg_q1604_init;
        else
          reg_q1604 <= reg_q1604_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2212_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2211 AND symb_decoder(16#0d#)) OR
 					(reg_q2211 AND symb_decoder(16#0a#));
reg_q2212_init <= '0' ;
	p_reg_q2212: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2212 <= reg_q2212_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2212 <= reg_q2212_init;
        else
          reg_q2212 <= reg_q2212_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q226_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q225 AND symb_decoder(16#0a#)) OR
 					(reg_q225 AND symb_decoder(16#0d#));
reg_q226_init <= '0' ;
	p_reg_q226: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q226 <= reg_q226_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q226 <= reg_q226_init;
        else
          reg_q226 <= reg_q226_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2125_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2124 AND symb_decoder(16#0d#)) OR
 					(reg_q2124 AND symb_decoder(16#0a#));
reg_q2125_init <= '0' ;
	p_reg_q2125: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2125 <= reg_q2125_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2125 <= reg_q2125_init;
        else
          reg_q2125 <= reg_q2125_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q47_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q46 AND symb_decoder(16#0a#)) OR
 					(reg_q46 AND symb_decoder(16#0d#));
reg_q47_init <= '0' ;
	p_reg_q47: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q47 <= reg_q47_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q47 <= reg_q47_init;
        else
          reg_q47 <= reg_q47_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1762_in <= (reg_q1760 AND symb_decoder(16#20#)) OR
 					(reg_q1760 AND symb_decoder(16#09#)) OR
 					(reg_q1760 AND symb_decoder(16#0a#)) OR
 					(reg_q1760 AND symb_decoder(16#0c#)) OR
 					(reg_q1760 AND symb_decoder(16#0d#));
reg_q1762_init <= '0' ;
	p_reg_q1762: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1762 <= reg_q1762_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1762 <= reg_q1762_init;
        else
          reg_q1762 <= reg_q1762_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1760_in <= (reg_q1758 AND symb_decoder(16#0c#)) OR
 					(reg_q1758 AND symb_decoder(16#20#)) OR
 					(reg_q1758 AND symb_decoder(16#09#)) OR
 					(reg_q1758 AND symb_decoder(16#0d#)) OR
 					(reg_q1758 AND symb_decoder(16#0a#));
reg_q1760_init <= '0' ;
	p_reg_q1760: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1760 <= reg_q1760_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1760 <= reg_q1760_init;
        else
          reg_q1760 <= reg_q1760_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q415_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q414 AND symb_decoder(16#0a#)) OR
 					(reg_q414 AND symb_decoder(16#0d#));
reg_q415_init <= '0' ;
	p_reg_q415: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q415 <= reg_q415_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q415 <= reg_q415_init;
        else
          reg_q415 <= reg_q415_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q179_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q178 AND symb_decoder(16#0a#)) OR
 					(reg_q178 AND symb_decoder(16#0d#));
reg_q179_init <= '0' ;
	p_reg_q179: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q179 <= reg_q179_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q179 <= reg_q179_init;
        else
          reg_q179 <= reg_q179_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1758_in <= (reg_q1756 AND symb_decoder(16#0a#)) OR
 					(reg_q1756 AND symb_decoder(16#09#)) OR
 					(reg_q1756 AND symb_decoder(16#0d#)) OR
 					(reg_q1756 AND symb_decoder(16#20#)) OR
 					(reg_q1756 AND symb_decoder(16#0c#));
reg_q1758_init <= '0' ;
	p_reg_q1758: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1758 <= reg_q1758_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1758 <= reg_q1758_init;
        else
          reg_q1758 <= reg_q1758_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q1750_in <= (reg_q1748 AND symb_decoder(16#0d#)) OR
 					(reg_q1748 AND symb_decoder(16#0c#)) OR
 					(reg_q1748 AND symb_decoder(16#09#)) OR
 					(reg_q1748 AND symb_decoder(16#0a#)) OR
 					(reg_q1748 AND symb_decoder(16#20#));
reg_q1750_init <= '0' ;
	p_reg_q1750: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q1750 <= reg_q1750_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q1750 <= reg_q1750_init;
        else
          reg_q1750 <= reg_q1750_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q2253_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q2252 AND symb_decoder(16#0d#)) OR
 					(reg_q2252 AND symb_decoder(16#0a#));
reg_q2253_init <= '0' ;
	p_reg_q2253: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q2253 <= reg_q2253_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q2253 <= reg_q2253_init;
        else
          reg_q2253 <= reg_q2253_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q263_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q262 AND symb_decoder(16#0a#)) OR
 					(reg_q262 AND symb_decoder(16#0d#));
reg_q263_init <= '0' ;
	p_reg_q263: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q263 <= reg_q263_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q263 <= reg_q263_init;
        else
          reg_q263 <= reg_q263_in;
        end if;
      end if;
    end if;
  end process;

	
reg_q92_in <= (reg_q2695 AND symb_decoder(16#0a#)) OR
 					(reg_q2695 AND symb_decoder(16#0d#)) OR
 					(reg_q91 AND symb_decoder(16#0a#)) OR
 					(reg_q91 AND symb_decoder(16#0d#));
reg_q92_init <= '0' ;
	p_reg_q92: process (CLK)
	begin
    if (rising_edge(CLK)) then
      if (RESET = '1') then
        reg_q92 <= reg_q92_init;
      elsif (INPUT_EN = '1') then
        if (initialize = '1') then
          reg_q92 <= reg_q92_init;
        else
          reg_q92 <= reg_q92_in;
        end if;
      end if;
    end if;
  end process;

	
FINAL <= reg_q2692 OR reg_q677 OR reg_q1357 OR reg_q222 OR reg_q887 OR reg_q1952 OR reg_q776 OR reg_q1108 OR reg_q2206 OR reg_q2530 OR reg_q1824 OR reg_q953 OR reg_q2249 OR reg_q175 OR reg_q2050 OR reg_q88 OR reg_q662 OR reg_q2088 OR reg_q1541 OR reg_q846 OR reg_q1010 OR reg_q2320 OR reg_q1047 OR reg_q2482 OR reg_q44 OR reg_q700 OR reg_q1641 OR reg_q884 OR reg_q886 OR reg_q1449 OR reg_q2693 OR reg_q1221 OR reg_q259 OR reg_q1882 OR reg_q1294 OR reg_q411 OR reg_q2499 OR reg_q450 OR reg_q1995 OR reg_q1600 OR reg_q1193 OR reg_q2381 OR reg_q711 OR reg_q2465 OR reg_q2516 OR reg_q1740 OR reg_q554 OR reg_q300 OR reg_q1518 OR reg_q2121 OR reg_q2613 OR reg_q811;

	end architecture;
	